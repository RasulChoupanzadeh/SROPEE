* netlist generated with reverse MNA (number of voltage nodes: n = 144 )

.subckt equivalent_circuit

.param Ip1=1.0
.param Ip2=0.0
.param Ip3=0.0
.param Ip4=0.0

R1_1 V1 0 32843.0402864659
L1_1 V1 0 -3.2683358511908536e-10
C1_1 V1 0 2.413122947767331e-20

R1_2 V1 V2 52746231.549958125
L1_2 V1 V2 3.377887859248032e-05
C1_2 V1 V2 5.218874220682939e-23

R1_3 V1 V3 55846958.12957377
L1_3 V1 V3 1.2773824244766557e-05
C1_3 V1 V3 6.340278024200601e-23

R1_4 V1 V4 1073903185.2679036
L1_4 V1 V4 -1.7089623545141273e-05
C1_4 V1 V4 -2.4779152142870276e-23

R1_5 V1 V5 39595823.58352275
L1_5 V1 V5 -4.953740355020192e-08
C1_5 V1 V5 4.7202834206554005e-22

R1_6 V1 V6 11876006.411692316
L1_6 V1 V6 -1.308532442027404e-07
C1_6 V1 V6 -4.8306810156974107e-23

R1_7 V1 V7 142854975.01257032
L1_7 V1 V7 -1.5661352116073642e-06
C1_7 V1 V7 -5.963528942100693e-23

R1_8 V1 V8 22347140.48280149
L1_8 V1 V8 -1.1242992224486767e-07
C1_8 V1 V8 -3.439074131351262e-24

R1_9 V1 V9 -3830371.283593005
L1_9 V1 V9 -4.2192042035348874e-08
C1_9 V1 V9 -7.0941876418658755e-22

R1_10 V1 V10 81862704.53255837
L1_10 V1 V10 -4.2902233061870526e-07
C1_10 V1 V10 -8.049765475240366e-23

R1_11 V1 V11 -11978107.580503395
L1_11 V1 V11 -1.8159068499283704e-07
C1_11 V1 V11 -3.066695818799467e-22

R1_12 V1 V12 17144316.841018423
L1_12 V1 V12 6.481633826966991e-07
C1_12 V1 V12 9.12617197836186e-23

R1_13 V1 V13 -23818939.320242733
L1_13 V1 V13 -4.1208014760443834e-07
C1_13 V1 V13 1.0315661260393875e-22

R1_14 V1 V14 -64085881.18066183
L1_14 V1 V14 -7.084755535098106e-08
C1_14 V1 V14 -9.240417432989018e-23

R1_15 V1 V15 -26148326.513522975
L1_15 V1 V15 9.030389371508235e-07
C1_15 V1 V15 9.819553969537997e-23

R1_16 V1 V16 28725601.65227746
L1_16 V1 V16 -1.7694226864621593e-07
C1_16 V1 V16 2.5280422695212385e-23

R1_17 V1 V17 -7737485.838298803
L1_17 V1 V17 -3.756981512569454e-08
C1_17 V1 V17 1.3260301880256477e-22

R1_18 V1 V18 28303821.530887716
L1_18 V1 V18 -1.1952584288634779e-07
C1_18 V1 V18 -9.044989230821744e-23

R1_19 V1 V19 32691149.42204199
L1_19 V1 V19 -3.377562771398995e-08
C1_19 V1 V19 -3.659451689476625e-23

R1_20 V1 V20 21018648.695964266
L1_20 V1 V20 2.3630958950740225e-06
C1_20 V1 V20 -4.667415912773751e-24

R1_21 V1 V21 -7721284.765304409
L1_21 V1 V21 -7.411191718861069e-09
C1_21 V1 V21 -3.7256520888592416e-22

R1_22 V1 V22 29979587.248830955
L1_22 V1 V22 5.593646770029751e-08
C1_22 V1 V22 7.818970239421136e-23

R1_23 V1 V23 24757414.871199075
L1_23 V1 V23 6.506306370383417e-08
C1_23 V1 V23 1.3888522168740076e-22

R1_24 V1 V24 -50949061.22582886
L1_24 V1 V24 6.775758599486506e-08
C1_24 V1 V24 3.22900875993766e-23

R1_25 V1 V25 -16037777.282747775
L1_25 V1 V25 -1.662041461838372e-08
C1_25 V1 V25 -1.1436112666839887e-22

R1_26 V1 V26 25348243.415124003
L1_26 V1 V26 3.381828792779876e-07
C1_26 V1 V26 2.5107777253852702e-23

R1_27 V1 V27 38167232.45303551
L1_27 V1 V27 -3.6556393978432413e-07
C1_27 V1 V27 -1.136375887012821e-23

R1_28 V1 V28 12785431.786010666
L1_28 V1 V28 -1.095841863446447e-07
C1_28 V1 V28 7.263239261721158e-23

R1_29 V1 V29 4767414.027291174
L1_29 V1 V29 -9.832199228978045e-09
C1_29 V1 V29 1.357856585738304e-21

R1_30 V1 V30 76634896.97649817
L1_30 V1 V30 1.548260879302392e-07
C1_30 V1 V30 2.5315726162596637e-22

R1_31 V1 V31 9285072.272722468
L1_31 V1 V31 2.5618761654576376e-07
C1_31 V1 V31 3.832001796214252e-22

R1_32 V1 V32 -32779524.522479124
L1_32 V1 V32 1.2775889139842765e-07
C1_32 V1 V32 1.8766193819271925e-22

R1_33 V1 V33 -1097104.8601660826
L1_33 V1 V33 9.457348506474313e-09
C1_33 V1 V33 -1.829969141161941e-21

R1_34 V1 V34 2862722.169757503
L1_34 V1 V34 -2.5454722643384352e-08
C1_34 V1 V34 6.365146291089391e-22

R1_35 V1 V35 -2297700.406509519
L1_35 V1 V35 1.926871479372199e-08
C1_35 V1 V35 -1.107599839494037e-21

R1_36 V1 V36 5657132.812822665
L1_36 V1 V36 -4.237479404587872e-08
C1_36 V1 V36 1.6736863499499677e-22

R1_37 V1 V37 394231.43870306155
L1_37 V1 V37 -3.23330206204262e-09
C1_37 V1 V37 3.547840122995965e-21

R1_38 V1 V38 4291661.665044182
L1_38 V1 V38 -4.751699414819809e-08
C1_38 V1 V38 4.445516001488064e-23

R1_39 V1 V39 462298.1560930216
L1_39 V1 V39 -4.038869785419193e-09
C1_39 V1 V39 3.3368816057279373e-21

R1_40 V1 V40 6443175.383367595
L1_40 V1 V40 -5.703214977069511e-08
C1_40 V1 V40 2.1014761525213256e-22

R1_41 V1 V41 -112448.69088801344
L1_41 V1 V41 1.0175553356385538e-09
C1_41 V1 V41 -1.0559029253680108e-20

R1_42 V1 V42 -162841.24951230598
L1_42 V1 V42 1.4093739335828762e-09
C1_42 V1 V42 -8.345320248889722e-21

R1_43 V1 V43 -339376.3408647539
L1_43 V1 V43 2.925824996808596e-09
C1_43 V1 V43 -4.329345820682894e-21

R1_44 V1 V44 -17097648.764627084
L1_44 V1 V44 5.888259096231997e-08
C1_44 V1 V44 -6.028264627530951e-22

R1_45 V1 V45 360380.5431202822
L1_45 V1 V45 -2.8881873726576103e-09
C1_45 V1 V45 7.311748305114879e-21

R1_46 V1 V46 4162729.48508862
L1_46 V1 V46 -2.2709836450352162e-08
C1_46 V1 V46 2.928240534139445e-21

R1_47 V1 V47 -2052720.7638654984
L1_47 V1 V47 2.99583985503418e-08
C1_47 V1 V47 1.2738224478480188e-21

R1_48 V1 V48 1840186.642111468
L1_48 V1 V48 -1.6472831726292553e-08
C1_48 V1 V48 6.176438458964502e-22

R1_49 V1 V49 1791480.8531026542
L1_49 V1 V49 -2.9357910007834206e-08
C1_49 V1 V49 -2.020744562568901e-21

R1_50 V1 V50 -1256178.4098370196
L1_50 V1 V50 1.0243753678731118e-08
C1_50 V1 V50 -1.77973650693799e-21

R1_51 V1 V51 747848.2572784391
L1_51 V1 V51 -6.840369517497027e-09
C1_51 V1 V51 1.499752578020112e-21

R1_52 V1 V52 -1776777.1076365134
L1_52 V1 V52 9.155495474922957e-09
C1_52 V1 V52 -5.050452816685941e-21

R1_53 V1 V53 1401450.5401522422
L1_53 V1 V53 -3.086642045333136e-08
C1_53 V1 V53 -2.450533124392461e-21

R1_54 V1 V54 -1462423.9967887627
L1_54 V1 V54 1.6513956637089873e-08
C1_54 V1 V54 -2.493356092492769e-22

R1_55 V1 V55 -685697.3590686657
L1_55 V1 V55 6.379258191962469e-09
C1_55 V1 V55 -1.570150640364598e-21

R1_56 V1 V56 -890912.1133302493
L1_56 V1 V56 8.538688153465243e-09
C1_56 V1 V56 -8.534795472954785e-22

R1_57 V1 V57 -101369.67336762362
L1_57 V1 V57 1.0535652746819109e-09
C1_57 V1 V57 1.3012843427554375e-21

R1_58 V1 V58 -506574.6802424742
L1_58 V1 V58 5.312088089828148e-09
C1_58 V1 V58 8.217926709205395e-22

R1_59 V1 V59 218549487.70672575
L1_59 V1 V59 -1.2639234483926334e-07
C1_59 V1 V59 9.512041226937073e-22

R1_60 V1 V60 -856518.4811434228
L1_60 V1 V60 8.655046604078236e-09
C1_60 V1 V60 2.5010242193934017e-22

R1_61 V1 V61 414693.04993939324
L1_61 V1 V61 -5.1712957171823615e-09
C1_61 V1 V61 -3.658685693583345e-21

R1_62 V1 V62 589978.7212859753
L1_62 V1 V62 -7.843412808408912e-09
C1_62 V1 V62 -3.550019608678625e-21

R1_63 V1 V63 -861267.4288823472
L1_63 V1 V63 7.55514553883804e-09
C1_63 V1 V63 -5.642881149048322e-22

R1_64 V1 V64 2062206.2643365266
L1_64 V1 V64 -1.9816868834711433e-08
C1_64 V1 V64 1.4140884122887155e-23

R1_65 V1 V65 -902269.7054904008
L1_65 V1 V65 1.0457102773831963e-08
C1_65 V1 V65 -1.5240041896174158e-21

R1_66 V1 V66 1078982.856216841
L1_66 V1 V66 -9.055580185247047e-09
C1_66 V1 V66 -6.7995055671782055e-22

R1_67 V1 V67 -3006771.9473003964
L1_67 V1 V67 6.115335281011892e-08
C1_67 V1 V67 -5.973656651318281e-22

R1_68 V1 V68 -1687446.096172972
L1_68 V1 V68 1.4081775678361734e-08
C1_68 V1 V68 -3.0949848369106717e-22

R1_69 V1 V69 -9052349.336861283
L1_69 V1 V69 2.5314172433446704e-06
C1_69 V1 V69 3.165917547203309e-22

R1_70 V1 V70 -818520.4335827638
L1_70 V1 V70 6.683864525975626e-09
C1_70 V1 V70 7.059462057177734e-22

R1_71 V1 V71 -727767.347049306
L1_71 V1 V71 6.867361355868218e-09
C1_71 V1 V71 6.687809793114298e-23

R1_72 V1 V72 -593519.4213894722
L1_72 V1 V72 5.793284048969634e-09
C1_72 V1 V72 4.981342879926672e-22

R1_73 V1 V73 -726154.7589221237
L1_73 V1 V73 7.215288979736387e-09
C1_73 V1 V73 -6.125561186311525e-23

R1_74 V1 V74 -2891028.526898926
L1_74 V1 V74 3.3267259781992426e-08
C1_74 V1 V74 4.338769862454509e-22

R1_75 V1 V75 2369252.524528409
L1_75 V1 V75 -1.9330174211316795e-08
C1_75 V1 V75 -5.992295544599074e-22

R1_76 V1 V76 949902.041866384
L1_76 V1 V76 -1.0057739135561543e-08
C1_76 V1 V76 1.707278966582769e-23

R1_77 V1 V77 3058278.529729552
L1_77 V1 V77 -4.309076197662409e-08
C1_77 V1 V77 -3.5382253676290063e-22

R1_78 V1 V78 1391651.3671950893
L1_78 V1 V78 -1.567165311201621e-08
C1_78 V1 V78 2.507708236569878e-22

R1_79 V1 V79 -1655684.456960762
L1_79 V1 V79 1.5286493817785337e-08
C1_79 V1 V79 -3.777140496523959e-22

R1_80 V1 V80 -1111502.6385740878
L1_80 V1 V80 9.7023428262992e-09
C1_80 V1 V80 -1.4105691276472498e-21

R1_81 V1 V81 -3180537.602439113
L1_81 V1 V81 4.129913181684029e-08
C1_81 V1 V81 8.96438420813439e-22

R1_82 V1 V82 4213911.322560159
L1_82 V1 V82 -8.034706818088767e-06
C1_82 V1 V82 -2.0193786368205814e-21

R1_83 V1 V83 -1195074.881561418
L1_83 V1 V83 1.133582390558548e-08
C1_83 V1 V83 -2.28981729995327e-22

R1_84 V1 V84 -2896270.3600111636
L1_84 V1 V84 6.071922646930573e-08
C1_84 V1 V84 1.6721240742569983e-21

R1_85 V1 V85 -4716795.362988825
L1_85 V1 V85 5.418665279685167e-08
C1_85 V1 V85 1.6934387107601344e-21

R1_86 V1 V86 3167690.7094888883
L1_86 V1 V86 -2.9874305022998514e-08
C1_86 V1 V86 1.1182630068786639e-21

R1_87 V1 V87 1454800.7496338664
L1_87 V1 V87 -1.129250010763071e-08
C1_87 V1 V87 1.6670581475315065e-21

R1_88 V1 V88 1333408.6381786799
L1_88 V1 V88 -1.334097291378488e-08
C1_88 V1 V88 -2.8313435982336516e-23

R1_89 V1 V89 -696053.1793750672
L1_89 V1 V89 6.169279638160765e-09
C1_89 V1 V89 -3.2425813593640005e-21

R1_90 V1 V90 -3443754.016485305
L1_90 V1 V90 2.8145720762940472e-08
C1_90 V1 V90 -4.242550665491922e-22

R1_91 V1 V91 -2152448.2586292406
L1_91 V1 V91 1.5608222667900244e-08
C1_91 V1 V91 -1.162473247827108e-21

R1_92 V1 V92 -1852608.8580222558
L1_92 V1 V92 1.5439603264186715e-08
C1_92 V1 V92 -1.139471929984049e-21

R1_93 V1 V93 2622670.7309702113
L1_93 V1 V93 1.167617541131826e-07
C1_93 V1 V93 -6.049666961194877e-22

R1_94 V1 V94 947833.9629595152
L1_94 V1 V94 -9.962710811890822e-09
C1_94 V1 V94 9.041944996253866e-22

R1_95 V1 V95 21650079.26286582
L1_95 V1 V95 1.827924944083196e-07
C1_95 V1 V95 -7.254236547176128e-22

R1_96 V1 V96 -11250386.797580313
L1_96 V1 V96 1.5425672539357736e-07
C1_96 V1 V96 -4.986318144763171e-22

R1_97 V1 V97 -1402340.6600916826
L1_97 V1 V97 1.072116986403982e-08
C1_97 V1 V97 -7.69347883344696e-23

R1_98 V1 V98 -607064.5392113003
L1_98 V1 V98 4.912116968108495e-09
C1_98 V1 V98 -1.3283257644824645e-21

R1_99 V1 V99 4664032.150325526
L1_99 V1 V99 -1.0278665190570852e-07
C1_99 V1 V99 1.437698019898957e-22

R1_100 V1 V100 21297772.30512869
L1_100 V1 V100 -6.71781006306996e-08
C1_100 V1 V100 3.1535463917973907e-22

R1_101 V1 V101 -613243.5837422243
L1_101 V1 V101 4.726112685613836e-09
C1_101 V1 V101 -3.3370622884155835e-21

R1_102 V1 V102 -811769.7445107052
L1_102 V1 V102 6.486068208600473e-09
C1_102 V1 V102 -2.1390115279035516e-21

R1_103 V1 V103 -1711390.404223821
L1_103 V1 V103 1.5624298467135227e-08
C1_103 V1 V103 -2.288524898723252e-22

R1_104 V1 V104 13303391.39292363
L1_104 V1 V104 -1.7121809589362698e-07
C1_104 V1 V104 -1.6238603341875793e-22

R1_105 V1 V105 1520260.1600383609
L1_105 V1 V105 -1.0568155787918216e-08
C1_105 V1 V105 1.0432962631107801e-21

R1_106 V1 V106 -6599588.6049648635
L1_106 V1 V106 6.231455521736393e-08
C1_106 V1 V106 -1.8795116212243766e-21

R1_107 V1 V107 -5269078.610892548
L1_107 V1 V107 3.5397918120351514e-08
C1_107 V1 V107 -2.491964509463407e-22

R1_108 V1 V108 1633455.7452578458
L1_108 V1 V108 -1.1238941884644267e-08
C1_108 V1 V108 3.1541871644972083e-21

R1_109 V1 V109 -6673955.560010386
L1_109 V1 V109 6.702242041768541e-08
C1_109 V1 V109 9.183449763874366e-22

R1_110 V1 V110 970856.8964386502
L1_110 V1 V110 -7.797211126303572e-09
C1_110 V1 V110 2.259856238863837e-21

R1_111 V1 V111 -1113128.6186594053
L1_111 V1 V111 1.3303789514789824e-08
C1_111 V1 V111 5.0524221383538e-22

R1_112 V1 V112 -398598.83013509435
L1_112 V1 V112 3.723047592324976e-09
C1_112 V1 V112 -2.1901313226740027e-21

R1_113 V1 V113 -1015356.0691484276
L1_113 V1 V113 1.0446145129559443e-08
C1_113 V1 V113 -8.756084885912234e-22

R1_114 V1 V114 -1530102.9699661992
L1_114 V1 V114 1.1903460519159497e-08
C1_114 V1 V114 -1.2037175627443795e-21

R1_115 V1 V115 16583845.931724163
L1_115 V1 V115 1.484636220815114e-07
C1_115 V1 V115 1.4978296218055053e-22

R1_116 V1 V116 1718584.5393454952
L1_116 V1 V116 -1.3878659353327415e-08
C1_116 V1 V116 2.0187361819794865e-21

R1_117 V1 V117 1119947.6290512253
L1_117 V1 V117 -1.1745499879125276e-08
C1_117 V1 V117 1.519833338256691e-21

R1_118 V1 V118 1746102.0132761206
L1_118 V1 V118 -1.1982264603760076e-08
C1_118 V1 V118 1.0237488980688586e-21

R1_119 V1 V119 -3778825.3223985434
L1_119 V1 V119 -1.0547361060473124e-07
C1_119 V1 V119 1.3733410814643733e-21

R1_120 V1 V120 576205.9242385216
L1_120 V1 V120 -6.306052011868391e-09
C1_120 V1 V120 3.0675857383731888e-22

R1_121 V1 V121 -453234.43848173926
L1_121 V1 V121 4.833080869366125e-09
C1_121 V1 V121 3.4703757983399676e-23

R1_122 V1 V122 -424233.647523545
L1_122 V1 V122 4.5385512982356074e-09
C1_122 V1 V122 1.0990766150164231e-22

R1_123 V1 V123 -2518279.590135756
L1_123 V1 V123 2.1894502670419714e-08
C1_123 V1 V123 -4.0099855604402247e-23

R1_124 V1 V124 -2819604.889022666
L1_124 V1 V124 3.052444856266174e-08
C1_124 V1 V124 4.6104087512844755e-23

R1_125 V1 V125 327769.9214363838
L1_125 V1 V125 -3.5311878594038258e-09
C1_125 V1 V125 8.312698623966552e-22

R1_126 V1 V126 1418220.9132129846
L1_126 V1 V126 -1.7228862400004603e-08
C1_126 V1 V126 1.2670541911761877e-23

R1_127 V1 V127 8128955.869139963
L1_127 V1 V127 -1.3452295617387937e-07
C1_127 V1 V127 -7.001757841663426e-24

R1_128 V1 V128 6548344.088671126
L1_128 V1 V128 -1.530649027022328e-07
C1_128 V1 V128 -1.2443805642341043e-22

R1_129 V1 V129 -7165131.749022486
L1_129 V1 V129 4.619249992666612e-08
C1_129 V1 V129 2.1281113815397027e-22

R1_130 V1 V130 2378555.7728720475
L1_130 V1 V130 -2.27471190023386e-08
C1_130 V1 V130 6.457571498907343e-22

R1_131 V1 V131 2283956.394284192
L1_131 V1 V131 -2.6784855144760162e-08
C1_131 V1 V131 4.8786070674253297e-23

R1_132 V1 V132 5165008.448073854
L1_132 V1 V132 -4.813070936466818e-08
C1_132 V1 V132 -2.6941937826629985e-23

R1_133 V1 V133 2410285.2858179854
L1_133 V1 V133 -2.2158932964802693e-08
C1_133 V1 V133 -2.5793530182793574e-22

R1_134 V1 V134 1320410.4780889803
L1_134 V1 V134 -9.9042655812203e-09
C1_134 V1 V134 2.935599814283753e-23

R1_135 V1 V135 174890734.50693277
L1_135 V1 V135 -1.664592548413168e-07
C1_135 V1 V135 2.350638429623671e-23

R1_136 V1 V136 4341093.021484864
L1_136 V1 V136 -5.0295088708230144e-08
C1_136 V1 V136 1.1367551946295155e-22

R1_137 V1 V137 596636.1469189586
L1_137 V1 V137 -6.807862584734692e-09
C1_137 V1 V137 1.571250984869896e-22

R1_138 V1 V138 937873.6466902666
L1_138 V1 V138 -9.380584728931863e-09
C1_138 V1 V138 -6.566343755858544e-23

R1_139 V1 V139 3377950.4252117067
L1_139 V1 V139 -2.0091401667643498e-07
C1_139 V1 V139 5.633436971709963e-23

R1_140 V1 V140 1596978.721386951
L1_140 V1 V140 -1.2307054864814829e-08
C1_140 V1 V140 4.1511677071981066e-22

R1_141 V1 V141 2755203.2282374115
L1_141 V1 V141 -3.86355875506668e-08
C1_141 V1 V141 3.11672732564251e-23

R1_142 V1 V142 2137022.6892037555
L1_142 V1 V142 -1.440619467229633e-08
C1_142 V1 V142 3.3014390853137595e-22

R1_143 V1 V143 -2167665.0018736925
L1_143 V1 V143 2.4099626346447332e-08
C1_143 V1 V143 6.344356053853806e-23

R1_144 V1 V144 -1011138.082841155
L1_144 V1 V144 1.2801632896228117e-08
C1_144 V1 V144 -5.950854938297829e-23

R2_2 V2 0 -16598.25391868675
L2_2 V2 0 1.3663402264917693e-10
C2_2 V2 0 -7.044628079862263e-20

R2_3 V2 V3 -464134765.32059276
L2_3 V2 V3 -7.466204891194608e-06
C2_3 V2 V3 6.627145159301912e-24

R2_4 V2 V4 267277822.4601467
L2_4 V2 V4 -9.78586723435825e-05
C2_4 V2 V4 -4.396703962040296e-24

R2_5 V2 V5 8028283.501464993
L2_5 V2 V5 4.543290452198718e-08
C2_5 V2 V5 -9.670518095498818e-22

R2_6 V2 V6 -1544735.3219846075
L2_6 V2 V6 5.470304876717784e-08
C2_6 V2 V6 4.42562826843636e-22

R2_7 V2 V7 6685375.822887481
L2_7 V2 V7 -2.8804526280247934e-07
C2_7 V2 V7 2.0917583703109228e-23

R2_8 V2 V8 76569505.08801322
L2_8 V2 V8 2.7149033490131643e-07
C2_8 V2 V8 -2.4106317762941435e-23

R2_9 V2 V9 2710494.3409146806
L2_9 V2 V9 1.8412755271663976e-08
C2_9 V2 V9 1.5281860752041144e-21

R2_10 V2 V10 -5118422.0215715915
L2_10 V2 V10 -1.2635475698150586e-08
C2_10 V2 V10 2.302536394970034e-22

R2_11 V2 V11 2867969.430692642
L2_11 V2 V11 1.2955060765796995e-08
C2_11 V2 V11 5.894670676772178e-22

R2_12 V2 V12 100840170.83277157
L2_12 V2 V12 5.701871011004324e-08
C2_12 V2 V12 -1.5502535712615888e-22

R2_13 V2 V13 6327252.496050549
L2_13 V2 V13 -1.0170040861802575e-07
C2_13 V2 V13 -2.876502192749191e-22

R2_14 V2 V14 -6777595.074071171
L2_14 V2 V14 -1.0380310324886455e-07
C2_14 V2 V14 1.2330785998677858e-22

R2_15 V2 V15 2251298.058627233
L2_15 V2 V15 -2.5671929919517613e-08
C2_15 V2 V15 -3.6660193318370126e-23

R2_16 V2 V16 -7202337.1700584395
L2_16 V2 V16 -5.60243604808933e-07
C2_16 V2 V16 -1.3179183846945767e-22

R2_17 V2 V17 2288610.393013536
L2_17 V2 V17 -2.780586227976885e-06
C2_17 V2 V17 -3.1566574191405653e-22

R2_18 V2 V18 -2485025.3889011526
L2_18 V2 V18 1.0078616789007417e-07
C2_18 V2 V18 -5.501667212536036e-23

R2_19 V2 V19 3910983.6697651646
L2_19 V2 V19 2.4263334655761937e-08
C2_19 V2 V19 -7.8262714310386e-23

R2_20 V2 V20 -39825031.14205639
L2_20 V2 V20 -5.856889388436775e-07
C2_20 V2 V20 -5.771153578390855e-24

R2_21 V2 V21 4704586.611669512
L2_21 V2 V21 3.634873959364357e-09
C2_21 V2 V21 8.058147179955419e-22

R2_22 V2 V22 -6480406.288501584
L2_22 V2 V22 -2.703871106860538e-09
C2_22 V2 V22 -7.581651425668904e-22

R2_23 V2 V23 -26434514.78845729
L2_23 V2 V23 4.471818625214553e-08
C2_23 V2 V23 -1.7341799865347526e-22

R2_24 V2 V24 -47566988.92132696
L2_24 V2 V24 4.130321793504151e-08
C2_24 V2 V24 -1.1407104137514046e-23

R2_25 V2 V25 3564830.666791173
L2_25 V2 V25 7.403573752816353e-09
C2_25 V2 V25 3.9999934483241542e-22

R2_26 V2 V26 -2972710.504762462
L2_26 V2 V26 -6.041342408524807e-09
C2_26 V2 V26 4.5384871381096e-23

R2_27 V2 V27 -13287617.712034905
L2_27 V2 V27 -3.3806564515322894e-08
C2_27 V2 V27 1.3449829035053727e-22

R2_28 V2 V28 -17023260.090950422
L2_28 V2 V28 -6.319677872373745e-08
C2_28 V2 V28 1.2392733180484079e-23

R2_29 V2 V29 -2249706.700506102
L2_29 V2 V29 4.3244590644072375e-09
C2_29 V2 V29 -2.9427958561612753e-21

R2_30 V2 V30 1233170.4111738794
L2_30 V2 V30 -4.066027482985572e-09
C2_30 V2 V30 2.5782879850381134e-22

R2_31 V2 V31 -14127195.687006332
L2_31 V2 V31 3.511163990359686e-08
C2_31 V2 V31 -9.317232461676088e-22

R2_32 V2 V32 -10646309.146970887
L2_32 V2 V32 3.939928465659243e-08
C2_32 V2 V32 -4.72914652924051e-22

R2_33 V2 V33 432027.7008673561
L2_33 V2 V33 -3.4787250811867813e-09
C2_33 V2 V33 3.641210790073506e-21

R2_34 V2 V34 -816318.474436411
L2_34 V2 V34 7.899618512580589e-09
C2_34 V2 V34 -1.5167958147867585e-21

R2_35 V2 V35 729387.9383414787
L2_35 V2 V35 -6.772531286588097e-09
C2_35 V2 V35 2.3951697290631125e-21

R2_36 V2 V36 -3328622.0332434173
L2_36 V2 V36 2.7905405333079584e-08
C2_36 V2 V36 -3.3169113553500066e-22

R2_37 V2 V37 -178663.0555793493
L2_37 V2 V37 1.458303821202749e-09
C2_37 V2 V37 -7.683483658593131e-21

R2_38 V2 V38 1587916.1815414936
L2_38 V2 V38 -7.642515927110843e-09
C2_38 V2 V38 1.5710121586914955e-21

R2_39 V2 V39 -221317.67168855786
L2_39 V2 V39 1.9652285513616747e-09
C2_39 V2 V39 -6.837905308735239e-21

R2_40 V2 V40 -3001746.4960525557
L2_40 V2 V40 1.8842513379704014e-08
C2_40 V2 V40 -4.941254565619937e-22

R2_41 V2 V41 49247.911961832004
L2_41 V2 V41 -4.4607928998383965e-10
C2_41 V2 V41 2.617055264637077e-20

R2_42 V2 V42 122694.11065692459
L2_42 V2 V42 -1.0353932664703243e-09
C2_42 V2 V42 9.951066634132869e-21

R2_43 V2 V43 127309.29923690995
L2_43 V2 V43 -1.1869877186078185e-09
C2_43 V2 V43 9.086756462852295e-21

R2_44 V2 V44 1703004.2519272552
L2_44 V2 V44 -1.4992431360822584e-08
C2_44 V2 V44 7.515250640227825e-22

R2_45 V2 V45 -176984.35014046598
L2_45 V2 V45 1.4178180117467436e-09
C2_45 V2 V45 -1.4337390904336163e-20

R2_46 V2 V46 1875053.9125895968
L2_46 V2 V46 -3.1710976907471624e-08
C2_46 V2 V46 -4.787270281385801e-21

R2_47 V2 V47 560710.2876326484
L2_47 V2 V47 -8.300297367826769e-09
C2_47 V2 V47 -1.3986926047105152e-21

R2_48 V2 V48 -2563629.1982271564
L2_48 V2 V48 1.914099989521306e-08
C2_48 V2 V48 -7.611719792772675e-23

R2_49 V2 V49 -846037.1180080662
L2_49 V2 V49 1.4292022172930286e-08
C2_49 V2 V49 4.728305324557671e-21

R2_50 V2 V50 471379.15730621567
L2_50 V2 V50 -4.615861451706547e-09
C2_50 V2 V50 2.7528600661129823e-21

R2_51 V2 V51 -300452.9568473322
L2_51 V2 V51 3.0323837681859175e-09
C2_51 V2 V51 -5.110969824578016e-22

R2_52 V2 V52 1400965.083674924
L2_52 V2 V52 -5.9601871220779164e-09
C2_52 V2 V52 9.835570064944916e-21

R2_53 V2 V53 2554631.3675525137
L2_53 V2 V53 -6.9021947016569995e-09
C2_53 V2 V53 8.643206251252378e-21

R2_54 V2 V54 865314.846285405
L2_54 V2 V54 -9.42256440579449e-09
C2_54 V2 V54 6.880268654585119e-22

R2_55 V2 V55 321664.3876069898
L2_55 V2 V55 -3.136056222330645e-09
C2_55 V2 V55 3.8452958382005874e-21

R2_56 V2 V56 327554.58315089374
L2_56 V2 V56 -2.9070545658741804e-09
C2_56 V2 V56 5.5003259336860595e-21

R2_57 V2 V57 49216.089046359804
L2_57 V2 V57 -5.131527616426603e-10
C2_57 V2 V57 -4.033912573610479e-21

R2_58 V2 V58 -827506.4776425986
L2_58 V2 V58 9.809594148151674e-09
C2_58 V2 V58 -3.5126096734057167e-22

R2_59 V2 V59 27796300.28888489
L2_59 V2 V59 3.653068393799374e-07
C2_59 V2 V59 -1.0293399464634224e-21

R2_60 V2 V60 300974.7463030751
L2_60 V2 V60 -3.0451431746869348e-09
C2_60 V2 V60 1.2270922882570377e-22

R2_61 V2 V61 -250164.55193084048
L2_61 V2 V61 3.903593080377951e-09
C2_61 V2 V61 1.0839784614991505e-20

R2_62 V2 V62 -311720.0541977106
L2_62 V2 V62 3.422959649097056e-09
C2_62 V2 V62 5.444558979968133e-21

R2_63 V2 V63 2636594.611546251
L2_63 V2 V63 -8.22070644053174e-09
C2_63 V2 V63 4.84501807547823e-21

R2_64 V2 V64 5671480.143446064
L2_64 V2 V64 -1.6381241997721204e-08
C2_64 V2 V64 3.8459458341606476e-21

R2_65 V2 V65 453114.14460881427
L2_65 V2 V65 -6.0611241631994355e-09
C2_65 V2 V65 2.5663627580293354e-21

R2_66 V2 V66 1255717.8386187893
L2_66 V2 V66 -9.085447378152784e-09
C2_66 V2 V66 4.725373041763146e-21

R2_67 V2 V67 -3403580.044240243
L2_67 V2 V67 9.366523973743265e-09
C2_67 V2 V67 8.31335266521186e-22

R2_68 V2 V68 1273954.2319084578
L2_68 V2 V68 -1.2988282408587683e-08
C2_68 V2 V68 4.938624386266307e-22

R2_69 V2 V69 8234214.678762466
L2_69 V2 V69 4.239728377153699e-08
C2_69 V2 V69 -1.4017200382807775e-22

R2_70 V2 V70 205968.96984990197
L2_70 V2 V70 -1.7589386423816162e-09
C2_70 V2 V70 4.163192380472793e-21

R2_71 V2 V71 128931.06884812684
L2_71 V2 V71 -1.1001238236469469e-09
C2_71 V2 V71 2.4865537491844655e-21

R2_72 V2 V72 476291.5462123885
L2_72 V2 V72 -5.176955511013495e-09
C2_72 V2 V72 -2.084248296899213e-22

R2_73 V2 V73 1022510.2570774391
L2_73 V2 V73 -9.617231588873826e-09
C2_73 V2 V73 3.75135559956275e-22

R2_74 V2 V74 990966.6970881205
L2_74 V2 V74 -8.300754061417645e-09
C2_74 V2 V74 1.1254457563304014e-21

R2_75 V2 V75 -478218.84398592287
L2_75 V2 V75 3.941761547504857e-09
C2_75 V2 V75 -2.1959845382717093e-21

R2_76 V2 V76 1122307.0544384886
L2_76 V2 V76 -5.688907768032162e-09
C2_76 V2 V76 6.3213367191721406e-21

R2_77 V2 V77 -10114124.502744783
L2_77 V2 V77 -2.7113059978931933e-08
C2_77 V2 V77 1.261043557598604e-21

R2_78 V2 V78 -3431177.9949026573
L2_78 V2 V78 -6.637408600142379e-08
C2_78 V2 V78 1.83768661068434e-21

R2_79 V2 V79 211093.6175813218
L2_79 V2 V79 -1.7716764738579702e-09
C2_79 V2 V79 9.484642945043628e-21

R2_80 V2 V80 -829907.5871838259
L2_80 V2 V80 7.725142024649827e-09
C2_80 V2 V80 -4.393678989714966e-21

R2_81 V2 V81 4833460.610357505
L2_81 V2 V81 -1.3959317263957953e-07
C2_81 V2 V81 -2.25401000589874e-21

R2_82 V2 V82 -378696.6270379321
L2_82 V2 V82 3.827650418532891e-09
C2_82 V2 V82 -1.618082008449578e-21

R2_83 V2 V83 14153934.345235303
L2_83 V2 V83 3.952698144026955e-08
C2_83 V2 V83 -5.7915287219281905e-21

R2_84 V2 V84 639120.2241219201
L2_84 V2 V84 -5.671901740138614e-09
C2_84 V2 V84 -4.345643215068273e-22

R2_85 V2 V85 380837.47446557845
L2_85 V2 V85 -3.055224942526626e-09
C2_85 V2 V85 3.0965926488334e-21

R2_86 V2 V86 -1767751.7340569
L2_86 V2 V86 1.34708347899092e-08
C2_86 V2 V86 -6.332337725368667e-22

R2_87 V2 V87 774153.5221306864
L2_87 V2 V87 -6.242667113050841e-09
C2_87 V2 V87 3.0563485666923476e-21

R2_88 V2 V88 -770886.0058899634
L2_88 V2 V88 6.984594501082451e-09
C2_88 V2 V88 4.364633550570707e-22

R2_89 V2 V89 389226.2360312805
L2_89 V2 V89 -3.5958768756603396e-09
C2_89 V2 V89 5.236711915808688e-21

R2_90 V2 V90 -288825.6917293818
L2_90 V2 V90 2.444910317211345e-09
C2_90 V2 V90 -6.996400956051701e-21

R2_91 V2 V91 -1099940.8942624545
L2_91 V2 V91 9.858527557154378e-09
C2_91 V2 V91 -1.2481756600327752e-21

R2_92 V2 V92 -5707805.203888551
L2_92 V2 V92 4.342241400794157e-08
C2_92 V2 V92 -8.387829832125654e-22

R2_93 V2 V93 2542132.6925973925
L2_93 V2 V93 -5.608766191563338e-09
C2_93 V2 V93 3.0349529353053125e-21

R2_94 V2 V94 -417238.27253422834
L2_94 V2 V94 4.210063027313488e-09
C2_94 V2 V94 -3.579185448698709e-21

R2_95 V2 V95 -711064.8500121612
L2_95 V2 V95 8.815387726630637e-09
C2_95 V2 V95 -1.525024733223549e-21

R2_96 V2 V96 -1278672.9531197501
L2_96 V2 V96 9.417478323931764e-09
C2_96 V2 V96 -1.5205162086537526e-21

R2_97 V2 V97 -1532216.1500385501
L2_97 V2 V97 1.2276552501471952e-08
C2_97 V2 V97 -2.8660256036305096e-21

R2_98 V2 V98 932136.0973392973
L2_98 V2 V98 -6.388878449839909e-09
C2_98 V2 V98 -2.1421599407796152e-21

R2_99 V2 V99 662271.595891302
L2_99 V2 V99 -4.576820161611853e-09
C2_99 V2 V99 1.3154583926917702e-21

R2_100 V2 V100 -3620074.734076392
L2_100 V2 V100 1.975604087122046e-08
C2_100 V2 V100 -7.187828008930672e-22

R2_101 V2 V101 385761.95747226477
L2_101 V2 V101 -3.191012291257192e-09
C2_101 V2 V101 3.684681868615182e-21

R2_102 V2 V102 -177330.24208946736
L2_102 V2 V102 1.5119123762088744e-09
C2_102 V2 V102 -1.5391083873859462e-20

R2_103 V2 V103 168587.25582617847
L2_103 V2 V103 -1.4726151192194105e-09
C2_103 V2 V103 1.2271382980792967e-20

R2_104 V2 V104 -32212211.807844173
L2_104 V2 V104 -9.540464479096833e-08
C2_104 V2 V104 3.0810693003202216e-22

R2_105 V2 V105 562622.9979444204
L2_105 V2 V105 -4.2980062352447665e-09
C2_105 V2 V105 5.2127435600287886e-21

R2_106 V2 V106 -231841.91554622815
L2_106 V2 V106 1.7458510491860731e-09
C2_106 V2 V106 -9.888173199460563e-21

R2_107 V2 V107 -179511.77746392312
L2_107 V2 V107 1.4058888078893292e-09
C2_107 V2 V107 -1.6962359107668757e-20

R2_108 V2 V108 301832.6461818642
L2_108 V2 V108 -2.112912716416447e-09
C2_108 V2 V108 7.038383773370728e-21

R2_109 V2 V109 355794.53949414956
L2_109 V2 V109 -2.848124242960218e-09
C2_109 V2 V109 4.964027886445002e-21

R2_110 V2 V110 -3464268.0376774133
L2_110 V2 V110 -2.747538929848018e-08
C2_110 V2 V110 3.4826823836330744e-21

R2_111 V2 V111 164250.8831963773
L2_111 V2 V111 -1.5731125505404492e-09
C2_111 V2 V111 8.214641532932116e-21

R2_112 V2 V112 -3045071.3614095068
L2_112 V2 V112 1.2050323761342258e-08
C2_112 V2 V112 -7.494184435857428e-21

R2_113 V2 V113 -1251155.8233431967
L2_113 V2 V113 9.315984692268823e-09
C2_113 V2 V113 -3.385975606833796e-21

R2_114 V2 V114 -856366.6128045991
L2_114 V2 V114 7.1040991248203455e-09
C2_114 V2 V114 -3.1674948866083203e-21

R2_115 V2 V115 -254934.3942535894
L2_115 V2 V115 2.589382646373891e-09
C2_115 V2 V115 -9.291883709235086e-21

R2_116 V2 V116 444973.4714868123
L2_116 V2 V116 -3.767002493812145e-09
C2_116 V2 V116 2.2043191568278886e-21

R2_117 V2 V117 -2814700.6096163853
L2_117 V2 V117 -4.185469215611147e-08
C2_117 V2 V117 3.388370866596649e-21

R2_118 V2 V118 729895.2549750117
L2_118 V2 V118 -6.9918186895843e-09
C2_118 V2 V118 2.585846186384332e-21

R2_119 V2 V119 265686.70720891684
L2_119 V2 V119 -2.7810211030035146e-09
C2_119 V2 V119 3.0567824825918253e-21

R2_120 V2 V120 -146513.7984994706
L2_120 V2 V120 1.6000793253187093e-09
C2_120 V2 V120 2.0467812714043383e-21

R2_121 V2 V121 264482.76033595146
L2_121 V2 V121 -3.0050895634151927e-09
C2_121 V2 V121 -1.6779652945761484e-21

R2_122 V2 V122 -788222.2012149282
L2_122 V2 V122 9.24193441955356e-09
C2_122 V2 V122 -7.101870329761073e-23

R2_123 V2 V123 -5662996.871146351
L2_123 V2 V123 9.640838853490311e-08
C2_123 V2 V123 9.922093548054283e-22

R2_124 V2 V124 620952.9997885637
L2_124 V2 V124 -5.791747841038982e-09
C2_124 V2 V124 1.0194014390911567e-21

R2_125 V2 V125 -146557.12619480497
L2_125 V2 V125 1.6595990064572327e-09
C2_125 V2 V125 -4.371275666678909e-22

R2_126 V2 V126 163676.89762727742
L2_126 V2 V126 -1.679394609950197e-09
C2_126 V2 V126 -1.6731475742395204e-21

R2_127 V2 V127 -156591.70670206586
L2_127 V2 V127 1.6418838389995597e-09
C2_127 V2 V127 -4.711570909985393e-22

R2_128 V2 V128 -1442126.8335706994
L2_128 V2 V128 1.8329562229095607e-08
C2_128 V2 V128 3.8830458788482714e-22

R2_129 V2 V129 -597310.5886082778
L2_129 V2 V129 6.976680446257762e-09
C2_129 V2 V129 -5.320522157666889e-22

R2_130 V2 V130 438796.3384612707
L2_130 V2 V130 -3.5025493709153994e-09
C2_130 V2 V130 3.185449204178414e-21

R2_131 V2 V131 12672879.619198516
L2_131 V2 V131 4.613007877909802e-08
C2_131 V2 V131 -4.777924834510119e-21

R2_132 V2 V132 783600.932023793
L2_132 V2 V132 -8.698437272476713e-09
C2_132 V2 V132 7.595286261282403e-23

R2_133 V2 V133 -549087.6298692769
L2_133 V2 V133 4.333239397375927e-09
C2_133 V2 V133 -2.843476007563872e-21

R2_134 V2 V134 -1730904.9303851097
L2_134 V2 V134 8.192784458480933e-09
C2_134 V2 V134 -6.598472092335081e-22

R2_135 V2 V135 -260791.95014478866
L2_135 V2 V135 2.5700606499259002e-09
C2_135 V2 V135 1.885468764016298e-21

R2_136 V2 V136 -1884444.8865981698
L2_136 V2 V136 2.1500653024480288e-08
C2_136 V2 V136 -1.426966751824732e-22

R2_137 V2 V137 -357480.7182527387
L2_137 V2 V137 4.858850612251273e-09
C2_137 V2 V137 1.4870162311944885e-21

R2_138 V2 V138 201317.10451913046
L2_138 V2 V138 -2.225484035061966e-09
C2_138 V2 V138 1.0416458921646887e-21

R2_139 V2 V139 -113141.81986529748
L2_139 V2 V139 1.254127848007131e-09
C2_139 V2 V139 -2.6546429234812566e-21

R2_140 V2 V140 886144.2434393744
L2_140 V2 V140 -8.041299693404997e-09
C2_140 V2 V140 8.689395121881005e-22

R2_141 V2 V141 1246471.2272817874
L2_141 V2 V141 -9.868186808966014e-09
C2_141 V2 V141 8.267536454015628e-22

R2_142 V2 V142 555900.4061520792
L2_142 V2 V142 -5.530922786317309e-09
C2_142 V2 V142 1.3892570909529958e-21

R2_143 V2 V143 278054.6255032842
L2_143 V2 V143 -2.892840451059142e-09
C2_143 V2 V143 -9.187927543732806e-22

R2_144 V2 V144 1908074.8441534229
L2_144 V2 V144 2.5888774497486817e-08
C2_144 V2 V144 2.0831310022760955e-22

R3_3 V3 0 -15844.578596616017
L3_3 V3 0 1.8272355419274677e-10
C3_3 V3 0 -2.9041228806181295e-20

R3_4 V3 V4 -200483705.4429442
L3_4 V3 V4 5.142119067086406e-06
C3_4 V3 V4 8.461394404944589e-23

R3_5 V3 V5 -7582035.937310421
L3_5 V3 V5 1.9769608986934794e-08
C3_5 V3 V5 -9.476079275745161e-22

R3_6 V3 V6 4342408.933865775
L3_6 V3 V6 9.63430492762005e-08
C3_6 V3 V6 -1.7058220852370324e-22

R3_7 V3 V7 -3818873.891842494
L3_7 V3 V7 8.4114925539224e-08
C3_7 V3 V7 2.382932193931356e-22

R3_8 V3 V8 -7187423.421906916
L3_8 V3 V8 3.931429368616709e-08
C3_8 V3 V8 -2.3056822287020202e-23

R3_9 V3 V9 1551110.8722753595
L3_9 V3 V9 2.3076536525274465e-08
C3_9 V3 V9 1.3024437641259908e-21

R3_10 V3 V10 9286339.852465441
L3_10 V3 V10 1.4205291528762048e-08
C3_10 V3 V10 1.8152640950080765e-22

R3_11 V3 V11 -114007061.30466205
L3_11 V3 V11 -2.350904455054028e-08
C3_11 V3 V11 6.761412238343776e-22

R3_12 V3 V12 -5255594.764994696
L3_12 V3 V12 1.214541027501861e-06
C3_12 V3 V12 -9.913232597739978e-23

R3_13 V3 V13 18964149.0046642
L3_13 V3 V13 4.371319920272657e-08
C3_13 V3 V13 -1.0272620133126183e-22

R3_14 V3 V14 5398147.698580737
L3_14 V3 V14 3.5547961897542845e-08
C3_14 V3 V14 1.0441744692681459e-22

R3_15 V3 V15 -4075408.290191935
L3_15 V3 V15 6.192489353649147e-08
C3_15 V3 V15 -3.570900656593216e-22

R3_16 V3 V16 35646793.89240865
L3_16 V3 V16 7.460792207805531e-08
C3_16 V3 V16 -8.659756184447211e-24

R3_17 V3 V17 4805995.670747269
L3_17 V3 V17 1.2502134114550082e-08
C3_17 V3 V17 -2.2380751083394938e-22

R3_18 V3 V18 5522033.552749715
L3_18 V3 V18 4.077530574634185e-08
C3_18 V3 V18 3.4498384618440172e-22

R3_19 V3 V19 -1577206.0028308171
L3_19 V3 V19 9.429771705416101e-09
C3_19 V3 V19 2.0457333707979247e-22

R3_20 V3 V20 -8623830.040035319
L3_20 V3 V20 -6.73890994567272e-07
C3_20 V3 V20 1.412165063930602e-23

R3_21 V3 V21 3345084.6969309254
L3_21 V3 V21 3.6214172272515943e-09
C3_21 V3 V21 7.69877105885032e-22

R3_22 V3 V22 -141061057.25780606
L3_22 V3 V22 4.430145439261143e-09
C3_22 V3 V22 3.1973773666167925e-22

R3_23 V3 V23 -7685888.5479354495
L3_23 V3 V23 -6.108962053537348e-09
C3_23 V3 V23 -4.401632183266665e-22

R3_24 V3 V24 12859126.741803357
L3_24 V3 V24 -1.4838441314602158e-08
C3_24 V3 V24 -1.0322491283374585e-22

R3_25 V3 V25 12702590.621892905
L3_25 V3 V25 8.462013452339146e-09
C3_25 V3 V25 1.8336902494041383e-22

R3_26 V3 V26 11804690.532153485
L3_26 V3 V26 7.535982079855664e-09
C3_26 V3 V26 -5.43784384871403e-23

R3_27 V3 V27 -23070219.47380599
L3_27 V3 V27 8.2941672225689e-08
C3_27 V3 V27 -1.568480450646483e-22

R3_28 V3 V28 -4659637.4044531
L3_28 V3 V28 2.679178458106228e-08
C3_28 V3 V28 -2.369848805813675e-22

R3_29 V3 V29 -2458511.7943269736
L3_29 V3 V29 5.044714302155815e-09
C3_29 V3 V29 -2.6468593568645882e-21

R3_30 V3 V30 -1418928.603132689
L3_30 V3 V30 5.630180888569598e-09
C3_30 V3 V30 -1.1022348204086299e-21

R3_31 V3 V31 -3242714.2962993006
L3_31 V3 V31 -1.3266677729285923e-08
C3_31 V3 V31 -2.2651463609693973e-22

R3_32 V3 V32 6360991.425298552
L3_32 V3 V32 -2.331797726253502e-08
C3_32 V3 V32 -2.8498962119338046e-22

R3_33 V3 V33 682746.2993852535
L3_33 V3 V33 -5.900258076337688e-09
C3_33 V3 V33 3.8738735723781894e-21

R3_34 V3 V34 -5909084.8823316125
L3_34 V3 V34 3.300347069014078e-08
C3_34 V3 V34 -1.0558768147355163e-21

R3_35 V3 V35 6858702.211873575
L3_35 V3 V35 -4.412633178427557e-08
C3_35 V3 V35 1.6683963349956909e-21

R3_36 V3 V36 -3169781.583271021
L3_36 V3 V36 2.122409208650935e-08
C3_36 V3 V36 -3.1695103878080993e-22

R3_37 V3 V37 -222983.9322918328
L3_37 V3 V37 1.809722098492942e-09
C3_37 V3 V37 -6.711334811566126e-21

R3_38 V3 V38 -660817.9300510808
L3_38 V3 V38 5.064060940147954e-09
C3_38 V3 V38 -1.6115405853439721e-21

R3_39 V3 V39 -229109.21134269456
L3_39 V3 V39 2.047620878858421e-09
C3_39 V3 V39 -5.954327270281073e-21

R3_40 V3 V40 -2122199.5277558817
L3_40 V3 V40 2.4483335507824276e-08
C3_40 V3 V40 -4.464050483746243e-22

R3_41 V3 V41 58822.46120692364
L3_41 V3 V41 -5.325833919285517e-10
C3_41 V3 V41 1.8705808099130436e-20

R3_42 V3 V42 60596.34477571149
L3_42 V3 V42 -5.33303669782374e-10
C3_42 V3 V42 2.277599993970785e-20

R3_43 V3 V43 232412.39582545086
L3_43 V3 V43 -1.7868148937735473e-09
C3_43 V3 V43 7.861235489485647e-21

R3_44 V3 V44 3166570.568100301
L3_44 V3 V44 -1.4619755682452954e-08
C3_44 V3 V44 2.4793918862780974e-21

R3_45 V3 V45 -204682.48815876464
L3_45 V3 V45 1.6140256431217932e-09
C3_45 V3 V45 -1.3688711125618173e-20

R3_46 V3 V46 -509510.0187093949
L3_46 V3 V46 3.863052717747449e-09
C3_46 V3 V46 -8.817292920882915e-21

R3_47 V3 V47 -10006727.737695472
L3_47 V3 V47 6.201871123925824e-08
C3_47 V3 V47 -4.023592215640593e-21

R3_48 V3 V48 -613808.8759834982
L3_48 V3 V48 5.5382851423399754e-09
C3_48 V3 V48 -2.351265515921468e-21

R3_49 V3 V49 -954287.0929767417
L3_49 V3 V49 1.2955216876450369e-08
C3_49 V3 V49 3.1363719801850418e-21

R3_50 V3 V50 795505.7748622794
L3_50 V3 V50 -5.279892201368324e-09
C3_50 V3 V50 4.97345577066646e-21

R3_51 V3 V51 -419184.963115637
L3_51 V3 V51 3.4675397693532136e-09
C3_51 V3 V51 -5.052915278747638e-21

R3_52 V3 V52 647127.4866938329
L3_52 V3 V52 -3.661773685884028e-09
C3_52 V3 V52 1.0728375476132046e-20

R3_53 V3 V53 -355883.84398830566
L3_53 V3 V53 4.706740296686624e-09
C3_53 V3 V53 2.506396597671162e-21

R3_54 V3 V54 669458.5591572055
L3_54 V3 V54 -7.2302013721335025e-09
C3_54 V3 V54 4.610418074519529e-22

R3_55 V3 V55 381437.28658959264
L3_55 V3 V55 -3.624313657945465e-09
C3_55 V3 V55 2.3291503248913716e-21

R3_56 V3 V56 622751.802327546
L3_56 V3 V56 -6.626157544030783e-09
C3_56 V3 V56 -1.0564648555475644e-21

R3_57 V3 V57 49482.63587540879
L3_57 V3 V57 -5.131045768990788e-10
C3_57 V3 V57 -1.7860327283771947e-21

R3_58 V3 V58 117414.88583564766
L3_58 V3 V58 -1.2353755734093221e-09
C3_58 V3 V58 -2.7205382920638094e-21

R3_59 V3 V59 -1585505.6477547626
L3_59 V3 V59 1.2596115923628796e-08
C3_59 V3 V59 -2.6550498455103774e-21

R3_60 V3 V60 564085.9573883748
L3_60 V3 V60 -5.825475733188812e-09
C3_60 V3 V60 -1.0095966146534556e-21

R3_61 V3 V61 -177233.23540710617
L3_61 V3 V61 1.993538839241726e-09
C3_61 V3 V61 5.218286404632372e-21

R3_62 V3 V62 -257390.1492615146
L3_62 V3 V62 3.961079398945447e-09
C3_62 V3 V62 8.704726525497408e-21

R3_63 V3 V63 257381.48283410768
L3_63 V3 V63 -2.5910333815441357e-09
C3_63 V3 V63 -2.064504135026238e-21

R3_64 V3 V64 -492342.950709017
L3_64 V3 V64 4.139188477828989e-09
C3_64 V3 V64 -2.8281306079720886e-21

R3_65 V3 V65 473557.64175882045
L3_65 V3 V65 -5.289539673603881e-09
C3_65 V3 V65 3.467463943719827e-21

R3_66 V3 V66 -306851.5569343401
L3_66 V3 V66 2.5049665775936397e-09
C3_66 V3 V66 -6.416054297562593e-22

R3_67 V3 V67 747766.9083950398
L3_67 V3 V67 -7.32703789039527e-09
C3_67 V3 V67 1.5575825201528048e-21

R3_68 V3 V68 600972.0305884632
L3_68 V3 V68 -4.806566343933524e-09
C3_68 V3 V68 2.844289950368463e-22

R3_69 V3 V69 1509893.7252553974
L3_69 V3 V69 -1.9311987023945347e-08
C3_69 V3 V69 -1.7246240274459697e-21

R3_70 V3 V70 1481717.0541831988
L3_70 V3 V70 -8.470102144879354e-09
C3_70 V3 V70 -4.6053892657329955e-21

R3_71 V3 V71 -960542.4885453265
L3_71 V3 V71 5.454321908812186e-09
C3_71 V3 V71 -2.2444534706295167e-21

R3_72 V3 V72 225961.77085152728
L3_72 V3 V72 -2.0276866491312885e-09
C3_72 V3 V72 -8.807102186155217e-22

R3_73 V3 V73 233300.05312961419
L3_73 V3 V73 -2.3546813921493124e-09
C3_73 V3 V73 -5.2649056177819156e-24

R3_74 V3 V74 2054853.547427481
L3_74 V3 V74 -1.7887879452089537e-07
C3_74 V3 V74 -3.072739975353162e-21

R3_75 V3 V75 8833638.417067504
L3_75 V3 V75 -2.9871114093662956e-07
C3_75 V3 V75 3.354951527247266e-21

R3_76 V3 V76 -224403.98574060362
L3_76 V3 V76 2.0525804091918767e-09
C3_76 V3 V76 -4.701820441733388e-21

R3_77 V3 V77 -965460.673339475
L3_77 V3 V77 9.139882063955042e-09
C3_77 V3 V77 3.043571290884243e-22

R3_78 V3 V78 -553483.4003650178
L3_78 V3 V78 5.712984713434503e-09
C3_78 V3 V78 -1.167250473149415e-21

R3_79 V3 V79 -670553.5422991186
L3_79 V3 V79 4.8726173563284136e-09
C3_79 V3 V79 -6.0666384631342475e-21

R3_80 V3 V80 230362.02445414977
L3_80 V3 V80 -2.0374931345141213e-09
C3_80 V3 V80 8.820268369171336e-21

R3_81 V3 V81 1207412.9028195292
L3_81 V3 V81 -1.523000077240393e-08
C3_81 V3 V81 -1.862336961261238e-21

R3_82 V3 V82 -3615855.9905302864
L3_82 V3 V82 -1.0258619215269268e-07
C3_82 V3 V82 4.4921586829671e-21

R3_83 V3 V83 492998.0049153543
L3_83 V3 V83 -4.618521401002722e-09
C3_83 V3 V83 2.602098828759712e-21

R3_84 V3 V84 -6696857.8311371105
L3_84 V3 V84 1.0764242470934646e-08
C3_84 V3 V84 -6.082089997775556e-21

R3_85 V3 V85 -938535.4901864799
L3_85 V3 V85 6.468163295801516e-09
C3_85 V3 V85 -7.847649701232085e-21

R3_86 V3 V86 -7090865.964732199
L3_86 V3 V86 -8.479412448559819e-08
C3_86 V3 V86 -1.579665395490337e-21

R3_87 V3 V87 -344758.47022236325
L3_87 V3 V87 2.6789831416025066e-09
C3_87 V3 V87 -6.197829820701138e-21

R3_88 V3 V88 -678743.110482549
L3_88 V3 V88 7.66612413348408e-09
C3_88 V3 V88 5.375105210099361e-22

R3_89 V3 V89 330731.03917372506
L3_89 V3 V89 -2.891859031049181e-09
C3_89 V3 V89 6.914604667519138e-21

R3_90 V3 V90 255265.19241387805
L3_90 V3 V90 -2.1471418882779423e-09
C3_90 V3 V90 7.55170031581837e-21

R3_91 V3 V91 1219918.4125613861
L3_91 V3 V91 -8.773945391836897e-09
C3_91 V3 V91 5.743406147250252e-22

R3_92 V3 V92 552483.9070724268
L3_92 V3 V92 -4.802203930528666e-09
C3_92 V3 V92 3.758474522182303e-21

R3_93 V3 V93 -663666.6112175363
L3_93 V3 V93 1.2384227320361147e-08
C3_93 V3 V93 2.0810570645627476e-22

R3_94 V3 V94 -668355.8178083878
L3_94 V3 V94 8.253898239850011e-09
C3_94 V3 V94 7.214835166542978e-22

R3_95 V3 V95 10167795.12258905
L3_95 V3 V95 -1.9211040361153595e-07
C3_95 V3 V95 1.591492116337809e-21

R3_96 V3 V96 960568.1426958954
L3_96 V3 V96 -7.57476480085614e-09
C3_96 V3 V96 2.949697994230911e-21

R3_97 V3 V97 274564.19231491064
L3_97 V3 V97 -2.0908117489051866e-09
C3_97 V3 V97 3.721273285993408e-21

R3_98 V3 V98 212698.12504622448
L3_98 V3 V98 -1.7831051166960517e-09
C3_98 V3 V98 5.074000599027945e-21

R3_99 V3 V99 -519885.54840081546
L3_99 V3 V99 4.860298760166138e-09
C3_99 V3 V99 -1.4080164076751723e-21

R3_100 V3 V100 12690456.21937371
L3_100 V3 V100 5.835880089524926e-07
C3_100 V3 V100 -4.786498224035493e-22

R3_101 V3 V101 288488.13647011964
L3_101 V3 V101 -2.1353116750131342e-09
C3_101 V3 V101 7.702770059094285e-21

R3_102 V3 V102 112965.36124906238
L3_102 V3 V102 -9.474998086440527e-10
C3_102 V3 V102 1.9637175818866485e-20

R3_103 V3 V103 -370072.13263995165
L3_103 V3 V103 3.091218091683128e-09
C3_103 V3 V103 -9.10253650164473e-21

R3_104 V3 V104 6122299.871522031
L3_104 V3 V104 -3.933695827707652e-08
C3_104 V3 V104 1.6181059865341334e-21

R3_105 V3 V105 -312724.53030764294
L3_105 V3 V105 2.251687696214766e-09
C3_105 V3 V105 -6.00818094519479e-21

R3_106 V3 V106 375587.6192235482
L3_106 V3 V106 -2.9222909174056123e-09
C3_106 V3 V106 1.0241156327063715e-20

R3_107 V3 V107 208297.34207327772
L3_107 V3 V107 -1.5802789860916302e-09
C3_107 V3 V107 1.3555297881919346e-20

R3_108 V3 V108 -210395.38875503646
L3_108 V3 V108 1.4807747728499846e-09
C3_108 V3 V108 -1.6854843744313108e-20

R3_109 V3 V109 -703627.2611471334
L3_109 V3 V109 5.162013130884403e-09
C3_109 V3 V109 -6.52313457759655e-21

R3_110 V3 V110 -404570.7676771607
L3_110 V3 V110 2.724721957864103e-09
C3_110 V3 V110 -7.154966457087435e-21

R3_111 V3 V111 -809399.2877592267
L3_111 V3 V111 5.275378374399838e-09
C3_111 V3 V111 -7.433390118871225e-21

R3_112 V3 V112 108370.7680946419
L3_112 V3 V112 -9.932491199880256e-10
C3_112 V3 V112 1.2856996437653444e-20

R3_113 V3 V113 256456.56717689612
L3_113 V3 V113 -2.5155227524140092e-09
C3_113 V3 V113 4.892535325429096e-21

R3_114 V3 V114 376382.9031032974
L3_114 V3 V114 -2.9068533205866427e-09
C3_114 V3 V114 4.523092103435752e-21

R3_115 V3 V115 357544.52235195815
L3_115 V3 V115 -3.201239518470979e-09
C3_115 V3 V115 6.5386897633515066e-21

R3_116 V3 V116 -257953.59973034274
L3_116 V3 V116 2.2016266065352634e-09
C3_116 V3 V116 -8.957671534582295e-21

R3_117 V3 V117 -361198.6253174661
L3_117 V3 V117 3.366670702273682e-09
C3_117 V3 V117 -7.714401574644935e-21

R3_118 V3 V118 -390643.72051342926
L3_118 V3 V118 2.913431185426188e-09
C3_118 V3 V118 -3.4178585229371674e-21

R3_119 V3 V119 -720986.4980290416
L3_119 V3 V119 4.177777837601663e-09
C3_119 V3 V119 -5.201925533444221e-21

R3_120 V3 V120 -1117870.9446688846
L3_120 V3 V120 1.2591474994128446e-08
C3_120 V3 V120 -2.5031894898186875e-21

R3_121 V3 V121 197168.96452689197
L3_121 V3 V121 -2.0778988325307367e-09
C3_121 V3 V121 7.981471228260445e-22

R3_122 V3 V122 102624.36404926426
L3_122 V3 V122 -1.1087853833822426e-09
C3_122 V3 V122 -4.319823569555905e-22

R3_123 V3 V123 611074.6494114053
L3_123 V3 V123 -5.437516408598367e-09
C3_123 V3 V123 -3.862940355347507e-22

R3_124 V3 V124 4276529.299351984
L3_124 V3 V124 4.086012389093889e-06
C3_124 V3 V124 -7.484372429549037e-22

R3_125 V3 V125 -172423.6957989443
L3_125 V3 V125 1.798832688138788e-09
C3_125 V3 V125 -2.2958512759304975e-21

R3_126 V3 V126 -131604.34053282684
L3_126 V3 V126 1.4302448892600144e-09
C3_126 V3 V126 9.684861196598488e-22

R3_127 V3 V127 213943.36210942763
L3_127 V3 V127 -2.205527275369618e-09
C3_127 V3 V127 2.5940508291314723e-22

R3_128 V3 V128 -5732074.363545385
L3_128 V3 V128 6.790026598660893e-06
C3_128 V3 V128 3.1290801967626665e-22

R3_129 V3 V129 533163.8817155148
L3_129 V3 V129 -5.2931423587675046e-09
C3_129 V3 V129 -3.9551619084050114e-22

R3_130 V3 V130 -311893.3306215056
L3_130 V3 V130 2.6263969763735506e-09
C3_130 V3 V130 -4.5138358818833375e-21

R3_131 V3 V131 -584773.8170789717
L3_131 V3 V131 7.850050525677751e-09
C3_131 V3 V131 3.6369571370304284e-21

R3_132 V3 V132 -555601.3709510724
L3_132 V3 V132 5.566020333435782e-09
C3_132 V3 V132 -4.591418789906383e-22

R3_133 V3 V133 -2217121.520779216
L3_133 V3 V133 2.9983865997289206e-08
C3_133 V3 V133 1.473985735128194e-21

R3_134 V3 V134 -444703.08803062333
L3_134 V3 V134 3.6140710844295038e-09
C3_134 V3 V134 7.668602049763361e-22

R3_135 V3 V135 327422.7723109326
L3_135 V3 V135 -3.4281475068779584e-09
C3_135 V3 V135 -1.6277506662336789e-21

R3_136 V3 V136 -2008735.7903697884
L3_136 V3 V136 2.5419764450515585e-08
C3_136 V3 V136 1.142702641644488e-22

R3_137 V3 V137 -262038.9561120554
L3_137 V3 V137 2.7435371047677364e-09
C3_137 V3 V137 -8.924501084506121e-22

R3_138 V3 V138 -126704.26381081539
L3_138 V3 V138 1.317539120267043e-09
C3_138 V3 V138 -8.432098322231441e-22

R3_139 V3 V139 169897.90238451218
L3_139 V3 V139 -1.638440476510434e-09
C3_139 V3 V139 1.4051284893225171e-21

R3_140 V3 V140 -303839.3563012372
L3_140 V3 V140 2.4930012583235193e-09
C3_140 V3 V140 -2.0381018500008405e-21

R3_141 V3 V141 -535540.5472058214
L3_141 V3 V141 5.917156847209993e-09
C3_141 V3 V141 -7.261928064416395e-22

R3_142 V3 V142 -322077.44293551013
L3_142 V3 V142 2.6160346762872783e-09
C3_142 V3 V142 -2.4703121811273372e-21

R3_143 V3 V143 -854021.6763022824
L3_143 V3 V143 8.074856096789057e-09
C3_143 V3 V143 3.6028070409078003e-22

R3_144 V3 V144 313270.5819174327
L3_144 V3 V144 -3.1507724614263237e-09
C3_144 V3 V144 -1.8147534775953028e-22

R4_4 V4 0 15786.89362155807
L4_4 V4 0 -3.108842053130248e-10
C4_4 V4 0 -3.0727748275177625e-21

R4_5 V4 V5 2972386.8168062186
L4_5 V4 V5 -2.789497053327826e-08
C4_5 V4 V5 6.262694348423861e-24

R4_6 V4 V6 3402583.164697048
L4_6 V4 V6 -2.882278590203419e-08
C4_6 V4 V6 -3.667282703538242e-22

R4_7 V4 V7 -24437578.007394675
L4_7 V4 V7 2.820284854947311e-06
C4_7 V4 V7 -1.4918217026106062e-22

R4_8 V4 V8 -140246.97416002175
L4_8 V4 V8 2.0935069591278653e-09
C4_8 V4 V8 1.8162003478949084e-21

R4_9 V4 V9 1174840.3520263867
L4_9 V4 V9 -1.1411317204456841e-08
C4_9 V4 V9 -1.2778761908127059e-21

R4_10 V4 V10 -648209.8083420771
L4_10 V4 V10 9.821472753206748e-09
C4_10 V4 V10 9.826560826086612e-22

R4_11 V4 V11 -424966.1276391337
L4_11 V4 V11 5.969632300538698e-09
C4_11 V4 V11 6.9808648288769045e-22

R4_12 V4 V12 -1199644.2649364127
L4_12 V4 V12 -1.3768868617690625e-09
C4_12 V4 V12 -2.3633514626167484e-22

R4_13 V4 V13 2881205.8142332914
L4_13 V4 V13 3.4374404746986827e-09
C4_13 V4 V13 3.469010105796554e-22

R4_14 V4 V14 3375112.286296263
L4_14 V4 V14 -2.3827642001629706e-09
C4_14 V4 V14 -8.836479252826053e-22

R4_15 V4 V15 12641783.224511584
L4_15 V4 V15 -2.869150288972372e-09
C4_15 V4 V15 -3.067306915573918e-22

R4_16 V4 V16 -606330.4343318718
L4_16 V4 V16 -4.942192323299023e-09
C4_16 V4 V16 1.8668255747402623e-22

R4_17 V4 V17 4502415.440851407
L4_17 V4 V17 -1.4014192411319498e-08
C4_17 V4 V17 -8.850520130440564e-24

R4_18 V4 V18 1804405.857391104
L4_18 V4 V18 3.133859809023345e-08
C4_18 V4 V18 -5.26633699347719e-22

R4_19 V4 V19 -1380224.5277734962
L4_19 V4 V19 4.453123930103176e-08
C4_19 V4 V19 -3.456310177860798e-22

R4_20 V4 V20 -155984.62124826718
L4_20 V4 V20 1.337146532657053e-09
C4_20 V4 V20 2.1134815460252628e-21

R4_21 V4 V21 4284606.224063099
L4_21 V4 V21 2.514005208736217e-08
C4_21 V4 V21 1.6238497796765973e-22

R4_22 V4 V22 -12059015.016705062
L4_22 V4 V22 1.1403378981215683e-08
C4_22 V4 V22 4.052924312573802e-24

R4_23 V4 V23 -1714677.7985984772
L4_23 V4 V23 6.143132593506808e-09
C4_23 V4 V23 2.2437664982313457e-22

R4_24 V4 V24 5809414.805588346
L4_24 V4 V24 -8.987465447276685e-10
C4_24 V4 V24 -2.9656341588395783e-21

R4_25 V4 V25 705631.3759640905
L4_25 V4 V25 -1.9114990268062746e-08
C4_25 V4 V25 8.254562811408631e-22

R4_26 V4 V26 5532282.919096174
L4_26 V4 V26 5.928020489897053e-09
C4_26 V4 V26 9.5948849429437e-22

R4_27 V4 V27 717179.1322114842
L4_27 V4 V27 1.2317785230424083e-07
C4_27 V4 V27 8.114759982379483e-22

R4_28 V4 V28 753946.0135149533
L4_28 V4 V28 -1.2667086473123914e-09
C4_28 V4 V28 -3.682518795326484e-22

R4_29 V4 V29 -1150187.2098915481
L4_29 V4 V29 5.07536279064635e-09
C4_29 V4 V29 -6.567609962173634e-23

R4_30 V4 V30 -598845.4483560851
L4_30 V4 V30 3.98665022744502e-09
C4_30 V4 V30 -2.183977530680712e-22

R4_31 V4 V31 -3544922.859254957
L4_31 V4 V31 9.00393141183924e-09
C4_31 V4 V31 -4.312190160652675e-22

R4_32 V4 V32 665026.0791109602
L4_32 V4 V32 -1.5705735162223998e-09
C4_32 V4 V32 4.543383381696751e-21

R4_33 V4 V33 713860.3610487519
L4_33 V4 V33 -6.402018930905312e-09
C4_33 V4 V33 -1.8961497451754076e-22

R4_34 V4 V34 2877868.25536519
L4_34 V4 V34 -1.8379024667038813e-08
C4_34 V4 V34 -7.666295957557646e-22

R4_35 V4 V35 319249.97591254604
L4_35 V4 V35 -2.1248779520284743e-09
C4_35 V4 V35 5.08349569010188e-22

R4_36 V4 V36 -294471.93551262096
L4_36 V4 V36 4.305130093069756e-09
C4_36 V4 V36 -3.4618366933083014e-21

R4_37 V4 V37 -922977.8985469976
L4_37 V4 V37 7.924453346597087e-09
C4_37 V4 V37 -1.3435843741770868e-21

R4_38 V4 V38 2882294.7985689724
L4_38 V4 V38 -4.022264960074238e-08
C4_38 V4 V38 -2.732541570552159e-21

R4_39 V4 V39 -617603.7846297303
L4_39 V4 V39 6.1621555191766216e-09
C4_39 V4 V39 -1.6944585757765977e-21

R4_40 V4 V40 628121.4573639828
L4_40 V4 V40 -2.617694560817053e-09
C4_40 V4 V40 1.835677145315138e-20

R4_41 V4 V41 7310449.645012031
L4_41 V4 V41 1.8642590872606075e-08
C4_41 V4 V41 -4.289330047143001e-22

R4_42 V4 V42 189652.13475949227
L4_42 V4 V42 -2.2920002810165896e-09
C4_42 V4 V42 3.39452742927052e-21

R4_43 V4 V43 -1524247.0209536196
L4_43 V4 V43 3.103391465543538e-08
C4_43 V4 V43 -9.138437187580732e-22

R4_44 V4 V44 -50474.9262134325
L4_44 V4 V44 4.833214229317767e-10
C4_44 V4 V44 -3.8188907507139514e-20

R4_45 V4 V45 296345.1350028815
L4_45 V4 V45 -3.1633283439399693e-09
C4_45 V4 V45 1.1441474653928097e-20

R4_46 V4 V46 -1213830.1960902044
L4_46 V4 V46 2.5621573128879973e-09
C4_46 V4 V46 -8.55136540057715e-21

R4_47 V4 V47 -558105.2212821179
L4_47 V4 V47 1.0297584012578165e-08
C4_47 V4 V47 1.1635486199806819e-21

R4_48 V4 V48 567270.9559929473
L4_48 V4 V48 -7.201788475620923e-09
C4_48 V4 V48 1.1895628185074077e-20

R4_49 V4 V49 -294007.73901964456
L4_49 V4 V49 5.435746843368572e-09
C4_49 V4 V49 -1.8975117617422265e-21

R4_50 V4 V50 460711.66255948826
L4_50 V4 V50 -5.96913645636656e-08
C4_50 V4 V50 1.2551787230279365e-21

R4_51 V4 V51 -389316.2620094816
L4_51 V4 V51 5.626483742955136e-09
C4_51 V4 V51 -2.5006497293807157e-21

R4_52 V4 V52 -1828671.0634715022
L4_52 V4 V52 3.2904272979096548e-09
C4_52 V4 V52 -1.6369550072636629e-21

R4_53 V4 V53 238688.50241582957
L4_53 V4 V53 -2.2667042870696063e-09
C4_53 V4 V53 9.365367399130481e-21

R4_54 V4 V54 577011.1880563076
L4_54 V4 V54 -5.669971950680042e-09
C4_54 V4 V54 5.131449304278634e-21

R4_55 V4 V55 3764801.7472489807
L4_55 V4 V55 6.041551020081754e-09
C4_55 V4 V55 1.15126764836065e-21

R4_56 V4 V56 -79075.04274711017
L4_56 V4 V56 7.064221990169343e-10
C4_56 V4 V56 -1.0570272072035845e-20

R4_57 V4 V57 527577.1771498076
L4_57 V4 V57 -3.9454289533766705e-09
C4_57 V4 V57 -3.221087465048645e-21

R4_58 V4 V58 174292.94939042183
L4_58 V4 V58 -1.3849218627471415e-09
C4_58 V4 V58 1.8044116097996722e-21

R4_59 V4 V59 1398971.513639106
L4_59 V4 V59 -7.497239811243652e-09
C4_59 V4 V59 8.584502491443297e-22

R4_60 V4 V60 -46912.870583558724
L4_60 V4 V60 5.151065494837879e-10
C4_60 V4 V60 -1.7740271053710406e-21

R4_61 V4 V61 776676.3090105671
L4_61 V4 V61 -5.814487159123931e-09
C4_61 V4 V61 6.3990459839074494e-21

R4_62 V4 V62 -259613.23654927232
L4_62 V4 V62 3.506206457421133e-09
C4_62 V4 V62 -1.3725699452320515e-21

R4_63 V4 V63 -309063.2846728074
L4_63 V4 V63 2.5341370442837903e-09
C4_63 V4 V63 -6.509631158017632e-21

R4_64 V4 V64 351512.88744780497
L4_64 V4 V64 -1.5009906640516124e-09
C4_64 V4 V64 -6.5147540150077205e-21

R4_65 V4 V65 -680673.1995037148
L4_65 V4 V65 6.559742346450412e-09
C4_65 V4 V65 1.1622217855430465e-23

R4_66 V4 V66 174685.56381769947
L4_66 V4 V66 -1.2041316731529185e-09
C4_66 V4 V66 5.711166711003817e-21

R4_67 V4 V67 -776913.8882518326
L4_67 V4 V67 1.1527654751334471e-08
C4_67 V4 V67 -4.171393061644509e-21

R4_68 V4 V68 -88352.91290120059
L4_68 V4 V68 7.423523211821534e-10
C4_68 V4 V68 7.511515404275132e-21

R4_69 V4 V69 133577.12225659628
L4_69 V4 V69 -1.1448013278777912e-09
C4_69 V4 V69 -4.91289346683489e-22

R4_70 V4 V70 6800292.676772209
L4_70 V4 V70 -3.465461425146203e-09
C4_70 V4 V70 1.2778715907491942e-20

R4_71 V4 V71 70631283.68640168
L4_71 V4 V71 5.068730890841065e-08
C4_71 V4 V71 2.471981860518001e-22

R4_72 V4 V72 1158590.0236719395
L4_72 V4 V72 -4.87091682604944e-09
C4_72 V4 V72 -6.87685009538325e-22

R4_73 V4 V73 2046227.1612223855
L4_73 V4 V73 -4.004144009279305e-09
C4_73 V4 V73 1.2097416176352936e-20

R4_74 V4 V74 894092.4092409122
L4_74 V4 V74 -7.046525462229954e-09
C4_74 V4 V74 2.780494015978183e-21

R4_75 V4 V75 -765728.6817879103
L4_75 V4 V75 5.758507660444744e-09
C4_75 V4 V75 -6.547120674170534e-21

R4_76 V4 V76 218787.1973360025
L4_76 V4 V76 -1.8886999738288205e-09
C4_76 V4 V76 1.2536456035338233e-20

R4_77 V4 V77 -221094.8021653315
L4_77 V4 V77 1.5791011125576946e-09
C4_77 V4 V77 -1.4897339550219562e-20

R4_78 V4 V78 338574.9944496311
L4_78 V4 V78 -3.4151680960668663e-09
C4_78 V4 V78 7.699278753004548e-21

R4_79 V4 V79 384835.6422167754
L4_79 V4 V79 -3.0038519063238023e-09
C4_79 V4 V79 8.216697117289998e-21

R4_80 V4 V80 -89259.11148026526
L4_80 V4 V80 7.076592944376643e-10
C4_80 V4 V80 -3.16540059121595e-20

R4_81 V4 V81 47138.45404378871
L4_81 V4 V81 -3.5112655875455627e-10
C4_81 V4 V81 5.9253855062896e-20

R4_82 V4 V82 -174057.1561862835
L4_82 V4 V82 1.3275985313281106e-09
C4_82 V4 V82 -1.881092302099836e-20

R4_83 V4 V83 -79268.31803318947
L4_83 V4 V83 6.077066301813772e-10
C4_83 V4 V83 -3.6139681204352966e-20

R4_84 V4 V84 -410932.9962987309
L4_84 V4 V84 3.0100803176390356e-09
C4_84 V4 V84 -2.8661556721414553e-21

R4_85 V4 V85 255213.5896075951
L4_85 V4 V85 -1.5443820275631534e-09
C4_85 V4 V85 1.273140104283698e-20

R4_86 V4 V86 4057138.564806704
L4_86 V4 V86 -3.048966084386301e-09
C4_86 V4 V86 -9.940108572863026e-22

R4_87 V4 V87 179837.5416021483
L4_87 V4 V87 -1.394063944972504e-09
C4_87 V4 V87 2.1869577116917148e-20

R4_88 V4 V88 190024.24503102523
L4_88 V4 V88 -1.6345329724044345e-09
C4_88 V4 V88 1.8478244699996876e-20

R4_89 V4 V89 -274110.6359389164
L4_89 V4 V89 1.9519959356533652e-09
C4_89 V4 V89 -1.1174145934120901e-20

R4_90 V4 V90 -1775748.1161976825
L4_90 V4 V90 9.964167072303478e-08
C4_90 V4 V90 -1.0871343543199352e-21

R4_91 V4 V91 -13002796.571166405
L4_91 V4 V91 3.3010369216073933e-08
C4_91 V4 V91 -5.884007426947282e-22

R4_92 V4 V92 -49294.32613122003
L4_92 V4 V92 3.974029622978194e-10
C4_92 V4 V92 -5.900881582151957e-20

R4_93 V4 V93 367741.6459806636
L4_93 V4 V93 -2.4856144509497707e-09
C4_93 V4 V93 6.403404496418327e-21

R4_94 V4 V94 107091.63732573751
L4_94 V4 V94 -8.680733974827567e-10
C4_94 V4 V94 2.6636169090688238e-20

R4_95 V4 V95 -647658.3351935808
L4_95 V4 V95 4.113102176517196e-09
C4_95 V4 V95 -7.599968274576103e-21

R4_96 V4 V96 -45391.08365754449
L4_96 V4 V96 3.478628772514738e-10
C4_96 V4 V96 -6.499771190433029e-20

R4_97 V4 V97 150186.98690612864
L4_97 V4 V97 -1.093019179398066e-09
C4_97 V4 V97 2.0163700467042772e-20

R4_98 V4 V98 -133108.0144599741
L4_98 V4 V98 9.579417388906623e-10
C4_98 V4 V98 -2.3530431749261578e-20

R4_99 V4 V99 415745.5833266776
L4_99 V4 V99 -3.44765948737867e-09
C4_99 V4 V99 8.729549830385856e-21

R4_100 V4 V100 114000.59565204472
L4_100 V4 V100 -1.0517017676147375e-09
C4_100 V4 V100 3.1153511226002497e-20

R4_101 V4 V101 -137729.8579567935
L4_101 V4 V101 1.0383197385653264e-09
C4_101 V4 V101 -2.4804528312345865e-20

R4_102 V4 V102 -950133.2591015425
L4_102 V4 V102 3.0853036356464634e-09
C4_102 V4 V102 -6.060925362390266e-21

R4_103 V4 V103 662453.4880996235
L4_103 V4 V103 -4.6803453888170836e-09
C4_103 V4 V103 7.009872989497981e-21

R4_104 V4 V104 -68589.29390438227
L4_104 V4 V104 5.932212338987878e-10
C4_104 V4 V104 -4.3309784769375465e-20

R4_105 V4 V105 95992.32003151182
L4_105 V4 V105 -8.477223058492894e-10
C4_105 V4 V105 3.345602013093944e-20

R4_106 V4 V106 -96358.16877828569
L4_106 V4 V106 7.565864879903329e-10
C4_106 V4 V106 -3.5418643242973895e-20

R4_107 V4 V107 -300778.9498688247
L4_107 V4 V107 2.15317720790056e-09
C4_107 V4 V107 -1.0298359069032539e-20

R4_108 V4 V108 106600.6141762814
L4_108 V4 V108 -9.02534373246663e-10
C4_108 V4 V108 3.5167890705710324e-20

R4_109 V4 V109 -91689.23692485824
L4_109 V4 V109 9.577311015055087e-10
C4_109 V4 V109 -4.114976232395383e-20

R4_110 V4 V110 119069.90009081452
L4_110 V4 V110 -8.850199817874288e-10
C4_110 V4 V110 3.0348153154285623e-20

R4_111 V4 V111 215178.6707597293
L4_111 V4 V111 -1.5880856116651451e-09
C4_111 V4 V111 1.909600260721872e-20

R4_112 V4 V112 -181739.57898982952
L4_112 V4 V112 1.2668999682098793e-09
C4_112 V4 V112 -2.3562240028745395e-20

R4_113 V4 V113 265349.51274737145
L4_113 V4 V113 -4.582895859055499e-09
C4_113 V4 V113 1.5387763260712844e-20

R4_114 V4 V114 -241506.5569785095
L4_114 V4 V114 1.5838760422605957e-09
C4_114 V4 V114 -2.332221597345819e-20

R4_115 V4 V115 -498706.4116264378
L4_115 V4 V115 3.767213176837696e-09
C4_115 V4 V115 -9.41552811696786e-21

R4_116 V4 V116 177964.76286367694
L4_116 V4 V116 -1.2693611863610075e-09
C4_116 V4 V116 2.1920344395347838e-20

R4_117 V4 V117 -1066580.173206302
L4_117 V4 V117 -5.2069241907425525e-08
C4_117 V4 V117 -9.395767217011761e-21

R4_118 V4 V118 -1514757.1249537324
L4_118 V4 V118 -4.2622835445708314e-08
C4_118 V4 V118 -7.713819970203972e-22

R4_119 V4 V119 118094.4204517851
L4_119 V4 V119 -9.262935139935767e-10
C4_119 V4 V119 3.458601241861496e-20

R4_120 V4 V120 217382.4818357329
L4_120 V4 V120 -1.9560064627262344e-09
C4_120 V4 V120 1.960598834829327e-20

R4_121 V4 V121 11956955.58639557
L4_121 V4 V121 -4.7635047836845035e-08
C4_121 V4 V121 -2.017460599048596e-21

R4_122 V4 V122 272671.9882141285
L4_122 V4 V122 -2.8617758465396056e-09
C4_122 V4 V122 -1.4916076081336594e-21

R4_123 V4 V123 479150.11300605745
L4_123 V4 V123 -4.479026236746943e-09
C4_123 V4 V123 -2.5841824579854525e-22

R4_124 V4 V124 321299.56382066634
L4_124 V4 V124 -3.961221506865028e-09
C4_124 V4 V124 1.8879126771478536e-20

R4_125 V4 V125 6168634.380630078
L4_125 V4 V125 -6.930231163781969e-09
C4_125 V4 V125 1.037632830552327e-21

R4_126 V4 V126 -268624.85510003
L4_126 V4 V126 2.450257697627556e-09
C4_126 V4 V126 -1.2531850219067476e-21

R4_127 V4 V127 371376.9762139727
L4_127 V4 V127 -5.898954598156403e-09
C4_127 V4 V127 5.059872392227317e-21

R4_128 V4 V128 396447.72949105396
L4_128 V4 V128 -5.586829434302591e-09
C4_128 V4 V128 -4.303168470655478e-21

R4_129 V4 V129 348840.1953505878
L4_129 V4 V129 -4.33454408653231e-09
C4_129 V4 V129 3.797636657393564e-21

R4_130 V4 V130 -8333778.062785924
L4_130 V4 V130 5.564262717279717e-08
C4_130 V4 V130 -6.622110899822908e-22

R4_131 V4 V131 -293696.63004944613
L4_131 V4 V131 2.8258069373551423e-09
C4_131 V4 V131 -6.179073139536321e-21

R4_132 V4 V132 820899.0500723992
L4_132 V4 V132 -3.555641136455742e-09
C4_132 V4 V132 9.136683786692658e-21

R4_133 V4 V133 -357262.95620533393
L4_133 V4 V133 2.557057518698972e-09
C4_133 V4 V133 -8.522460582434967e-21

R4_134 V4 V134 -1856761.9385447644
L4_134 V4 V134 1.4472652984920086e-08
C4_134 V4 V134 -7.864920672648091e-23

R4_135 V4 V135 473611.2118755299
L4_135 V4 V135 -6.028201890604522e-09
C4_135 V4 V135 3.0740295400670435e-21

R4_136 V4 V136 1324151.809030022
L4_136 V4 V136 -1.788453987007506e-08
C4_136 V4 V136 2.171977052273406e-21

R4_137 V4 V137 613328.3365683822
L4_137 V4 V137 -1.5212824499258936e-08
C4_137 V4 V137 1.108840737284475e-20

R4_138 V4 V138 -344652.99946104037
L4_138 V4 V138 2.6576928318748964e-09
C4_138 V4 V138 8.566964440072764e-21

R4_139 V4 V139 681210.688956758
L4_139 V4 V139 -5.8470988018808915e-09
C4_139 V4 V139 -2.161048408890155e-21

R4_140 V4 V140 683938.0602857488
L4_140 V4 V140 -4.244220050900778e-09
C4_140 V4 V140 1.5819092623265472e-21

R4_141 V4 V141 -647255.8244867182
L4_141 V4 V141 9.546281989358019e-09
C4_141 V4 V141 1.5260220111241854e-21

R4_142 V4 V142 53137990.025273144
L4_142 V4 V142 1.1582479680562114e-08
C4_142 V4 V142 5.3369315467474154e-21

R4_143 V4 V143 -2249089.2991456212
L4_143 V4 V143 8.731317190286272e-09
C4_143 V4 V143 2.0477063206657653e-21

R4_144 V4 V144 5495129.018577243
L4_144 V4 V144 4.08100163870233e-09
C4_144 V4 V144 -3.580585951838305e-21

R5_5 V5 0 858.8135290597778
L5_5 V5 0 -4.987102308527547e-13
C5_5 V5 0 -6.174601043946447e-19

R5_6 V5 V6 991390.507499064
L5_6 V5 V6 -2.265211815936951e-10
C5_6 V5 V6 8.854576034742471e-22

R5_7 V5 V7 580348.0781299584
L5_7 V5 V7 -3.249510960190535e-09
C5_7 V5 V7 9.434662104028838e-22

R5_8 V5 V8 -319093.98064241017
L5_8 V5 V8 -1.7617252905808556e-10
C5_8 V5 V8 3.55179588979021e-22

R5_9 V5 V9 66544.59419078132
L5_9 V5 V9 -5.2052594775024706e-11
C5_9 V5 V9 1.2885067922701199e-20

R5_10 V5 V10 129268.96739250285
L5_10 V5 V10 -4.3185250124270433e-10
C5_10 V5 V10 1.6617545839310247e-21

R5_11 V5 V11 87244.03790850777
L5_11 V5 V11 -2.0933008031266174e-10
C5_11 V5 V11 5.867705705219233e-21

R5_12 V5 V12 -894716.1295059356
L5_12 V5 V12 6.785994430267609e-10
C5_12 V5 V12 -1.5908631105810588e-21

R5_13 V5 V13 -89869.59110598927
L5_13 V5 V13 -7.595103185738952e-10
C5_13 V5 V13 -3.1554158299038816e-21

R5_14 V5 V14 -504927.3173222829
L5_14 V5 V14 -9.354001585507514e-11
C5_14 V5 V14 8.648147816999356e-22

R5_15 V5 V15 -195555.67170080013
L5_15 V5 V15 -1.8426710659707098e-08
C5_15 V5 V15 -2.6588144620539592e-21

R5_16 V5 V16 -388600.6798158074
L5_16 V5 V16 -2.5994445161807447e-10
C5_16 V5 V16 -6.84722048113226e-22

R5_17 V5 V17 -34058.1047134944
L5_17 V5 V17 -5.301970762546698e-11
C5_17 V5 V17 -7.410271849731504e-21

R5_18 V5 V18 2605026.729079143
L5_18 V5 V18 -1.8929864523795036e-10
C5_18 V5 V18 1.5267411491527453e-21

R5_19 V5 V19 -60797.209497330994
L5_19 V5 V19 -5.2210601226145536e-11
C5_19 V5 V19 -2.7471095935863757e-21

R5_20 V5 V20 506517.6859081943
L5_20 V5 V20 1.09335496299042e-09
C5_20 V5 V20 9.32618120809727e-22

R5_21 V5 V21 39330.1716474382
L5_21 V5 V21 -9.97686657903912e-12
C5_21 V5 V21 1.6191335009093347e-20

R5_22 V5 V22 -294242.4919334115
L5_22 V5 V22 8.163496644532626e-11
C5_22 V5 V22 -2.8095265061904294e-21

R5_23 V5 V23 -222943.94238764475
L5_23 V5 V23 9.438288969943372e-11
C5_23 V5 V23 -3.3267096856773584e-21

R5_24 V5 V24 -1341983.2973148206
L5_24 V5 V24 1.0264565836299891e-10
C5_24 V5 V24 -9.259715105469734e-22

R5_25 V5 V25 -30222.42942070447
L5_25 V5 V25 -2.4913690369609994e-11
C5_25 V5 V25 -1.1968790868410529e-21

R5_26 V5 V26 504657.23348136403
L5_26 V5 V26 4.966350566840845e-10
C5_26 V5 V26 -1.415685239803965e-23

R5_27 V5 V27 205259.27997335466
L5_27 V5 V27 -4.227464415372454e-10
C5_27 V5 V27 3.809568353476624e-22

R5_28 V5 V28 -1643476.937286475
L5_28 V5 V28 -1.5609785869861788e-10
C5_28 V5 V28 -1.080912845431664e-21

R5_29 V5 V29 120236.69620156403
L5_29 V5 V29 -1.2999549606973689e-11
C5_29 V5 V29 -3.3154536820824035e-20

R5_30 V5 V30 899575.4186185261
L5_30 V5 V30 3.0434691531364977e-10
C5_30 V5 V30 -3.467788272589393e-21

R5_31 V5 V31 158147.71093184245
L5_31 V5 V31 5.445092359578178e-10
C5_31 V5 V31 -8.28131120444471e-21

R5_32 V5 V32 431509.0207482572
L5_32 V5 V32 2.503257201563696e-10
C5_32 V5 V32 -2.6127307178848213e-21

R5_33 V5 V33 -23630.660686288866
L5_33 V5 V33 1.319992341733803e-11
C5_33 V5 V33 3.517172188073632e-20

R5_34 V5 V34 40327.032152321284
L5_34 V5 V34 -3.466010866618466e-11
C5_34 V5 V34 -1.207002887597591e-20

R5_35 V5 V35 -43710.845276361295
L5_35 V5 V35 2.5866343118774708e-11
C5_35 V5 V35 1.86582823235369e-20

R5_36 V5 V36 120629.19239877237
L5_36 V5 V36 -6.127139608265703e-11
C5_36 V5 V36 -3.1747967218763168e-21

R5_37 V5 V37 -14984.343716108478
L5_37 V5 V37 -5.071890036039024e-12
C5_37 V5 V37 -8.144730808742436e-20

R5_38 V5 V38 -87241.08466842493
L5_38 V5 V38 -8.893155523166639e-11
C5_38 V5 V38 -1.5840196353326897e-21

R5_39 V5 V39 -22440.956256845
L5_39 V5 V39 -6.277485519621775e-12
C5_39 V5 V39 -7.02275834849336e-20

R5_40 V5 V40 -62769.64831787369
L5_40 V5 V40 -1.0187536446527059e-10
C5_40 V5 V40 -4.276950230454871e-21

R5_41 V5 V41 -113196.90770797928
L5_41 V5 V41 1.5759502409191027e-12
C5_41 V5 V41 2.4398511168125983e-19

R5_42 V5 V42 19325.754310760814
L5_42 V5 V42 2.1773746403766194e-12
C5_42 V5 V42 1.8113233847955733e-19

R5_43 V5 V43 37779.934447615575
L5_43 V5 V43 4.494645056793645e-12
C5_43 V5 V43 9.494886941201744e-20

R5_44 V5 V44 53046.69673819033
L5_44 V5 V44 8.25708873116171e-11
C5_44 V5 V44 8.348234484969353e-21

R5_45 V5 V45 -5620.608507045548
L5_45 V5 V45 -4.4382918272001024e-12
C5_45 V5 V45 -1.744462114592776e-19

R5_46 V5 V46 -8185.471227500612
L5_46 V5 V46 -3.475919479314238e-11
C5_46 V5 V46 -7.200797526002005e-20

R5_47 V5 V47 -12687.33883237855
L5_47 V5 V47 5.0366083672299764e-11
C5_47 V5 V47 -2.728728532806237e-20

R5_48 V5 V48 147904.50842171762
L5_48 V5 V48 -2.526189954476457e-11
C5_48 V5 V48 -9.97815007396678e-21

R5_49 V5 V49 25561.292793389504
L5_49 V5 V49 -8.131184909105563e-11
C5_49 V5 V49 4.7505344461134264e-20

R5_50 V5 V50 -24475.333206341624
L5_50 V5 V50 1.3956335900174148e-11
C5_50 V5 V50 3.7390717413882834e-20

R5_51 V5 V51 39332.55107912229
L5_51 V5 V51 -1.0379180434754164e-11
C5_51 V5 V51 -3.3483127782409e-20

R5_52 V5 V52 71354.02162294924
L5_52 V5 V52 1.0925692367989756e-11
C5_52 V5 V52 1.154881242119258e-19

R5_53 V5 V53 -20089.445543289483
L5_53 V5 V53 5.718498040267285e-10
C5_53 V5 V53 5.87960127930703e-20

R5_54 V5 V54 -13580.866802175175
L5_54 V5 V54 2.3413753682636062e-11
C5_54 V5 V54 7.879252581226536e-21

R5_55 V5 V55 -16166.261472225273
L5_55 V5 V55 9.378121546351602e-12
C5_55 V5 V55 3.56328145090925e-20

R5_56 V5 V56 -24385.347410806346
L5_56 V5 V56 1.2986966359448862e-11
C5_56 V5 V56 2.4990070677453004e-20

R5_57 V5 V57 -1659.3099737936725
L5_57 V5 V57 1.65146620513807e-12
C5_57 V5 V57 -2.8219359219974654e-20

R5_58 V5 V58 -6892.2259084235
L5_58 V5 V58 8.350629056260215e-12
C5_58 V5 V58 -1.6214094248219125e-20

R5_59 V5 V59 -19745.747994243542
L5_59 V5 V59 -2.0893960430488883e-10
C5_59 V5 V59 -1.892686982137172e-20

R5_60 V5 V60 -10469.490989334789
L5_60 V5 V60 1.3169388631754668e-11
C5_60 V5 V60 -5.6770374891591665e-21

R5_61 V5 V61 4645.427864180235
L5_61 V5 V61 -8.874281370556565e-12
C5_61 V5 V61 8.455609603049775e-20

R5_62 V5 V62 4409.032630563449
L5_62 V5 V62 -1.308133788459353e-11
C5_62 V5 V62 7.461669719090532e-20

R5_63 V5 V63 18933.440436507783
L5_63 V5 V63 1.3028490994509583e-11
C5_63 V5 V63 1.204669305220798e-20

R5_64 V5 V64 -37172.90542114425
L5_64 V5 V64 -3.6226067505758937e-11
C5_64 V5 V64 4.347443808027652e-21

R5_65 V5 V65 -3141.8013550079154
L5_65 V5 V65 1.0811741382609301e-11
C5_65 V5 V65 3.245274401639012e-20

R5_66 V5 V66 -3058.7066069655216
L5_66 V5 V66 -3.1281105951217256e-11
C5_66 V5 V66 2.222967005965743e-20

R5_67 V5 V67 -17583.70194072909
L5_67 V5 V67 6.433952477278784e-11
C5_67 V5 V67 1.3006092901090824e-20

R5_68 V5 V68 -134539.09569508012
L5_68 V5 V68 2.1964477708273167e-11
C5_68 V5 V68 7.466930183035478e-21

R5_69 V5 V69 15894.561779982203
L5_69 V5 V69 -1.1212778566004465e-10
C5_69 V5 V69 -8.753572045814547e-21

R5_70 V5 V70 9238.273712124492
L5_70 V5 V70 1.2925142945056885e-11
C5_70 V5 V70 -2.3346732528590123e-21

R5_71 V5 V71 19359.788302345012
L5_71 V5 V71 1.2388386200919898e-11
C5_71 V5 V71 -4.236576339737123e-22

R5_72 V5 V72 6972.783076075042
L5_72 V5 V72 1.1762592228167277e-11
C5_72 V5 V72 -8.09493771580586e-21

R5_73 V5 V73 18510.775805922185
L5_73 V5 V73 1.314206506123107e-11
C5_73 V5 V73 6.58222828930948e-21

R5_74 V5 V74 14310.890870866739
L5_74 V5 V74 1.218241506319499e-10
C5_74 V5 V74 -1.19755655920354e-20

R5_75 V5 V75 -14664.609989555793
L5_75 V5 V75 -4.493881073535587e-11
C5_75 V5 V75 1.463970260275909e-20

R5_76 V5 V76 -15343.053588354176
L5_76 V5 V76 -1.9542686813053906e-11
C5_76 V5 V76 1.399018912046788e-20

R5_77 V5 V77 -36350.53428635226
L5_77 V5 V77 -1.2452136765282342e-10
C5_77 V5 V77 6.902168776685461e-21

R5_78 V5 V78 -92714.34778065978
L5_78 V5 V78 -2.7554811022484278e-11
C5_78 V5 V78 1.6262527071359466e-21

R5_79 V5 V79 20695.50047814798
L5_79 V5 V79 2.7856665099573477e-11
C5_79 V5 V79 4.507981356344964e-21

R5_80 V5 V80 23239.988279583315
L5_80 V5 V80 1.5628897262103394e-11
C5_80 V5 V80 7.727910302399977e-21

R5_81 V5 V81 48369.73170899046
L5_81 V5 V81 1.4226885233208357e-10
C5_81 V5 V81 -7.057279527827001e-21

R5_82 V5 V82 -109759.01305655272
L5_82 V5 V82 7.701054029106554e-11
C5_82 V5 V82 1.661008292830703e-20

R5_83 V5 V83 73693.81689907494
L5_83 V5 V83 1.9279737616834965e-11
C5_83 V5 V83 5.170416801774679e-21

R5_84 V5 V84 64380.20945334605
L5_84 V5 V84 -5.24218311614153e-10
C5_84 V5 V84 -1.1175064059358957e-20

R5_85 V5 V85 29162.6912776333
L5_85 V5 V85 -1.5076109056884191e-09
C5_85 V5 V85 -1.1516258059307624e-20

R5_86 V5 V86 73905.57334629718
L5_86 V5 V86 -3.808397222471722e-11
C5_86 V5 V86 -9.810570644790703e-21

R5_87 V5 V87 -85738.96397706954
L5_87 V5 V87 -1.648110760218388e-11
C5_87 V5 V87 -8.858794985472327e-21

R5_88 V5 V88 100978.964249082
L5_88 V5 V88 -2.240229406878102e-11
C5_88 V5 V88 2.193036239810135e-21

R5_89 V5 V89 -185291.47259330144
L5_89 V5 V89 8.901833352245007e-12
C5_89 V5 V89 2.6654783108815313e-20

R5_90 V5 V90 -255669.0976322931
L5_90 V5 V90 4.171323948755962e-11
C5_90 V5 V90 2.6486237075253965e-21

R5_91 V5 V91 105004.42296930193
L5_91 V5 V91 2.2701567428670387e-11
C5_91 V5 V91 1.2618699559554493e-20

R5_92 V5 V92 115511.43980697944
L5_92 V5 V92 2.29576600606472e-11
C5_92 V5 V92 9.854917913828347e-21

R5_93 V5 V93 9296.12933874876
L5_93 V5 V93 3.246511182663285e-10
C5_93 V5 V93 7.192506489091625e-21

R5_94 V5 V94 26518.29234073515
L5_94 V5 V94 -1.5190835776227006e-11
C5_94 V5 V94 -9.177405233996752e-21

R5_95 V5 V95 47985.007045140126
L5_95 V5 V95 1.8039817335343509e-10
C5_95 V5 V95 6.591874721785694e-21

R5_96 V5 V96 -1150319.6548551843
L5_96 V5 V96 1.789114977921746e-10
C5_96 V5 V96 1.5499831987828752e-21

R5_97 V5 V97 -96490.52252927498
L5_97 V5 V97 1.6955042424078562e-11
C5_97 V5 V97 -9.635482036037375e-22

R5_98 V5 V98 -26954.36589316911
L5_98 V5 V98 7.458561804744667e-12
C5_98 V5 V98 1.1448313040157584e-20

R5_99 V5 V99 90891.72542671215
L5_99 V5 V99 -1.7127978415580772e-10
C5_99 V5 V99 -1.5446107799588066e-21

R5_100 V5 V100 -158493.6910038964
L5_100 V5 V100 -9.244576393562225e-11
C5_100 V5 V100 -1.2737916732334611e-21

R5_101 V5 V101 32319.612790887688
L5_101 V5 V101 7.031776514180716e-12
C5_101 V5 V101 2.621105120910575e-20

R5_102 V5 V102 71098.15857074349
L5_102 V5 V102 9.727824202583617e-12
C5_102 V5 V102 1.616781471859665e-20

R5_103 V5 V103 534188.2792311846
L5_103 V5 V103 2.550212887446738e-11
C5_103 V5 V103 7.742237257668377e-21

R5_104 V5 V104 63971.16515184944
L5_104 V5 V104 -2.368302657451725e-10
C5_104 V5 V104 -4.045015198772486e-23

R5_105 V5 V105 -57670.528400318384
L5_105 V5 V105 -1.6052991937428495e-11
C5_105 V5 V105 -9.077042938205775e-21

R5_106 V5 V106 29577.35657803269
L5_106 V5 V106 6.972813327302782e-11
C5_106 V5 V106 1.452663798078109e-20

R5_107 V5 V107 -77505.31942660492
L5_107 V5 V107 4.951744064663001e-11
C5_107 V5 V107 -1.3518691878071887e-21

R5_108 V5 V108 -16523.44227275048
L5_108 V5 V108 -1.5615588582026958e-11
C5_108 V5 V108 -2.2228672150859864e-20

R5_109 V5 V109 -30900.532221886882
L5_109 V5 V109 1.3106823796020687e-10
C5_109 V5 V109 -7.832072393004881e-21

R5_110 V5 V110 -105004.64322473112
L5_110 V5 V110 -1.1425501711413665e-11
C5_110 V5 V110 -1.7630699770185596e-20

R5_111 V5 V111 -17755.640200623166
L5_111 V5 V111 2.1966309907301267e-11
C5_111 V5 V111 9.33733226393788e-22

R5_112 V5 V112 -13091.3507698348
L5_112 V5 V112 5.646902121001693e-12
C5_112 V5 V112 1.7078003642906146e-20

R5_113 V5 V113 -22317.187942853525
L5_113 V5 V113 1.5601165212486712e-11
C5_113 V5 V113 6.835289086518655e-21

R5_114 V5 V114 56907.12829848429
L5_114 V5 V114 1.8135185433477797e-11
C5_114 V5 V114 8.255109227398404e-21

R5_115 V5 V115 58374.93835957076
L5_115 V5 V115 3.1748948149756264e-10
C5_115 V5 V115 -1.7194022285449524e-21

R5_116 V5 V116 -212339.84476028406
L5_116 V5 V116 -1.8942673385353875e-11
C5_116 V5 V116 -1.253113560602434e-20

R5_117 V5 V117 51270.64456991395
L5_117 V5 V117 -1.719729495614924e-11
C5_117 V5 V117 -1.2451616460385107e-20

R5_118 V5 V118 1140101.8609005918
L5_118 V5 V118 -1.752499606344041e-11
C5_118 V5 V118 -6.751000063683003e-21

R5_119 V5 V119 -13366.476646260242
L5_119 V5 V119 -1.1233235033247703e-10
C5_119 V5 V119 -9.574036369713243e-21

R5_120 V5 V120 10204.821918320557
L5_120 V5 V120 -9.814368537267449e-12
C5_120 V5 V120 -1.3862595255807256e-21

R5_121 V5 V121 -6718.950259535794
L5_121 V5 V121 7.454740655469391e-12
C5_121 V5 V121 -3.7785315907489054e-22

R5_122 V5 V122 -6344.444426511977
L5_122 V5 V122 7.037535870653589e-12
C5_122 V5 V122 -6.656368615802763e-22

R5_123 V5 V123 -204939.18174920097
L5_123 V5 V123 3.539516064768798e-11
C5_123 V5 V123 -1.8538268421784627e-22

R5_124 V5 V124 -86040.32139328081
L5_124 V5 V124 4.9955789896178035e-11
C5_124 V5 V124 6.89422385790499e-22

R5_125 V5 V125 5431.514965085472
L5_125 V5 V125 -5.39906692153871e-12
C5_125 V5 V125 -3.3819908493087506e-21

R5_126 V5 V126 14832.829133072077
L5_126 V5 V126 -2.5580226091356307e-11
C5_126 V5 V126 1.7126178346536683e-21

R5_127 V5 V127 3053288.033271902
L5_127 V5 V127 -2.794538909751424e-10
C5_127 V5 V127 5.382957599484584e-22

R5_128 V5 V128 142413.5051413554
L5_128 V5 V128 -3.7195593805162506e-10
C5_128 V5 V128 7.616215002864285e-22

R5_129 V5 V129 134022.1930980775
L5_129 V5 V129 8.2032564604041e-11
C5_129 V5 V129 -2.8677889825462056e-21

R5_130 V5 V130 -155936.42186869256
L5_130 V5 V130 -3.5528478922016074e-11
C5_130 V5 V130 -3.8571247689984016e-21

R5_131 V5 V131 39631.032554228106
L5_131 V5 V131 -4.213761826457299e-11
C5_131 V5 V131 -1.3322703911626283e-22

R5_132 V5 V132 81995.51017270745
L5_132 V5 V132 -7.41958027543954e-11
C5_132 V5 V132 -6.992089247646697e-22

R5_133 V5 V133 30407.527053705457
L5_133 V5 V133 -3.4333868835475414e-11
C5_133 V5 V133 5.761803611375925e-21

R5_134 V5 V134 59139.51534748704
L5_134 V5 V134 -1.556772626604057e-11
C5_134 V5 V134 3.517362015749886e-21

R5_135 V5 V135 -89904.62528119303
L5_135 V5 V135 -3.13289689688268e-10
C5_135 V5 V135 1.0207221009908744e-21

R5_136 V5 V136 71623.39786569188
L5_136 V5 V136 -7.64028008418665e-11
C5_136 V5 V136 -1.8797739782563792e-22

R5_137 V5 V137 8791.997994337687
L5_137 V5 V137 -1.0520116212995968e-11
C5_137 V5 V137 -2.519974348177449e-21

R5_138 V5 V138 13644.473755417257
L5_138 V5 V138 -1.4462045438736837e-11
C5_138 V5 V138 4.160394661948146e-21

R5_139 V5 V139 71521.00518698701
L5_139 V5 V139 -6.786446859365793e-10
C5_139 V5 V139 -3.574126658233496e-21

R5_140 V5 V140 -421253.5275002841
L5_140 V5 V140 -1.926306093489689e-11
C5_140 V5 V140 -6.650192340821118e-21

R5_141 V5 V141 32274.079386277026
L5_141 V5 V141 -5.910275394788071e-11
C5_141 V5 V141 -1.4007681274822488e-22

R5_142 V5 V142 -41518.669530981686
L5_142 V5 V142 -2.3290537386955285e-11
C5_142 V5 V142 -4.971301893849911e-21

R5_143 V5 V143 -61756.191650909306
L5_143 V5 V143 3.993964615100077e-11
C5_143 V5 V143 1.830396242402363e-21

R5_144 V5 V144 -24773.296045269726
L5_144 V5 V144 2.1083886277255074e-11
C5_144 V5 V144 6.893404850099129e-21

R6_6 V6 0 2717.2812046152353
L6_6 V6 0 1.7973947220856997e-12
C6_6 V6 0 1.4188828326199288e-19

R6_7 V6 V7 389924.7439279369
L6_7 V6 V7 -1.937336208466521e-09
C6_7 V6 V7 5.502001954020769e-22

R6_8 V6 V8 5767747.970153708
L6_8 V6 V8 -2.426252341094827e-10
C6_8 V6 V8 5.5062317547109225e-22

R6_9 V6 V9 -526891.2222454277
L6_9 V6 V9 5.8372245985148e-10
C6_9 V6 V9 -2.6135003428887672e-21

R6_10 V6 V10 2707378.737843721
L6_10 V6 V10 -3.162610492988564e-11
C6_10 V6 V10 1.0919801015085467e-21

R6_11 V6 V11 2502959.571642687
L6_11 V6 V11 3.9730082289156645e-11
C6_11 V6 V11 -1.1048695529823775e-21

R6_12 V6 V12 -1680964.9417464389
L6_12 V6 V12 1.2545615050805592e-10
C6_12 V6 V12 -4.3481557147463205e-22

R6_13 V6 V13 569270.9281542347
L6_13 V6 V13 -2.405474291268187e-10
C6_13 V6 V13 1.2836661174120677e-21

R6_14 V6 V14 -1560544.1598931903
L6_14 V6 V14 -6.582826788206654e-11
C6_14 V6 V14 -2.3782542436256824e-22

R6_15 V6 V15 205275.43758191238
L6_15 V6 V15 -8.671701447778938e-11
C6_15 V6 V15 1.0575185081458106e-22

R6_16 V6 V16 -1398004.7389937905
L6_16 V6 V16 -1.9125793169646568e-10
C6_16 V6 V16 2.72823409009155e-22

R6_17 V6 V17 351737.3099392306
L6_17 V6 V17 -5.799325554408697e-11
C6_17 V6 V17 1.559435627644987e-21

R6_18 V6 V18 -250776.98050922083
L6_18 V6 V18 -2.5482567881093555e-10
C6_18 V6 V18 1.4832834070513032e-22

R6_19 V6 V19 -5643010.845310859
L6_19 V6 V19 -3.697184938933312e-10
C6_19 V6 V19 1.1772678664113832e-21

R6_20 V6 V20 -823393.1109424843
L6_20 V6 V20 1.8416638071752477e-09
C6_20 V6 V20 3.7909890507694374e-22

R6_21 V6 V21 -356289.18337197625
L6_21 V6 V21 1.6528034052449552e-10
C6_21 V6 V21 -1.9581324592800423e-21

R6_22 V6 V22 375463.9446778319
L6_22 V6 V22 -8.321208715383839e-12
C6_22 V6 V22 3.3627014490468434e-21

R6_23 V6 V23 -711644.0813469662
L6_23 V6 V23 5.624745904623516e-11
C6_23 V6 V23 -8.182121674949471e-22

R6_24 V6 V24 -1387397.993265652
L6_24 V6 V24 5.784208889177837e-11
C6_24 V6 V24 -4.329871154292987e-22

R6_25 V6 V25 162648.20460183136
L6_25 V6 V25 1.2834765283065634e-10
C6_25 V6 V25 -3.760066100574181e-22

R6_26 V6 V26 1239685.1451376507
L6_26 V6 V26 -1.6838214586590524e-11
C6_26 V6 V26 9.598571816247621e-22

R6_27 V6 V27 201966.22429559918
L6_27 V6 V27 -7.383814470941875e-11
C6_27 V6 V27 1.4739375552510425e-22

R6_28 V6 V28 492805.9273401314
L6_28 V6 V28 -8.123463875037502e-11
C6_28 V6 V28 -6.605834986554627e-22

R6_29 V6 V29 -252031.15026227158
L6_29 V6 V29 6.838415061393829e-11
C6_29 V6 V29 4.79281512380139e-21

R6_30 V6 V30 459832.7387640071
L6_30 V6 V30 -1.2738937652308256e-11
C6_30 V6 V30 -4.319964254699583e-21

R6_31 V6 V31 -414738.0760533878
L6_31 V6 V31 6.94911599410197e-11
C6_31 V6 V31 3.1432873267914007e-21

R6_32 V6 V32 -392167.20966001134
L6_32 V6 V32 7.498907080426499e-11
C6_32 V6 V32 1.5727041731863447e-21

R6_33 V6 V33 109023.28291965861
L6_33 V6 V33 -3.511717674251194e-11
C6_33 V6 V33 -2.6313970171438495e-21

R6_34 V6 V34 -231667.96933818597
L6_34 V6 V34 6.50751598692695e-11
C6_34 V6 V34 4.117762615347914e-21

R6_35 V6 V35 76981.24864471515
L6_35 V6 V35 -6.472401553807937e-11
C6_35 V6 V35 -2.1989071045846525e-21

R6_36 V6 V36 819065.0580182319
L6_36 V6 V36 -3.248478137209975e-10
C6_36 V6 V36 -5.529657211257053e-22

R6_37 V6 V37 204500.10597388266
L6_37 V6 V37 3.131021925499893e-11
C6_37 V6 V37 1.2069498571136175e-20

R6_38 V6 V38 -54888.206788993004
L6_38 V6 V38 -1.8577328127139163e-11
C6_38 V6 V38 -1.3934706356583608e-20

R6_39 V6 V39 -664449.9798310978
L6_39 V6 V39 7.713547670011343e-11
C6_39 V6 V39 9.675796521594165e-21

R6_40 V6 V40 -407029.0873025103
L6_40 V6 V40 1.3791707230247753e-10
C6_40 V6 V40 5.0641807319105186e-21

R6_41 V6 V41 -96292.66923635647
L6_41 V6 V41 -8.106797754138459e-12
C6_41 V6 V41 -5.3428392337060333e-20

R6_42 V6 V42 52505.47091722444
L6_42 V6 V42 8.7598697329256e-12
C6_42 V6 V42 2.6653066031983762e-20

R6_43 V6 V43 55610.708017966324
L6_43 V6 V43 -1.7668183265901787e-11
C6_43 V6 V43 -2.3203930113589926e-20

R6_44 V6 V44 133620.61317326268
L6_44 V6 V44 -1.1511813784951951e-10
C6_44 V6 V44 -7.360039171604321e-21

R6_45 V6 V45 90849.00793741428
L6_45 V6 V45 6.197359674767828e-11
C6_45 V6 V45 2.064810865327604e-20

R6_46 V6 V46 -269338.47016647144
L6_46 V6 V46 -2.954370687782755e-11
C6_46 V6 V46 -1.2031561041178189e-20

R6_47 V6 V47 19289.00405621872
L6_47 V6 V47 -4.71698397945658e-11
C6_47 V6 V47 1.3197817663343249e-20

R6_48 V6 V48 76511.3374854073
L6_48 V6 V48 -4.905170518755641e-11
C6_48 V6 V48 2.07479131714439e-21

R6_49 V6 V49 -52749.20283570598
L6_49 V6 V49 8.662384818453811e-10
C6_49 V6 V49 -6.963723368039733e-21

R6_50 V6 V50 -716227.5506561177
L6_50 V6 V50 -1.903037616413512e-10
C6_50 V6 V50 -4.261226146084863e-22

R6_51 V6 V51 58245.74314808206
L6_51 V6 V51 1.4225343421322517e-10
C6_51 V6 V51 -2.1445403253375962e-20

R6_52 V6 V52 -83928.38527460594
L6_52 V6 V52 8.639154784727175e-11
C6_52 V6 V52 -1.2368517080298027e-20

R6_53 V6 V53 -289397.64818393753
L6_53 V6 V53 -1.4893205428967124e-11
C6_53 V6 V53 -1.8269620666680585e-20

R6_54 V6 V54 188620.59962592114
L6_54 V6 V54 2.0470238435285105e-09
C6_54 V6 V54 8.95231971926437e-21

R6_55 V6 V55 -57556.38793108768
L6_55 V6 V55 -1.8885792398370095e-10
C6_55 V6 V55 -8.121491308895176e-21

R6_56 V6 V56 -76462.36476739848
L6_56 V6 V56 -2.3243810605858065e-11
C6_56 V6 V56 -1.8229887960420135e-20

R6_57 V6 V57 11147.671857551111
L6_57 V6 V57 -1.9652887453598487e-11
C6_57 V6 V57 6.538569490781065e-21

R6_58 V6 V58 -9436.002598856554
L6_58 V6 V58 7.580224861873263e-12
C6_58 V6 V58 -5.0535653050412976e-21

R6_59 V6 V59 102559.65900523918
L6_59 V6 V59 -1.5250090118789825e-10
C6_59 V6 V59 -1.6063332168890376e-21

R6_60 V6 V60 39767.19562013825
L6_60 V6 V60 -2.892717750320697e-11
C6_60 V6 V60 -2.5931131053082593e-21

R6_61 V6 V61 -22447.960195263266
L6_61 V6 V61 -2.6875538705437005e-11
C6_61 V6 V61 -1.8298244824298713e-20

R6_62 V6 V62 90424.76115554532
L6_62 V6 V62 5.0388640886974e-11
C6_62 V6 V62 1.2690041464547822e-21

R6_63 V6 V63 -11931.298900040709
L6_63 V6 V63 3.1003626910129705e-11
C6_63 V6 V63 -2.418265258225482e-20

R6_64 V6 V64 -44047.7044016744
L6_64 V6 V64 -1.8934275697011292e-11
C6_64 V6 V64 -1.5837353741408693e-20

R6_65 V6 V65 45799.499285038095
L6_65 V6 V65 2.1986667356744295e-10
C6_65 V6 V65 -1.320812970213747e-21

R6_66 V6 V66 -21673.431338322433
L6_66 V6 V66 -1.0395487195120103e-11
C6_66 V6 V66 -3.8890891009873925e-21

R6_67 V6 V67 8938.549210426456
L6_67 V6 V67 3.219982083869962e-11
C6_67 V6 V67 -1.0637758230569332e-20

R6_68 V6 V68 44343.212734908826
L6_68 V6 V68 6.292333591422458e-11
C6_68 V6 V68 -2.071756237964705e-21

R6_69 V6 V69 22695.526010728405
L6_69 V6 V69 3.962503870192932e-10
C6_69 V6 V69 -3.413075086016795e-21

R6_70 V6 V70 -22485.27481730858
L6_70 V6 V70 -1.1296137483078932e-11
C6_70 V6 V70 -9.654825505039087e-21

R6_71 V6 V71 -6859.659297135293
L6_71 V6 V71 -5.665247132036655e-12
C6_71 V6 V71 -4.843076032832565e-21

R6_72 V6 V72 22545.266046516736
L6_72 V6 V72 3.083093974456965e-11
C6_72 V6 V72 -1.697320895863448e-21

R6_73 V6 V73 18920.714248017073
L6_73 V6 V73 2.6780189644976715e-11
C6_73 V6 V73 2.5404892109854847e-22

R6_74 V6 V74 25420.84415348017
L6_74 V6 V74 -3.5994308984121204e-11
C6_74 V6 V74 3.0700850289590775e-21

R6_75 V6 V75 6930093.143691913
L6_75 V6 V75 1.9228553706399334e-11
C6_75 V6 V75 4.345051618924338e-21

R6_76 V6 V76 274368.7537972383
L6_76 V6 V76 -8.35240087128797e-12
C6_76 V6 V76 -5.368913769336892e-21

R6_77 V6 V77 2284925.8766471995
L6_77 V6 V77 -3.87608315830156e-11
C6_77 V6 V77 -2.917187148425833e-22

R6_78 V6 V78 98360.16844006021
L6_78 V6 V78 -2.210616843357265e-11
C6_78 V6 V78 -3.755968155130441e-21

R6_79 V6 V79 -425272.09227637056
L6_79 V6 V79 -6.8424894611286246e-12
C6_79 V6 V79 -1.8021636931969257e-20

R6_80 V6 V80 5859475.04787937
L6_80 V6 V80 9.406784197711225e-12
C6_80 V6 V80 1.3676110408710045e-20

R6_81 V6 V81 3356602.922018091
L6_81 V6 V81 8.661606339956834e-11
C6_81 V6 V81 7.081722425277742e-21

R6_82 V6 V82 58769.37453902046
L6_82 V6 V82 1.1774193174431827e-11
C6_82 V6 V82 7.943488357732381e-21

R6_83 V6 V83 -29888.660776283126
L6_83 V6 V83 1.389002349973839e-11
C6_83 V6 V83 1.3232967903894442e-20

R6_84 V6 V84 36942.766534901515
L6_84 V6 V84 -1.894133823175056e-11
C6_84 V6 V84 -6.059052690730031e-21

R6_85 V6 V85 163251.60977196932
L6_85 V6 V85 -1.0005546263521012e-11
C6_85 V6 V85 -1.1095855447513534e-20

R6_86 V6 V86 31511.050525473674
L6_86 V6 V86 -5.181899821571759e-10
C6_86 V6 V86 -4.9274884952532015e-21

R6_87 V6 V87 1099031.7512987137
L6_87 V6 V87 -9.222800541084118e-12
C6_87 V6 V87 -8.052373658232319e-21

R6_88 V6 V88 597046.1616447805
L6_88 V6 V88 1.1244684317423956e-09
C6_88 V6 V88 1.5711394839440274e-21

R6_89 V6 V89 135116.16246217652
L6_89 V6 V89 1.0723873775945671e-10
C6_89 V6 V89 8.438324348257936e-22

R6_90 V6 V90 -29707.60909235316
L6_90 V6 V90 6.372410472354634e-12
C6_90 V6 V90 1.989211686898449e-20

R6_91 V6 V91 -103016.83735791857
L6_91 V6 V91 1.3728077547103403e-11
C6_91 V6 V91 1.2132201993666229e-20

R6_92 V6 V92 -12644906.664358368
L6_92 V6 V92 2.0759892097933538e-11
C6_92 V6 V92 4.033783047723434e-21

R6_93 V6 V93 -124814.64989596547
L6_93 V6 V93 -1.9288745561097332e-11
C6_93 V6 V93 -4.256239077570975e-21

R6_94 V6 V94 22358.828254157135
L6_94 V6 V94 7.362369199145838e-11
C6_94 V6 V94 2.9905770480890125e-21

R6_95 V6 V95 -53172.39959226367
L6_95 V6 V95 2.423241398760357e-11
C6_95 V6 V95 6.051473705796475e-21

R6_96 V6 V96 -193847.42082110464
L6_96 V6 V96 2.5049009550888704e-11
C6_96 V6 V96 -3.5462599860052173e-22

R6_97 V6 V97 -55741.60749471209
L6_97 V6 V97 1.1940178217432845e-11
C6_97 V6 V97 8.306817607876813e-21

R6_98 V6 V98 -29905.00478137014
L6_98 V6 V98 1.2896942491601086e-11
C6_98 V6 V98 6.952423263505857e-21

R6_99 V6 V99 17152.887499563887
L6_99 V6 V99 -1.2784420325076435e-11
C6_99 V6 V99 -2.0444029707534366e-21

R6_100 V6 V100 131054.50940108046
L6_100 V6 V100 1.6462849000421846e-10
C6_100 V6 V100 5.469040655483335e-21

R6_101 V6 V101 74546.459676566
L6_101 V6 V101 3.2965016076375094e-11
C6_101 V6 V101 4.840496182042566e-22

R6_102 V6 V102 -57094.52009191547
L6_102 V6 V102 3.1521949181993893e-12
C6_102 V6 V102 3.7034026974455437e-20

R6_103 V6 V103 -115872.9299913934
L6_103 V6 V103 -5.44566339124764e-12
C6_103 V6 V103 -2.382580994245728e-20

R6_104 V6 V104 68366.87784512223
L6_104 V6 V104 -1.181517991008385e-10
C6_104 V6 V104 -1.9906143176285087e-21

R6_105 V6 V105 1059614.2910879331
L6_105 V6 V105 -7.288861995862878e-12
C6_105 V6 V105 -9.832564136003007e-21

R6_106 V6 V106 32599.909547295603
L6_106 V6 V106 4.948559297701947e-12
C6_106 V6 V106 2.3256324070222982e-20

R6_107 V6 V107 33891.79776861471
L6_107 V6 V107 3.882676037955582e-12
C6_107 V6 V107 3.349704888274505e-20

R6_108 V6 V108 -20857.283847598264
L6_108 V6 V108 -4.665965389781014e-12
C6_108 V6 V108 -2.0018160388276054e-20

R6_109 V6 V109 -232775.75475060983
L6_109 V6 V109 -9.225015936130503e-12
C6_109 V6 V109 -1.5540236004224496e-20

R6_110 V6 V110 -10662.206527794533
L6_110 V6 V110 -1.0891947861357e-11
C6_110 V6 V110 -1.5431661720535102e-20

R6_111 V6 V111 15822.128212804475
L6_111 V6 V111 -6.016564006623341e-12
C6_111 V6 V111 -1.2617503981459555e-20

R6_112 V6 V112 -17748.409080124773
L6_112 V6 V112 5.03265545143109e-12
C6_112 V6 V112 1.6027243211959112e-20

R6_113 V6 V113 -23265.70193296145
L6_113 V6 V113 1.0427017885313158e-11
C6_113 V6 V113 1.1054467226205236e-20

R6_114 V6 V114 -42016.36873089815
L6_114 V6 V114 9.928140851308034e-12
C6_114 V6 V114 5.35503876142985e-21

R6_115 V6 V115 -29008.56131790045
L6_115 V6 V115 7.48620840433063e-12
C6_115 V6 V115 2.094882165740499e-20

R6_116 V6 V116 38812.3879355556
L6_116 V6 V116 -7.617877078160774e-12
C6_116 V6 V116 -1.535128732804451e-20

R6_117 V6 V117 -18261.19942380572
L6_117 V6 V117 -1.6101590326632274e-11
C6_117 V6 V117 -1.4343293999275825e-20

R6_118 V6 V118 49531.03063362472
L6_118 V6 V118 -1.012399763069992e-11
C6_118 V6 V118 -1.1810923507517637e-20

R6_119 V6 V119 19513.48016683199
L6_119 V6 V119 -7.983958677988026e-12
C6_119 V6 V119 -9.588748870782264e-21

R6_120 V6 V120 -4155.710133161452
L6_120 V6 V120 9.280322721697414e-12
C6_120 V6 V120 -2.4257926062237937e-21

R6_121 V6 V121 -90931.72804868929
L6_121 V6 V121 4.6734761966324164e-11
C6_121 V6 V121 2.7380028620571756e-21

R6_122 V6 V122 -3205.4316523762486
L6_122 V6 V122 5.805963388158391e-12
C6_122 V6 V122 -1.0602860218292528e-21

R6_123 V6 V123 -15355.214092749453
L6_123 V6 V123 3.1428881747826807e-11
C6_123 V6 V123 -1.9360814066430086e-21

R6_124 V6 V124 61578.90451861479
L6_124 V6 V124 -2.7995811562910684e-11
C6_124 V6 V124 -1.8859748351699754e-21

R6_125 V6 V125 -13980.398426670325
L6_125 V6 V125 4.648157801977915e-11
C6_125 V6 V125 -3.747108360524082e-21

R6_126 V6 V126 2418.753020021475
L6_126 V6 V126 -4.332489516951325e-12
C6_126 V6 V126 2.797288282845244e-21

R6_127 V6 V127 -3189.357876701097
L6_127 V6 V127 5.09163106633867e-12
C6_127 V6 V127 1.4023790878097276e-21

R6_128 V6 V128 -36937.88929416062
L6_128 V6 V128 6.91359087221871e-11
C6_128 V6 V128 -9.418650146886576e-22

R6_129 V6 V129 -8555.337356149646
L6_129 V6 V129 1.5968003093321368e-11
C6_129 V6 V129 4.786643803084709e-22

R6_130 V6 V130 13157.519481637592
L6_130 V6 V130 -8.108590864002682e-12
C6_130 V6 V130 -7.296950190302448e-21

R6_131 V6 V131 9293.466727488541
L6_131 V6 V131 -8.603675169441611e-11
C6_131 V6 V131 6.046184103012433e-21

R6_132 V6 V132 12598.208887242201
L6_132 V6 V132 -1.996233561105141e-11
C6_132 V6 V132 -2.3921027931253843e-22

R6_133 V6 V133 52146.80777334516
L6_133 V6 V133 2.063831649857205e-11
C6_133 V6 V133 6.01352099277973e-21

R6_134 V6 V134 17421.998079154724
L6_134 V6 V134 -4.52655804611314e-11
C6_134 V6 V134 4.321272816265743e-22

R6_135 V6 V135 -4641.456635904884
L6_135 V6 V135 8.167300168295577e-12
C6_135 V6 V135 -3.1956517959482893e-21

R6_136 V6 V136 -157701.2449255253
L6_136 V6 V136 3.2607084642342603e-10
C6_136 V6 V136 -1.537147395510087e-22

R6_137 V6 V137 -45963.667516537775
L6_137 V6 V137 -4.312822168525741e-11
C6_137 V6 V137 -1.60519942207134e-22

R6_138 V6 V138 2893.437655780819
L6_138 V6 V138 -4.695118174466064e-12
C6_138 V6 V138 -1.4771053551542699e-21

R6_139 V6 V139 -2471.253422971517
L6_139 V6 V139 3.824435810616292e-12
C6_139 V6 V139 3.8870996077192076e-21

R6_140 V6 V140 10145.97348088649
L6_140 V6 V140 -1.0619101673344898e-11
C6_140 V6 V140 -1.6017187681126946e-21

R6_141 V6 V141 13716.692132204187
L6_141 V6 V141 -1.9712315467916392e-11
C6_141 V6 V141 -9.763892166891697e-22

R6_142 V6 V142 9804.302265432145
L6_142 V6 V142 -9.572516328324277e-12
C6_142 V6 V142 -4.874874424952951e-22

R6_143 V6 V143 7547.619681083487
L6_143 V6 V143 -1.1682235433620051e-11
C6_143 V6 V143 -3.810938352207933e-21

R6_144 V6 V144 -21809.27768638132
L6_144 V6 V144 1.6651515729816056e-11
C6_144 V6 V144 4.516285373617723e-21

R7_7 V7 0 -6872.122236299772
L7_7 V7 0 2.1774333483226157e-11
C7_7 V7 0 3.286471211197698e-20

R7_8 V7 V8 -16109452.947425468
L7_8 V7 V8 -4.4045249686092025e-09
C7_8 V7 V8 3.407377204194663e-22

R7_9 V7 V9 -994260.7654383436
L7_9 V7 V9 1.6096607675093097e-09
C7_9 V7 V9 -1.1365901957814053e-21

R7_10 V7 V10 -3009031.9518033406
L7_10 V7 V10 1.2436827682291853e-10
C7_10 V7 V10 -7.773273579458783e-22

R7_11 V7 V11 -902252.6046462466
L7_11 V7 V11 -1.2488698316616398e-10
C7_11 V7 V11 -3.9093654026672853e-22

R7_12 V7 V12 3392117.6614329545
L7_12 V7 V12 1.0941984509904736e-10
C7_12 V7 V12 -8.326456767861883e-22

R7_13 V7 V13 1963330.6602243674
L7_13 V7 V13 1.988955543154934e-10
C7_13 V7 V13 -2.9028429575363555e-22

R7_14 V7 V14 2975527.1365161426
L7_14 V7 V14 -8.087346248832908e-11
C7_14 V7 V14 1.113976427211883e-21

R7_15 V7 V15 -736002.7930382423
L7_15 V7 V15 -3.0446359699312275e-10
C7_15 V7 V15 4.873243339618168e-22

R7_16 V7 V16 1171866.133987327
L7_16 V7 V16 -3.6721207549480275e-10
C7_16 V7 V16 3.622695157500106e-22

R7_17 V7 V17 532249.8413450432
L7_17 V7 V17 -3.342092930463255e-10
C7_17 V7 V17 6.349684499158122e-22

R7_18 V7 V18 3378229.499234503
L7_18 V7 V18 3.980466294149521e-10
C7_18 V7 V18 -3.2446923750536223e-22

R7_19 V7 V19 -137321.44255080723
L7_19 V7 V19 6.222009540016689e-11
C7_19 V7 V19 -2.5640959637819822e-21

R7_20 V7 V20 3211514.0931152473
L7_20 V7 V20 -2.7086931863614538e-09
C7_20 V7 V20 2.303203178391437e-22

R7_21 V7 V21 -815972.5857579486
L7_21 V7 V21 1.759614303810972e-10
C7_21 V7 V21 -1.3810181570670914e-21

R7_22 V7 V22 -1629203.3344045272
L7_22 V7 V22 3.242643903522539e-11
C7_22 V7 V22 -7.860791666660886e-22

R7_23 V7 V23 269162.4528020847
L7_23 V7 V23 -1.7597246956489372e-11
C7_23 V7 V23 2.6018732053614872e-21

R7_24 V7 V24 4632437.64616598
L7_24 V7 V24 -3.7242213858288013e-10
C7_24 V7 V24 -1.2811541790353575e-23

R7_25 V7 V25 519157.9378959867
L7_25 V7 V25 2.320255684317352e-10
C7_25 V7 V25 -4.75649202908608e-22

R7_26 V7 V26 -37995383.58975987
L7_26 V7 V26 4.455950384579855e-11
C7_26 V7 V26 -1.265884820728642e-21

R7_27 V7 V27 -225880.64314305974
L7_27 V7 V27 -1.2885716597365382e-10
C7_27 V7 V27 7.07877916362168e-22

R7_28 V7 V28 -12309837.178794362
L7_28 V7 V28 -9.694018272633836e-10
C7_28 V7 V28 4.112888174921294e-23

R7_29 V7 V29 818040.457356515
L7_29 V7 V29 1.386798754654841e-10
C7_29 V7 V29 3.426033980295179e-21

R7_30 V7 V30 -744121.5267540693
L7_30 V7 V30 4.026732479848282e-11
C7_30 V7 V30 1.9382969959778446e-21

R7_31 V7 V31 -1153353.7451835927
L7_31 V7 V31 -3.757239116689359e-11
C7_31 V7 V31 -7.036193167942266e-21

R7_32 V7 V32 816168.8822863541
L7_32 V7 V32 -7.616134741849861e-10
C7_32 V7 V32 4.927309718535706e-22

R7_33 V7 V33 -221909.72193745108
L7_33 V7 V33 -2.363263464237067e-10
C7_33 V7 V33 -6.927588853525061e-21

R7_34 V7 V34 278316.81370309775
L7_34 V7 V34 -1.2105881885672437e-10
C7_34 V7 V34 -5.936861586938442e-23

R7_35 V7 V35 -51248.018203713225
L7_35 V7 V35 3.5552279269557495e-11
C7_35 V7 V35 3.825041905661483e-21

R7_36 V7 V36 548018.8230738005
L7_36 V7 V36 -3.1152929631487123e-10
C7_36 V7 V36 9.699547349767616e-25

R7_37 V7 V37 45810.67133782604
L7_37 V7 V37 -9.113287219167967e-11
C7_37 V7 V37 6.810248845985698e-21

R7_38 V7 V38 -5416065.175339236
L7_38 V7 V38 4.091714388428566e-11
C7_38 V7 V38 6.6652567167081876e-21

R7_39 V7 V39 -2032045.4172455308
L7_39 V7 V39 -7.389848305600647e-10
C7_39 V7 V39 -4.7173496207017235e-21

R7_40 V7 V40 -384028.651980721
L7_40 V7 V40 1.2712333378790132e-10
C7_40 V7 V40 1.6528614599903358e-21

R7_41 V7 V41 581993.416294007
L7_41 V7 V41 -2.2403774213706624e-11
C7_41 V7 V41 -2.577433367981328e-20

R7_42 V7 V42 -177872.91797735202
L7_42 V7 V42 -1.1357446548461287e-11
C7_42 V7 V42 -3.531168696134048e-20

R7_43 V7 V43 -147276.306235123
L7_43 V7 V43 9.910629740880093e-11
C7_43 V7 V43 4.117784672487961e-21

R7_44 V7 V44 1177531.0668937312
L7_44 V7 V44 -3.6173835437529605e-11
C7_44 V7 V44 -1.5015118389943708e-20

R7_45 V7 V45 29480.18415279399
L7_45 V7 V45 -2.993491199835325e-11
C7_45 V7 V45 -2.541490559297167e-21

R7_46 V7 V46 69606.47591748543
L7_46 V7 V46 2.0162914641883092e-11
C7_46 V7 V46 3.850270731552419e-20

R7_47 V7 V47 -30448.41524535383
L7_47 V7 V47 3.805525402307545e-11
C7_47 V7 V47 7.090202468349993e-21

R7_48 V7 V48 60202.203019694716
L7_48 V7 V48 1.2771579459488326e-10
C7_48 V7 V48 6.189539098430381e-21

R7_49 V7 V49 23725.065635969942
L7_49 V7 V49 2.931135647773406e-10
C7_49 V7 V49 5.447465470713298e-21

R7_50 V7 V50 -23586.960983719946
L7_50 V7 V50 -3.047638320327636e-10
C7_50 V7 V50 -1.669145739809829e-20

R7_51 V7 V51 -421986.79075445223
L7_51 V7 V51 8.386765398001164e-11
C7_51 V7 V51 9.606768991488968e-21

R7_52 V7 V52 -162465.94720070888
L7_52 V7 V52 -7.890318806378223e-11
C7_52 V7 V52 -1.3343451310019014e-20

R7_53 V7 V53 -446842.00609163597
L7_53 V7 V53 1.273992806084766e-10
C7_53 V7 V53 -4.183367195216749e-21

R7_54 V7 V54 501542.82819905743
L7_54 V7 V54 -1.867912525949439e-10
C7_54 V7 V54 -3.489267174084538e-21

R7_55 V7 V55 32513.727232846428
L7_55 V7 V55 7.054776161339371e-11
C7_55 V7 V55 5.3493765391510005e-21

R7_56 V7 V56 500995.2066029979
L7_56 V7 V56 1.3299297567434673e-10
C7_56 V7 V56 1.5031760743401686e-21

R7_57 V7 V57 40825.76974022743
L7_57 V7 V57 -2.3323505474234627e-11
C7_57 V7 V57 2.796735555595591e-21

R7_58 V7 V58 17116.69397536545
L7_58 V7 V58 -1.5045173042466808e-11
C7_58 V7 V58 4.350632026320946e-21

R7_59 V7 V59 -17950.949530831756
L7_59 V7 V59 3.328911708227523e-11
C7_59 V7 V59 2.942183467212818e-21

R7_60 V7 V60 444903.90933340404
L7_60 V7 V60 -7.629629568485322e-09
C7_60 V7 V60 1.513845317184609e-21

R7_61 V7 V61 -841801.0374857618
L7_61 V7 V61 6.097161101312313e-11
C7_61 V7 V61 -8.143728106947479e-21

R7_62 V7 V62 -23875.29690479606
L7_62 V7 V62 1.036550787525756e-10
C7_62 V7 V62 -1.1091440318836341e-20

R7_63 V7 V63 51508.59319688509
L7_63 V7 V63 -7.142353851191682e-11
C7_63 V7 V63 6.155905873949205e-21

R7_64 V7 V64 196593.85220481385
L7_64 V7 V64 5.095386928132418e-11
C7_64 V7 V64 2.1477297676863575e-21

R7_65 V7 V65 48843.158827425636
L7_65 V7 V65 1.7084510289553418e-10
C7_65 V7 V65 -3.3535816878355402e-21

R7_66 V7 V66 23779.145268262906
L7_66 V7 V66 -6.550541185890962e-11
C7_66 V7 V66 -1.8669559960370945e-21

R7_67 V7 V67 -30598.504754595357
L7_67 V7 V67 -1.5577091011633907e-10
C7_67 V7 V67 1.6373574555149344e-21

R7_68 V7 V68 425700.4699847109
L7_68 V7 V68 -9.070557814611722e-11
C7_68 V7 V68 7.537421875881469e-22

R7_69 V7 V69 1384189.9855356298
L7_69 V7 V69 -7.651759736909387e-11
C7_69 V7 V69 2.7379122079539696e-22

R7_70 V7 V70 -116990.22599173237
L7_70 V7 V70 2.1677133609193827e-10
C7_70 V7 V70 1.321048223217954e-21

R7_71 V7 V71 33080.92241107257
L7_71 V7 V71 2.385237539744751e-11
C7_71 V7 V71 9.618106385199979e-22

R7_72 V7 V72 -33196.87057845426
L7_72 V7 V72 -3.72146770270598e-11
C7_72 V7 V72 -7.378533140807139e-22

R7_73 V7 V73 -64876.70107272671
L7_73 V7 V73 -5.945261627426726e-11
C7_73 V7 V73 -2.1152396676684084e-22

R7_74 V7 V74 -109306.79270163148
L7_74 V7 V74 7.439762236922255e-11
C7_74 V7 V74 2.9234837830929326e-21

R7_75 V7 V75 109131.61114919338
L7_75 V7 V75 -1.5052279087134175e-10
C7_75 V7 V75 -3.185028658984086e-22

R7_76 V7 V76 127786.90029994644
L7_76 V7 V76 3.531120368892674e-11
C7_76 V7 V76 2.577298996450231e-22

R7_77 V7 V77 371408.6001620291
L7_77 V7 V77 1.6219005896151408e-10
C7_77 V7 V77 -2.3861461624606597e-21

R7_78 V7 V78 -166884.58842626022
L7_78 V7 V78 -5.0464768507020103e-11
C7_78 V7 V78 -3.2552279868252428e-21

R7_79 V7 V79 -474722.2524871733
L7_79 V7 V79 2.726710971381538e-11
C7_79 V7 V79 4.991171511053463e-21

R7_80 V7 V80 -123374.94757836072
L7_80 V7 V80 -2.503969491735318e-11
C7_80 V7 V80 -8.622255475689591e-21

R7_81 V7 V81 938735.5348229271
L7_81 V7 V81 2.1437880080715536e-10
C7_81 V7 V81 5.356699585212411e-21

R7_82 V7 V82 356923.44488182326
L7_82 V7 V82 1.2621886619244873e-11
C7_82 V7 V82 9.973183934882795e-21

R7_83 V7 V83 101435.46272112196
L7_83 V7 V83 2.3274749046354047e-11
C7_83 V7 V83 5.388124450538454e-21

R7_84 V7 V84 -130922.07328855337
L7_84 V7 V84 4.76710155584027e-11
C7_84 V7 V84 5.784213954866899e-21

R7_85 V7 V85 -221719.31554352396
L7_85 V7 V85 1.338452689799417e-10
C7_85 V7 V85 3.852673518846957e-21

R7_86 V7 V86 -93792.49591070044
L7_86 V7 V86 -2.580885231494283e-11
C7_86 V7 V86 -3.2407798909374298e-21

R7_87 V7 V87 -9129707.889539897
L7_87 V7 V87 -1.3171178081438363e-10
C7_87 V7 V87 -1.0087712557709469e-21

R7_88 V7 V88 -474197.6109762409
L7_88 V7 V88 -7.737134046180828e-11
C7_88 V7 V88 -1.125255962658666e-21

R7_89 V7 V89 -422091.1210721385
L7_89 V7 V89 2.849893865714535e-10
C7_89 V7 V89 -2.8035505209936834e-21

R7_90 V7 V90 107469.67799162898
L7_90 V7 V90 -1.9188619640891233e-11
C7_90 V7 V90 -6.900497853676639e-21

R7_91 V7 V91 134439.96349531593
L7_91 V7 V91 1.2093266577309577e-11
C7_91 V7 V91 1.2875040663260253e-20

R7_92 V7 V92 1787493.3453119865
L7_92 V7 V92 1.12570009465591e-10
C7_92 V7 V92 -2.675122611470714e-21

R7_93 V7 V93 -95509.88496204215
L7_93 V7 V93 -2.3936357550936917e-09
C7_93 V7 V93 -1.4608703145679528e-21

R7_94 V7 V94 -57635.63529514622
L7_94 V7 V94 -3.4985842183574814e-11
C7_94 V7 V94 -3.016845963682151e-21

R7_95 V7 V95 170869.49570571654
L7_95 V7 V95 2.3290992582843472e-11
C7_95 V7 V95 5.749570625251138e-21

R7_96 V7 V96 -281434.4561829367
L7_96 V7 V96 -4.2988208262631296e-11
C7_96 V7 V96 -4.682226663226604e-21

R7_97 V7 V97 182255.74788751002
L7_97 V7 V97 -1.5200222672810728e-11
C7_97 V7 V97 -5.1961918058702056e-21

R7_98 V7 V98 71592.85374570474
L7_98 V7 V98 -8.137528984494663e-09
C7_98 V7 V98 -4.853992427305911e-22

R7_99 V7 V99 -60201.6520036921
L7_99 V7 V99 4.806245757084245e-11
C7_99 V7 V99 7.608895720256063e-22

R7_100 V7 V100 3014299.7339453097
L7_100 V7 V100 -1.2379180912045063e-10
C7_100 V7 V100 8.448538113502596e-22

R7_101 V7 V101 -108754.78309654196
L7_101 V7 V101 8.240615191023721e-11
C7_101 V7 V101 -2.546385875644945e-21

R7_102 V7 V102 148879.7287022845
L7_102 V7 V102 -1.2707773628009951e-11
C7_102 V7 V102 -1.1189489727058612e-20

R7_103 V7 V103 174958.59758215107
L7_103 V7 V103 1.735245745604996e-11
C7_103 V7 V103 8.883662757021751e-21

R7_104 V7 V104 -166184.57704514317
L7_104 V7 V104 -3.710387569792469e-11
C7_104 V7 V104 -6.738862168056957e-21

R7_105 V7 V105 -394331.8534450448
L7_105 V7 V105 -2.985972866400976e-10
C7_105 V7 V105 -1.145903101333574e-21

R7_106 V7 V106 -134969.6641756392
L7_106 V7 V106 2.8473906437264195e-11
C7_106 V7 V106 3.515572891104488e-21

R7_107 V7 V107 -139035.9008991732
L7_107 V7 V107 -1.8008293233088014e-11
C7_107 V7 V107 -6.675433629961413e-21

R7_108 V7 V108 47715.52985902778
L7_108 V7 V108 1.9681134959604486e-11
C7_108 V7 V108 1.2422738951495617e-20

R7_109 V7 V109 168710.1778733273
L7_109 V7 V109 7.483657411777028e-11
C7_109 V7 V109 -8.278927481949354e-23

R7_110 V7 V110 36683.41862136241
L7_110 V7 V110 -2.528145683060147e-11
C7_110 V7 V110 -5.3298354265316776e-21

R7_111 V7 V111 -92699.33660098517
L7_111 V7 V111 4.681333666252454e-11
C7_111 V7 V111 1.4815767841643505e-21

R7_112 V7 V112 36845.93863689642
L7_112 V7 V112 -2.1765179668240222e-11
C7_112 V7 V112 -6.667905945465855e-21

R7_113 V7 V113 91805.33102452703
L7_113 V7 V113 -8.771246730715607e-11
C7_113 V7 V113 4.373884328175471e-22

R7_114 V7 V114 94047.32052021065
L7_114 V7 V114 1.2376415616361414e-10
C7_114 V7 V114 3.834786106011827e-21

R7_115 V7 V115 102195.59930451633
L7_115 V7 V115 -3.6189347782351034e-11
C7_115 V7 V115 -5.2718747147254695e-21

R7_116 V7 V116 -132612.37853853204
L7_116 V7 V116 3.3857399885065514e-11
C7_116 V7 V116 8.030186406793379e-21

R7_117 V7 V117 70433.53893739675
L7_117 V7 V117 2.3528300698533535e-10
C7_117 V7 V117 3.2618998593725477e-21

R7_118 V7 V118 -157827.97654345387
L7_118 V7 V118 -1.0209177353698657e-10
C7_118 V7 V118 -4.212220125236594e-21

R7_119 V7 V119 -82416.68812727567
L7_119 V7 V119 -1.2209572909995416e-10
C7_119 V7 V119 -2.146970551998551e-21

R7_120 V7 V120 16898.24216342345
L7_120 V7 V120 -4.007054433039441e-11
C7_120 V7 V120 1.7094590105981995e-21

R7_121 V7 V121 45320.77383625221
L7_121 V7 V121 -1.0507497308833504e-10
C7_121 V7 V121 1.5744093492087705e-21

R7_122 V7 V122 9263.814917759964
L7_122 V7 V122 -1.5556278563363453e-11
C7_122 V7 V122 -1.0110590625467491e-22

R7_123 V7 V123 37936.69444173085
L7_123 V7 V123 -5.914086188421155e-11
C7_123 V7 V123 -2.6000742894839816e-21

R7_124 V7 V124 113963.19815244107
L7_124 V7 V124 -4.542348964021835e-09
C7_124 V7 V124 -5.368105646893511e-23

R7_125 V7 V125 4773984.963280387
L7_125 V7 V125 1.6329060517788014e-10
C7_125 V7 V125 8.833636932959718e-22

R7_126 V7 V126 -7853.473147587993
L7_126 V7 V126 1.3277272839022859e-11
C7_126 V7 V126 -5.397367102022194e-22

R7_127 V7 V127 11187.996148302647
L7_127 V7 V127 -1.917021437100968e-11
C7_127 V7 V127 -4.868614256914507e-22

R7_128 V7 V128 -368054.2570519834
L7_128 V7 V128 1.7817363379447365e-10
C7_128 V7 V128 -1.5639596640411196e-21

R7_129 V7 V129 22011.421613811915
L7_129 V7 V129 -5.924527173729647e-11
C7_129 V7 V129 -5.748741730917361e-22

R7_130 V7 V130 -29511.066188996174
L7_130 V7 V130 2.855507173181479e-11
C7_130 V7 V130 1.3067842166392185e-21

R7_131 V7 V131 -22284.781912468006
L7_131 V7 V131 9.727266204471711e-11
C7_131 V7 V131 -1.5892123359216155e-21

R7_132 V7 V132 -43324.73581014188
L7_132 V7 V132 4.427296470470372e-11
C7_132 V7 V132 1.7177782972230566e-21

R7_133 V7 V133 -96742.53916341435
L7_133 V7 V133 5.450660355345182e-11
C7_133 V7 V133 2.473151203736658e-21

R7_134 V7 V134 -55705.045757281165
L7_134 V7 V134 7.494186780620028e-11
C7_134 V7 V134 -1.818547567709213e-21

R7_135 V7 V135 15807.255752473788
L7_135 V7 V135 -2.7418871394103732e-11
C7_135 V7 V135 9.969854381091338e-22

R7_136 V7 V136 -128155.15034604029
L7_136 V7 V136 1.2982031658806744e-09
C7_136 V7 V136 3.8266350297463536e-22

R7_137 V7 V137 -298866.8464898969
L7_137 V7 V137 1.3531802687077695e-10
C7_137 V7 V137 -8.303424664012147e-22

R7_138 V7 V138 -8929.660253649296
L7_138 V7 V138 1.362626129046779e-11
C7_138 V7 V138 3.0911046091700035e-23

R7_139 V7 V139 8779.869892316663
L7_139 V7 V139 -1.4283184799228888e-11
C7_139 V7 V139 -3.0025095749977424e-22

R7_140 V7 V140 -31139.52607787607
L7_140 V7 V140 3.142540974080192e-11
C7_140 V7 V140 1.626857101905856e-21

R7_141 V7 V141 -61002.131132061186
L7_141 V7 V141 7.90973801819971e-11
C7_141 V7 V141 -3.183256342387678e-22

R7_142 V7 V142 -22629.52528089517
L7_142 V7 V142 3.7537761358504815e-11
C7_142 V7 V142 -1.6662357406275034e-22

R7_143 V7 V143 -25209.907807995965
L7_143 V7 V143 4.2523663737875506e-11
C7_143 V7 V143 8.806357920498471e-22

R7_144 V7 V144 55646.70223526638
L7_144 V7 V144 -4.8370663902092065e-11
C7_144 V7 V144 -1.0280516563899402e-21

R8_8 V8 0 1650.8112016107175
L8_8 V8 0 -2.1249471933777578e-12
C8_8 V8 0 -7.38656517681341e-20

R8_9 V8 V9 -2076899.844905396
L8_9 V8 V9 -9.749003069464712e-11
C8_9 V8 V9 4.126935841695693e-22

R8_10 V8 V10 444615.06512890273
L8_10 V8 V10 3.037512680869789e-10
C8_10 V8 V10 -8.414189984494337e-22

R8_11 V8 V11 440038.9901083219
L8_11 V8 V11 6.655063849481068e-11
C8_11 V8 V11 -4.857918364869378e-22

R8_12 V8 V12 -811874.4344137333
L8_12 V8 V12 -1.1421884868424972e-11
C8_12 V8 V12 5.037595020151696e-21

R8_13 V8 V13 -1291438.2927572245
L8_13 V8 V13 2.916806107360469e-11
C8_13 V8 V13 -1.697140026381009e-21

R8_14 V8 V14 -347689.44167592033
L8_14 V8 V14 -1.976956483659689e-11
C8_14 V8 V14 1.288208299595974e-21

R8_15 V8 V15 -506874.32911461376
L8_15 V8 V15 -2.407360732429114e-11
C8_15 V8 V15 1.2479667422832626e-21

R8_16 V8 V16 -220322.0652474704
L8_16 V8 V16 -3.443565015209514e-11
C8_16 V8 V16 -1.6123191451171175e-22

R8_17 V8 V17 -204088.22221078892
L8_17 V8 V17 -8.299838212846262e-11
C8_17 V8 V17 -6.237018495559951e-22

R8_18 V8 V18 1123399.542395622
L8_18 V8 V18 2.4942967518839797e-10
C8_18 V8 V18 7.660732568162388e-22

R8_19 V8 V19 -248748.85916453935
L8_19 V8 V19 -3.0444534598171316e-10
C8_19 V8 V19 4.99889533357954e-22

R8_20 V8 V20 -56640.8882630768
L8_20 V8 V20 1.3863395646168986e-11
C8_20 V8 V20 -1.0871404986437149e-20

R8_21 V8 V21 358407.5851547658
L8_21 V8 V21 -1.0055891682916121e-10
C8_21 V8 V21 9.091628107002316e-22

R8_22 V8 V22 -937049.457907178
L8_22 V8 V22 -9.050228801557116e-10
C8_22 V8 V22 -6.145345472602184e-22

R8_23 V8 V23 -576748.4892508158
L8_23 V8 V23 4.0885673059541504e-11
C8_23 V8 V23 -1.7303823924217338e-21

R8_24 V8 V24 283121.40714875667
L8_24 V8 V24 -7.891650364030228e-12
C8_24 V8 V24 5.118668699164949e-21

R8_25 V8 V25 -468523.78781950666
L8_25 V8 V25 -1.1513639754850658e-10
C8_25 V8 V25 -1.0921117817721394e-21

R8_26 V8 V26 536874.6990580817
L8_26 V8 V26 7.684497418001625e-11
C8_26 V8 V26 -2.0563606092356416e-21

R8_27 V8 V27 237511.17929234155
L8_27 V8 V27 3.576055378516151e-10
C8_27 V8 V27 -1.980305170512541e-21

R8_28 V8 V28 -77251.91701169408
L8_28 V8 V28 -1.1068470118877637e-11
C8_28 V8 V28 2.218818026555192e-23

R8_29 V8 V29 440178.2616049681
L8_29 V8 V29 9.562048849219727e-11
C8_29 V8 V29 -6.223979447113205e-22

R8_30 V8 V30 -3521316.854558
L8_30 V8 V30 5.727292932816414e-11
C8_30 V8 V30 1.360712301824391e-21

R8_31 V8 V31 180761.47495027503
L8_31 V8 V31 6.350831043096537e-11
C8_31 V8 V31 6.0166664602161565e-21

R8_32 V8 V32 37994.95009447567
L8_32 V8 V32 -1.3335950418920252e-11
C8_32 V8 V32 -1.1680131764592813e-20

R8_33 V8 V33 -171681.50856991037
L8_33 V8 V33 -1.572671790277124e-10
C8_33 V8 V33 1.9950668195874993e-21

R8_34 V8 V34 260191.79944795917
L8_34 V8 V34 -1.389007734372577e-10
C8_34 V8 V34 2.0985789234763985e-21

R8_35 V8 V35 396397.6600937132
L8_35 V8 V35 -2.16902690844391e-11
C8_35 V8 V35 -3.1096549019195755e-21

R8_36 V8 V36 -16321.273297070207
L8_36 V8 V36 4.081276687305451e-11
C8_36 V8 V36 4.486422315292144e-21

R8_37 V8 V37 -141263.27659202914
L8_37 V8 V37 -9.171885180513437e-11
C8_37 V8 V37 4.791761692019686e-22

R8_38 V8 V38 6051073.42995887
L8_38 V8 V38 -1.1918349070292222e-10
C8_38 V8 V38 6.61306834021032e-21

R8_39 V8 V39 -231998.72762686483
L8_39 V8 V39 -2.0527734974719605e-10
C8_39 V8 V39 8.437950909464026e-21

R8_40 V8 V40 -64419.71146668557
L8_40 V8 V40 -1.9169783389724573e-11
C8_40 V8 V40 -6.531801513966538e-20

R8_41 V8 V41 -67607.93771540346
L8_41 V8 V41 1.1280285398283106e-11
C8_41 V8 V41 1.6811490256798934e-20

R8_42 V8 V42 1431553.6542070562
L8_42 V8 V42 2.5542422852110236e-11
C8_42 V8 V42 -7.386990578737206e-21

R8_43 V8 V43 -346968.434204263
L8_43 V8 V43 3.500144889885696e-11
C8_43 V8 V43 -9.471649129807977e-23

R8_44 V8 V44 -52650.913244579395
L8_44 V8 V44 4.5292159803717215e-12
C8_44 V8 V44 1.1662304938723573e-19

R8_45 V8 V45 -283853.8470180034
L8_45 V8 V45 -1.5680098685526882e-11
C8_45 V8 V45 -2.958051428299705e-20

R8_46 V8 V46 144123.65956010416
L8_46 V8 V46 2.775504559116291e-11
C8_46 V8 V46 1.2817280218744134e-20

R8_47 V8 V47 -28604.599073962563
L8_47 V8 V47 1.2627151179602216e-10
C8_47 V8 V47 -7.149777322884613e-21

R8_48 V8 V48 -8298.786239503816
L8_48 V8 V48 -6.999893125742868e-11
C8_48 V8 V48 -3.092060999600937e-20

R8_49 V8 V49 -468272.9386013031
L8_49 V8 V49 8.092329684489041e-11
C8_49 V8 V49 2.965861572379671e-21

R8_50 V8 V50 334579.1824836636
L8_50 V8 V50 8.09713487292471e-11
C8_50 V8 V50 5.713501327918731e-21

R8_51 V8 V51 -237955.9269666473
L8_51 V8 V51 3.211419339253652e-10
C8_51 V8 V51 1.6261458420071655e-21

R8_52 V8 V52 27746.262967680155
L8_52 V8 V52 2.1544557614795374e-11
C8_52 V8 V52 1.6666960144739884e-20

R8_53 V8 V53 -18211.087860002794
L8_53 V8 V53 -2.1287033714278832e-11
C8_53 V8 V53 -2.3636499595333064e-20

R8_54 V8 V54 -37360.75397581315
L8_54 V8 V54 -8.533199989880882e-11
C8_54 V8 V54 -1.1353429267611464e-20

R8_55 V8 V55 -76056.92128217274
L8_55 V8 V55 3.0538668633914954e-11
C8_55 V8 V55 -2.1617017541479383e-21

R8_56 V8 V56 9778.852229428772
L8_56 V8 V56 7.380962163042894e-12
C8_56 V8 V56 5.31489082960292e-20

R8_57 V8 V57 -13730.866616661737
L8_57 V8 V57 1.7329706637966648e-11
C8_57 V8 V57 2.4045829431295093e-21

R8_58 V8 V58 38031.36157175519
L8_58 V8 V58 -2.1777472485923276e-11
C8_58 V8 V58 -5.457125202981445e-21

R8_59 V8 V59 94334.24845027241
L8_59 V8 V59 -5.147188441836812e-11
C8_59 V8 V59 -2.1896580837428745e-21

R8_60 V8 V60 -3767.9445113696993
L8_60 V8 V60 4.8367322123541e-12
C8_60 V8 V60 -3.3898164354460645e-21

R8_61 V8 V61 29941.016789349982
L8_61 V8 V61 -2.453742908853346e-11
C8_61 V8 V61 -2.7941500717045297e-21

R8_62 V8 V62 -119355.6987763383
L8_62 V8 V62 5.211568278541507e-11
C8_62 V8 V62 3.2057966094870078e-21

R8_63 V8 V63 201717.1925801302
L8_63 V8 V63 1.8073283934556912e-11
C8_63 V8 V63 6.39753048401867e-21

R8_64 V8 V64 -436722.8667941061
L8_64 V8 V64 -1.2998807305745178e-11
C8_64 V8 V64 2.0889468698095788e-20

R8_65 V8 V65 -20065.110496965634
L8_65 V8 V65 3.712537716330648e-11
C8_65 V8 V65 1.1046811519563713e-21

R8_66 V8 V66 -21264.491196264185
L8_66 V8 V66 -1.026369182217188e-11
C8_66 V8 V66 1.2868018082053371e-21

R8_67 V8 V67 -232666.03726797647
L8_67 V8 V67 6.684633824491298e-11
C8_67 V8 V67 5.783646717322974e-21

R8_68 V8 V68 -15645.556636241075
L8_68 V8 V68 7.1940856285669195e-12
C8_68 V8 V68 2.506208283914742e-21

R8_69 V8 V69 24727.411328853937
L8_69 V8 V69 -1.1677145271238123e-11
C8_69 V8 V69 -1.0504678983647205e-20

R8_70 V8 V70 -211350.7528995445
L8_70 V8 V70 -2.7636590322196862e-11
C8_70 V8 V70 -5.83374294190947e-21

R8_71 V8 V71 -71964.78626451132
L8_71 V8 V71 -3.50881965600163e-10
C8_71 V8 V71 -1.8304368332453956e-21

R8_72 V8 V72 31957.99953311039
L8_72 V8 V72 -1.6437969173282796e-10
C8_72 V8 V72 3.0004680022153514e-21

R8_73 V8 V73 -822532.9793237209
L8_73 V8 V73 -4.953586747158659e-11
C8_73 V8 V73 -1.1159970387816564e-20

R8_74 V8 V74 53951.4510431169
L8_74 V8 V74 -5.5117706050539585e-11
C8_74 V8 V74 -4.733008312971603e-21

R8_75 V8 V75 -229327.9148975548
L8_75 V8 V75 4.5933652527410725e-11
C8_75 V8 V75 9.483424432884956e-21

R8_76 V8 V76 -97616.70030566286
L8_76 V8 V76 -1.3124100177245702e-11
C8_76 V8 V76 -7.080877938852084e-21

R8_77 V8 V77 65365.715185518195
L8_77 V8 V77 1.4948747754851492e-11
C8_77 V8 V77 1.2228413182903815e-20

R8_78 V8 V78 15805137.757325465
L8_78 V8 V78 -2.637987449789389e-11
C8_78 V8 V78 -3.068810655882826e-21

R8_79 V8 V79 152975.02914090862
L8_79 V8 V79 -2.1552474386967465e-11
C8_79 V8 V79 -1.0373853619274482e-20

R8_80 V8 V80 63319.72922838336
L8_80 V8 V80 5.690383721156429e-12
C8_80 V8 V80 3.536512770885832e-20

R8_81 V8 V81 -34703.69458902581
L8_81 V8 V81 -3.1934959255158628e-12
C8_81 V8 V81 -6.088914261089106e-20

R8_82 V8 V82 -146836.08028734257
L8_82 V8 V82 1.144060520192028e-11
C8_82 V8 V82 1.8171057297887545e-21

R8_83 V8 V83 156685.42055971833
L8_83 V8 V83 5.226989537564244e-12
C8_83 V8 V83 2.893395869375289e-20

R8_84 V8 V84 92174.44833518553
L8_84 V8 V84 3.598264028033025e-11
C8_84 V8 V84 4.6467900977858074e-21

R8_85 V8 V85 345606.71090629837
L8_85 V8 V85 -1.2215057759422084e-11
C8_85 V8 V85 -9.372704659280669e-21

R8_86 V8 V86 145647.12952467677
L8_86 V8 V86 -2.6427488713799124e-11
C8_86 V8 V86 8.575917385220803e-21

R8_87 V8 V87 -209173.69647467244
L8_87 V8 V87 -1.0122142412391486e-11
C8_87 V8 V87 -8.983099202422732e-21

R8_88 V8 V88 -220831.72810181874
L8_88 V8 V88 -1.3504181933864809e-11
C8_88 V8 V88 -1.3445881788268969e-20

R8_89 V8 V89 1769953.8777679105
L8_89 V8 V89 1.3663285122994132e-11
C8_89 V8 V89 8.696906686774885e-21

R8_90 V8 V90 -910455.4194322503
L8_90 V8 V90 5.2202167011886594e-11
C8_90 V8 V90 7.745829860079218e-21

R8_91 V8 V91 -331598.03151334653
L8_91 V8 V91 1.232151815897317e-10
C8_91 V8 V91 -1.3229893908277096e-20

R8_92 V8 V92 51795.02599913019
L8_92 V8 V92 3.478985221018479e-12
C8_92 V8 V92 5.778731134088437e-20

R8_93 V8 V93 137441.60389354877
L8_93 V8 V93 -2.1436546185129702e-11
C8_93 V8 V93 -6.037615440596411e-21

R8_94 V8 V94 -262156.6086090543
L8_94 V8 V94 -7.575179712968937e-12
C8_94 V8 V94 -2.335692160887817e-20

R8_95 V8 V95 -1008664.7986005896
L8_95 V8 V95 3.3939984880981995e-11
C8_95 V8 V95 -1.1057635692891844e-21

R8_96 V8 V96 31942.886224652317
L8_96 V8 V96 3.0828142255790166e-12
C8_96 V8 V96 6.421020901960336e-20

R8_97 V8 V97 -576034.5245262218
L8_97 V8 V97 -1.1986737236568916e-11
C8_97 V8 V97 -1.3002963967448891e-20

R8_98 V8 V98 406696.8797520272
L8_98 V8 V98 7.09465805571547e-12
C8_98 V8 V98 1.820231245384402e-20

R8_99 V8 V99 -652510.9458049074
L8_99 V8 V99 -2.4584419077967798e-11
C8_99 V8 V99 -8.806918493414989e-21

R8_100 V8 V100 -142856.93525921047
L8_100 V8 V100 -9.21200837556695e-12
C8_100 V8 V100 -2.4811911108161093e-20

R8_101 V8 V101 574181.0447719148
L8_101 V8 V101 7.626571716232531e-12
C8_101 V8 V101 1.517036236654703e-20

R8_102 V8 V102 95677.20374605194
L8_102 V8 V102 1.2193508889540093e-11
C8_102 V8 V102 8.660476645558073e-21

R8_103 V8 V103 218018.34718691002
L8_103 V8 V103 -2.5734103260472165e-11
C8_103 V8 V103 -8.340734952882235e-21

R8_104 V8 V104 65316.2208982283
L8_104 V8 V104 5.331660265156866e-12
C8_104 V8 V104 5.466124905611005e-20

R8_105 V8 V105 -83170.4555424008
L8_105 V8 V105 -6.65605731731993e-12
C8_105 V8 V105 -2.963968538990521e-20

R8_106 V8 V106 88659.33371002163
L8_106 V8 V106 6.104186171349781e-12
C8_106 V8 V106 2.278324985778466e-20

R8_107 V8 V107 -1761886.9272790991
L8_107 V8 V107 1.2691966782303314e-11
C8_107 V8 V107 1.106146226641309e-20

R8_108 V8 V108 -405051.45173303667
L8_108 V8 V108 -6.3195805292057925e-12
C8_108 V8 V108 -3.2944386279216375e-20

R8_109 V8 V109 710548.8091259506
L8_109 V8 V109 8.950399179195294e-12
C8_109 V8 V109 4.732411197468093e-20

R8_110 V8 V110 5147812.981726497
L8_110 V8 V110 -6.827282228900113e-12
C8_110 V8 V110 -1.6147223653473145e-20

R8_111 V8 V111 -1069409.693839078
L8_111 V8 V111 -1.2210507963038134e-11
C8_111 V8 V111 -1.5397221989621665e-20

R8_112 V8 V112 -278592.6327197484
L8_112 V8 V112 7.444242480125658e-12
C8_112 V8 V112 1.5338405142377326e-20

R8_113 V8 V113 -180976.5737734351
L8_113 V8 V113 -1.0278050271433159e-10
C8_113 V8 V113 -1.5313729222769512e-20

R8_114 V8 V114 32393.125762564807
L8_114 V8 V114 1.1211307977345037e-11
C8_114 V8 V114 9.987053424095672e-21

R8_115 V8 V115 98570.10743284426
L8_115 V8 V115 2.3149279554296122e-11
C8_115 V8 V115 9.654177058672303e-21

R8_116 V8 V116 -182068.92027551835
L8_116 V8 V116 -9.041100760505859e-12
C8_116 V8 V116 -2.174512384757532e-20

R8_117 V8 V117 134324.87355783457
L8_117 V8 V117 -8.12005920213395e-11
C8_117 V8 V117 7.352701490568763e-21

R8_118 V8 V118 408279.2494520508
L8_118 V8 V118 -5.5013696761573564e-11
C8_118 V8 V118 8.686996028983903e-21

R8_119 V8 V119 -32847.482123334834
L8_119 V8 V119 -7.454932768492458e-12
C8_119 V8 V119 -2.455939144895537e-20

R8_120 V8 V120 197929.64558397862
L8_120 V8 V120 -1.5268058874374465e-11
C8_120 V8 V120 -1.981098493111321e-20

R8_121 V8 V121 -106298.07037120979
L8_121 V8 V121 5.5436347184521133e-11
C8_121 V8 V121 -2.755582714762998e-22

R8_122 V8 V122 358809.0908291126
L8_122 V8 V122 1.9772721570004523e-09
C8_122 V8 V122 2.2477834201449768e-21

R8_123 V8 V123 27607.531806162722
L8_123 V8 V123 -5.7609150080516115e-11
C8_123 V8 V123 -2.5825567780086263e-22

R8_124 V8 V124 47226.521485269346
L8_124 V8 V124 -2.822413257522855e-11
C8_124 V8 V124 -2.346525473111714e-20

R8_125 V8 V125 50397.67720444473
L8_125 V8 V125 -2.436852191551153e-11
C8_125 V8 V125 4.992593515144472e-22

R8_126 V8 V126 -179568.5186409118
L8_126 V8 V126 6.090399632321689e-11
C8_126 V8 V126 4.610795814145629e-22

R8_127 V8 V127 -513865.88974753045
L8_127 V8 V127 -1.647617698879646e-09
C8_127 V8 V127 -5.513684895540461e-21

R8_128 V8 V128 -76169.59502196473
L8_128 V8 V128 -1.0004116476902413e-10
C8_128 V8 V128 -9.75179195317477e-22

R8_129 V8 V129 22975.413483427492
L8_129 V8 V129 -5.0858448464966134e-11
C8_129 V8 V129 -6.2749423744912596e-21

R8_130 V8 V130 -19626.756190282442
L8_130 V8 V130 -1.3454767154084475e-10
C8_130 V8 V130 -5.071766432038832e-21

R8_131 V8 V131 -23777.31662499669
L8_131 V8 V131 2.6627534076029447e-11
C8_131 V8 V131 4.8410834735523846e-21

R8_132 V8 V132 -66106.81171685604
L8_132 V8 V132 -2.4566909655460433e-11
C8_132 V8 V132 -1.1779502079414156e-20

R8_133 V8 V133 -508254.7791682202
L8_133 V8 V133 2.3296313369861132e-11
C8_133 V8 V133 7.609085207799893e-21

R8_134 V8 V134 -303380.3098877164
L8_134 V8 V134 -2.867620593187542e-10
C8_134 V8 V134 4.661495083586535e-22

R8_135 V8 V135 318533.6592866913
L8_135 V8 V135 -1.4485036349693628e-10
C8_135 V8 V135 -4.080891184173862e-21

R8_136 V8 V136 471402.48892976163
L8_136 V8 V136 -1.3235422435293672e-10
C8_136 V8 V136 2.837995303828149e-21

R8_137 V8 V137 70203.15235494672
L8_137 V8 V137 -3.972054578896074e-11
C8_137 V8 V137 -8.89974903734013e-21

R8_138 V8 V138 -32039.60405049693
L8_138 V8 V138 1.209804289621861e-10
C8_138 V8 V138 -7.157476352451243e-21

R8_139 V8 V139 215979.83422243505
L8_139 V8 V139 1.830060489951692e-10
C8_139 V8 V139 2.0712983946479167e-21

R8_140 V8 V140 -66628.96692205647
L8_140 V8 V140 -2.5359747031314298e-11
C8_140 V8 V140 -1.1419382845915696e-21

R8_141 V8 V141 36895.69093901992
L8_141 V8 V141 -8.372365225453529e-10
C8_141 V8 V141 3.0780407400355433e-21

R8_142 V8 V142 -22249.879841688016
L8_142 V8 V142 -2.5378785670526816e-10
C8_142 V8 V142 -7.70586410283678e-21

R8_143 V8 V143 -63074.01534955186
L8_143 V8 V143 1.1314482285075122e-10
C8_143 V8 V143 -3.240344333546299e-21

R8_144 V8 V144 -1556113.630169789
L8_144 V8 V144 2.3058080759870573e-11
C8_144 V8 V144 -2.998826025612436e-21

R9_9 V9 0 -4806.867903142079
L9_9 V9 0 -5.353919861214214e-13
C9_9 V9 0 9.69487694232049e-19

R9_10 V9 V10 -217093.25765607922
L9_10 V9 V10 -5.1989800124840263e-11
C9_10 V9 V10 -2.0067526249676494e-21

R9_11 V9 V11 -112036.09398842748
L9_11 V9 V11 -7.586890616956034e-11
C9_11 V9 V11 -9.750941163293252e-21

R9_12 V9 V12 784265.4140148715
L9_12 V9 V12 4.958901070823464e-11
C9_12 V9 V12 2.3300117178822357e-21

R9_13 V9 V13 129227.34141118568
L9_13 V9 V13 -2.1293196346543148e-10
C9_13 V9 V13 5.511012607111629e-21

R9_14 V9 V14 726617.4048774291
L9_14 V9 V14 -4.5504940329544064e-11
C9_14 V9 V14 -2.8807165630561256e-21

R9_15 V9 V15 223039.58196688717
L9_15 V9 V15 -2.088688323779266e-10
C9_15 V9 V15 3.3479786213080875e-21

R9_16 V9 V16 473361.3360381707
L9_16 V9 V16 -4.069093573461812e-10
C9_16 V9 V16 1.1926562134256176e-21

R9_17 V9 V17 48127.55290979155
L9_17 V9 V17 -2.706861682122414e-11
C9_17 V9 V17 1.054292500317027e-20

R9_18 V9 V18 -1136793.1576059272
L9_18 V9 V18 -1.9421744503956906e-10
C9_18 V9 V18 -2.6126937487332936e-21

R9_19 V9 V19 87277.0843223081
L9_19 V9 V19 -5.3265617021267115e-11
C9_19 V9 V19 3.548753119849358e-21

R9_20 V9 V20 -3062926.4089521854
L9_20 V9 V20 -4.0591235225157097e-10
C9_20 V9 V20 1.004660871182293e-21

R9_21 V9 V21 -37080.49024163336
L9_21 V9 V21 -4.385518363117206e-12
C9_21 V9 V21 -1.860847311493799e-20

R9_22 V9 V22 217564.2346243229
L9_22 V9 V22 -8.677741619796539e-11
C9_22 V9 V22 4.814891838190558e-21

R9_23 V9 V23 272357.71753507253
L9_23 V9 V23 4.673871564030096e-11
C9_23 V9 V23 4.1098176057338056e-21

R9_24 V9 V24 7988180.310550582
L9_24 V9 V24 3.0114426046572384e-11
C9_24 V9 V24 -5.057398626556419e-22

R9_25 V9 V25 47865.94593450308
L9_25 V9 V25 -2.1333384066658664e-11
C9_25 V9 V25 -8.510096440388585e-21

R9_26 V9 V26 -593501.7098995969
L9_26 V9 V26 -6.997567018821944e-11
C9_26 V9 V26 -7.801080556589156e-22

R9_27 V9 V27 -695202.5673233353
L9_27 V9 V27 -8.703290126404357e-11
C9_27 V9 V27 -2.247454420170348e-21

R9_28 V9 V28 304612.4348410923
L9_28 V9 V28 -9.499871565757733e-10
C9_28 V9 V28 2.714583017566133e-22

R9_29 V9 V29 94395.3407334287
L9_29 V9 V29 -5.328757410350793e-12
C9_29 V9 V29 5.4185628335760335e-20

R9_30 V9 V30 1219906.0130436744
L9_30 V9 V30 -3.429332433189499e-11
C9_30 V9 V30 6.785165752159046e-21

R9_31 V9 V31 2750793.738723926
L9_31 V9 V31 -3.8397634923160187e-10
C9_31 V9 V31 1.5925834594543062e-20

R9_32 V9 V32 -217429.69946417617
L9_32 V9 V32 1.6696121479233506e-10
C9_32 V9 V32 9.28118737861513e-21

R9_33 V9 V33 113632.51762787065
L9_33 V9 V33 7.076668004915854e-12
C9_33 V9 V33 -4.2780947791665085e-20

R9_34 V9 V34 -112154.99321494317
L9_34 V9 V34 -1.7409091383092147e-11
C9_34 V9 V34 1.5007024984642698e-20

R9_35 V9 V35 111169.93934359781
L9_35 V9 V35 1.1093055363792345e-11
C9_35 V9 V35 -2.5954014166934643e-20

R9_36 V9 V36 181885.4705686117
L9_36 V9 V36 -3.340958706250411e-11
C9_36 V9 V36 6.5568506840010045e-22

R9_37 V9 V37 12514.23227163757
L9_37 V9 V37 -7.35761206576286e-12
C9_37 V9 V37 1.2869901836186816e-19

R9_38 V9 V38 438700.1876011256
L9_38 V9 V38 4.1585887263291876e-10
C9_38 V9 V38 -4.7074402897525766e-21

R9_39 V9 V39 17468.9168947968
L9_39 V9 V39 -7.718689642067157e-12
C9_39 V9 V39 1.0779283339717276e-19

R9_40 V9 V40 84713.58505191393
L9_40 V9 V40 6.17756189420297e-11
C9_40 V9 V40 2.1977905640615342e-20

R9_41 V9 V41 -7337.127382823305
L9_41 V9 V41 1.9320635512736047e-12
C9_41 V9 V41 -3.9568084833191185e-19

R9_42 V9 V42 -8586.565769700028
L9_42 V9 V42 2.2635892089787713e-12
C9_42 V9 V42 -2.688157676287855e-19

R9_43 V9 V43 -16313.110570210029
L9_43 V9 V43 5.0877080329629976e-12
C9_43 V9 V43 -1.5613716535944301e-19

R9_44 V9 V44 -93426.49764444091
L9_44 V9 V44 -1.1734566038437518e-10
C9_44 V9 V44 -3.363253081494927e-20

R9_45 V9 V45 5526.909495544675
L9_45 V9 V45 -4.988103234766978e-12
C9_45 V9 V45 3.028470584507199e-19

R9_46 V9 V46 11019.065047978262
L9_46 V9 V46 -2.2075655055852833e-11
C9_46 V9 V46 9.579097067376738e-20

R9_47 V9 V47 14831.839358323767
L9_47 V9 V47 -1.1094956735951453e-10
C9_47 V9 V47 4.344135007015311e-20

R9_48 V9 V48 46481.376920033756
L9_48 V9 V48 -2.37310997002408e-11
C9_48 V9 V48 2.116334044318701e-20

R9_49 V9 V49 -21371.145687020904
L9_49 V9 V49 1.0913658777069886e-11
C9_49 V9 V49 -7.874993531820794e-20

R9_50 V9 V50 164533.48522606087
L9_50 V9 V50 6.5499956662126585e-12
C9_50 V9 V50 -5.509768876424246e-20

R9_51 V9 V51 98682.75955539386
L9_51 V9 V51 -9.522710780471648e-12
C9_51 V9 V51 4.55829218970559e-20

R9_52 V9 V52 -15195.334537538623
L9_52 V9 V52 3.304007665216594e-12
C9_52 V9 V52 -1.8584109370311576e-19

R9_53 V9 V53 94722.01874095897
L9_53 V9 V53 4.242049864501559e-12
C9_53 V9 V53 -8.930137600445536e-20

R9_54 V9 V54 28237.8034810549
L9_54 V9 V54 1.2801071479905012e-11
C9_54 V9 V54 -7.76562718099171e-21

R9_55 V9 V55 295539.0631217737
L9_55 V9 V55 6.9088667124855356e-12
C9_55 V9 V55 -6.06724121688982e-20

R9_56 V9 V56 -54044.22802951166
L9_56 V9 V56 1.91340991422057e-11
C9_56 V9 V56 -5.709666676194558e-20

R9_57 V9 V57 3304.910641317613
L9_57 V9 V57 2.3024319659310554e-12
C9_57 V9 V57 3.72016291193611e-20

R9_58 V9 V58 23269.483097513712
L9_58 V9 V58 7.873216707915626e-12
C9_58 V9 V58 2.300782250112295e-20

R9_59 V9 V59 26199.379262670787
L9_59 V9 V59 -5.061260989676794e-10
C9_59 V9 V59 2.866618343551561e-20

R9_60 V9 V60 11804.511565112569
L9_60 V9 V60 2.3159639586558198e-11
C9_60 V9 V60 7.099627460294414e-21

R9_61 V9 V61 -6834.3813429709135
L9_61 V9 V61 3.581867887989736e-11
C9_61 V9 V61 -1.2465615271039422e-19

R9_62 V9 V62 -7724.56175429871
L9_62 V9 V62 -3.800166803017312e-10
C9_62 V9 V62 -1.0857350309647764e-19

R9_63 V9 V63 -16633.218670885442
L9_63 V9 V63 -3.931341936210806e-11
C9_63 V9 V63 -3.374384102820847e-20

R9_64 V9 V64 129886.55376500191
L9_64 V9 V64 3.7882472660814896e-11
C9_64 V9 V64 -1.6427953444752787e-20

R9_65 V9 V65 6600.748567922992
L9_65 V9 V65 2.4536467652070046e-12
C9_65 V9 V65 -4.420627773616518e-20

R9_66 V9 V66 6369.114908035692
L9_66 V9 V66 2.589561227205454e-12
C9_66 V9 V66 -2.3578707148768388e-20

R9_67 V9 V67 20007.47346222199
L9_67 V9 V67 1.3822920408085247e-11
C9_67 V9 V67 -2.4172072070143498e-20

R9_68 V9 V68 98402.39005325342
L9_68 V9 V68 4.746161997520881e-11
C9_68 V9 V68 -1.3527085965854474e-20

R9_69 V9 V69 -48545.094652972955
L9_69 V9 V69 -1.0807347430386912e-11
C9_69 V9 V69 8.484322320808093e-21

R9_70 V9 V70 -14635.000135286835
L9_70 V9 V70 -6.467568532831935e-12
C9_70 V9 V70 6.322242994190249e-21

R9_71 V9 V71 -14881.783921905077
L9_71 V9 V71 -8.676325572616003e-12
C9_71 V9 V71 -3.811797447203253e-21

R9_72 V9 V72 -14834.709802488842
L9_72 V9 V72 -5.020625089720752e-12
C9_72 V9 V72 8.269372403895612e-21

R9_73 V9 V73 -46885.80304850888
L9_73 V9 V73 -1.54150538095984e-11
C9_73 V9 V73 -6.071916730910549e-21

R9_74 V9 V74 -42542.6625818599
L9_74 V9 V74 -8.494530348162235e-12
C9_74 V9 V74 1.3076649348980871e-20

R9_75 V9 V75 33479.14864230783
L9_75 V9 V75 9.156813546841176e-12
C9_75 V9 V75 -2.3190035189024256e-20

R9_76 V9 V76 28999.699529515983
L9_76 V9 V76 1.3265505101348824e-11
C9_76 V9 V76 -1.194366117882867e-20

R9_77 V9 V77 112432.89310061838
L9_77 V9 V77 1.9315993923956713e-11
C9_77 V9 V77 -1.521575601560935e-20

R9_78 V9 V78 71213.57043630198
L9_78 V9 V78 5.907775639253907e-11
C9_78 V9 V78 8.666135860718132e-21

R9_79 V9 V79 -36207.25569367842
L9_79 V9 V79 -1.5117719368962025e-11
C9_79 V9 V79 -1.1784593298396068e-20

R9_80 V9 V80 -36267.23510267277
L9_80 V9 V80 3.1495259806578e-11
C9_80 V9 V80 -1.9778741300849915e-20

R9_81 V9 V81 -5100227.861570401
L9_81 V9 V81 -2.5098136894104257e-11
C9_81 V9 V81 3.667002541681437e-20

R9_82 V9 V82 -7343767.9793881355
L9_82 V9 V82 6.468732609552297e-12
C9_82 V9 V82 -4.93492052239262e-20

R9_83 V9 V83 -33390.53919603078
L9_83 V9 V83 -4.325020197173929e-11
C9_83 V9 V83 -3.1262463593070566e-20

R9_84 V9 V84 -262151.5315633999
L9_84 V9 V84 -6.429521390288138e-12
C9_84 V9 V84 1.0062616007174746e-20

R9_85 V9 V85 -78466.50182122487
L9_85 V9 V85 -6.71605568201693e-12
C9_85 V9 V85 2.3432786087863657e-20

R9_86 V9 V86 131528.61434612278
L9_86 V9 V86 -1.5155175891500257e-11
C9_86 V9 V86 2.1537546273160205e-20

R9_87 V9 V87 68088.36240032299
L9_87 V9 V87 -9.737753550996215e-12
C9_87 V9 V87 3.054278046721135e-20

R9_88 V9 V88 222027.44592221457
L9_88 V9 V88 7.942701717285573e-11
C9_88 V9 V88 1.0172790062412382e-20

R9_89 V9 V89 -113982.63820819101
L9_89 V9 V89 5.727195231122362e-12
C9_89 V9 V89 -4.4778883628390177e-20

R9_90 V9 V90 -137239.28194693523
L9_90 V9 V90 1.4355252836944737e-11
C9_90 V9 V90 5.154252810346365e-21

R9_91 V9 V91 -53854.19004115482
L9_91 V9 V91 1.2853747403805315e-11
C9_91 V9 V91 -3.5649688404234196e-20

R9_92 V9 V92 -55810.61392047037
L9_92 V9 V92 3.7234812910282475e-11
C9_92 V9 V92 -4.2585244352804006e-20

R9_93 V9 V93 -22415.61349979753
L9_93 V9 V93 -3.4373505978158194e-11
C9_93 V9 V93 -4.711887312432049e-21

R9_94 V9 V94 94168.72487514577
L9_94 V9 V94 -2.19667870486887e-11
C9_94 V9 V94 3.1400119711854817e-20

R9_95 V9 V95 -58523.665974589494
L9_95 V9 V95 3.4656838452146187e-11
C9_95 V9 V95 -2.0511304518787602e-20

R9_96 V9 V96 -109069.02341608636
L9_96 V9 V96 -6.505131231140233e-11
C9_96 V9 V96 -3.0440037142344204e-20

R9_97 V9 V97 -356024.22993310075
L9_97 V9 V97 1.3284206755001574e-11
C9_97 V9 V97 1.7326935542757356e-20

R9_98 V9 V98 -63900.58864351982
L9_98 V9 V98 6.85820176037982e-12
C9_98 V9 V98 -3.054890933146321e-20

R9_99 V9 V99 83852.52173691647
L9_99 V9 V99 -7.128150868897797e-11
C9_99 V9 V99 5.000309672016683e-21

R9_100 V9 V100 110856.0992836712
L9_100 V9 V100 -1.8812758126016207e-10
C9_100 V9 V100 1.7962128466933627e-20

R9_101 V9 V101 -35698.0676348208
L9_101 V9 V101 5.718945841228615e-12
C9_101 V9 V101 -5.327797336168463e-20

R9_102 V9 V102 -44433.94241231065
L9_102 V9 V102 5.155674100496367e-12
C9_102 V9 V102 -1.462611577543334e-20

R9_103 V9 V103 -73935.83747638708
L9_103 V9 V103 -3.4453547978008415e-11
C9_103 V9 V103 -1.4963209735127322e-20

R9_104 V9 V104 -208943.04812371838
L9_104 V9 V104 -2.810226035288829e-11
C9_104 V9 V104 -1.410599563752646e-20

R9_105 V9 V105 46276.285965896204
L9_105 V9 V105 -1.2758948901921599e-11
C9_105 V9 V105 3.486380639184152e-20

R9_106 V9 V106 -68681.17083425405
L9_106 V9 V106 1.3090779026586713e-11
C9_106 V9 V106 -5.0521770023567676e-20

R9_107 V9 V107 100097.75554645565
L9_107 V9 V107 1.0932784205081832e-11
C9_107 V9 V107 5.945998179721743e-21

R9_108 V9 V108 51669.377401245845
L9_108 V9 V108 -6.2811060086754915e-12
C9_108 V9 V108 4.3575373957932456e-20

R9_109 V9 V109 131459.0909355125
L9_109 V9 V109 -1.7572831782062204e-11
C9_109 V9 V109 -8.597380476828556e-21

R9_110 V9 V110 -231685.51618063878
L9_110 V9 V110 -7.903477978458883e-12
C9_110 V9 V110 5.461090531130701e-20

R9_111 V9 V111 31335.41540812046
L9_111 V9 V111 -4.8784889989783154e-11
C9_111 V9 V111 8.40120556868415e-21

R9_112 V9 V112 -145003.30987425803
L9_112 V9 V112 4.397150342450268e-12
C9_112 V9 V112 -3.1269721581726213e-20

R9_113 V9 V113 1359787.6031173624
L9_113 V9 V113 9.412914190404752e-12
C9_113 V9 V113 -4.650269229637603e-21

R9_114 V9 V114 -36827.83632682322
L9_114 V9 V114 1.4515777860278024e-11
C9_114 V9 V114 -3.054765124658347e-20

R9_115 V9 V115 -64667.72064768887
L9_115 V9 V115 6.199149139570944e-11
C9_115 V9 V115 6.635921340262386e-21

R9_116 V9 V116 58163.545936673705
L9_116 V9 V116 -7.568289029525778e-12
C9_116 V9 V116 2.817550371281938e-20

R9_117 V9 V117 -64816.790376654026
L9_117 V9 V117 -1.0088720627398885e-11
C9_117 V9 V117 1.2195038324777474e-20

R9_118 V9 V118 74747.09659127165
L9_118 V9 V118 -9.52171244337994e-12
C9_118 V9 V118 1.9389173872463793e-20

R9_119 V9 V119 19510.152937504106
L9_119 V9 V119 -2.113916484163893e-11
C9_119 V9 V119 3.6925664104692496e-20

R9_120 V9 V120 -11345.469421237629
L9_120 V9 V120 -2.035534349226992e-11
C9_120 V9 V120 9.14042770007854e-21

R9_121 V9 V121 27214.156404212594
L9_121 V9 V121 7.765585349916088e-12
C9_121 V9 V121 -1.4489194287133895e-21

R9_122 V9 V122 -29892.550195767555
L9_122 V9 V122 5.919615706700608e-12
C9_122 V9 V122 1.2548966805799327e-21

R9_123 V9 V123 -40696.38056270413
L9_123 V9 V123 4.3372067310636375e-11
C9_123 V9 V123 5.935200475457555e-22

R9_124 V9 V124 534277.6760478953
L9_124 V9 V124 3.978214343453881e-10
C9_124 V9 V124 6.914069207578022e-21

R9_125 V9 V125 -14686.71130532583
L9_125 V9 V125 -5.52764448393126e-12
C9_125 V9 V125 1.1535141655321366e-20

R9_126 V9 V126 12075.64905154164
L9_126 V9 V126 -8.79805945739768e-12
C9_126 V9 V126 -1.872558577639778e-21

R9_127 V9 V127 -12861.665827233186
L9_127 V9 V127 1.6886610977971393e-11
C9_127 V9 V127 5.529682875866017e-22

R9_128 V9 V128 -135359.46390633276
L9_128 V9 V128 5.350725164118129e-11
C9_128 V9 V128 -1.961991810623693e-21

R9_129 V9 V129 -24200.364913091078
L9_129 V9 V129 9.737033376678863e-11
C9_129 V9 V129 1.9578441342682875e-21

R9_130 V9 V130 29328.79530060148
L9_130 V9 V130 -1.8996424997911246e-11
C9_130 V9 V130 5.368108776800116e-21

R9_131 V9 V131 36584.69799909666
L9_131 V9 V131 -3.835009877797132e-11
C9_131 V9 V131 7.768771416276745e-22

R9_132 V9 V132 51330.226732167976
L9_132 V9 V132 -5.0033982352819155e-11
C9_132 V9 V132 2.6269972167672644e-21

R9_133 V9 V133 -173954.73293958497
L9_133 V9 V133 -4.4209652335109925e-11
C9_133 V9 V133 -1.5372776138017854e-20

R9_134 V9 V134 68050.39571471956
L9_134 V9 V134 -1.8947043820060638e-11
C9_134 V9 V134 -1.7201397727921763e-22

R9_135 V9 V135 -19774.78095042547
L9_135 V9 V135 2.7417521983875537e-11
C9_135 V9 V135 -1.5212396107151164e-21

R9_136 V9 V136 -165468.28313367863
L9_136 V9 V136 -7.924950464027989e-11
C9_136 V9 V136 1.4834021271501227e-21

R9_137 V9 V137 -23979.901950338164
L9_137 V9 V137 -1.1258352921919969e-11
C9_137 V9 V137 9.481475640245276e-21

R9_138 V9 V138 14652.796444611567
L9_138 V9 V138 -8.28268656775317e-12
C9_138 V9 V138 -4.4794880339484475e-21

R9_139 V9 V139 -9473.093264901478
L9_139 V9 V139 1.2150746842959074e-11
C9_139 V9 V139 3.747278158946924e-21

R9_140 V9 V140 25693.61406589521
L9_140 V9 V140 -1.7005128078498952e-11
C9_140 V9 V140 8.738932196421856e-21

R9_141 V9 V141 204066.37448957778
L9_141 V9 V141 -3.349638137385971e-11
C9_141 V9 V141 -3.506146271804068e-22

R9_142 V9 V142 19605.45460342889
L9_142 V9 V142 -2.3048937406718498e-11
C9_142 V9 V142 6.356086821671733e-21

R9_143 V9 V143 25589.721847331584
L9_143 V9 V143 -5.0660316764807166e-11
C9_143 V9 V143 8.386875667349955e-22

R9_144 V9 V144 -309610.71427554067
L9_144 V9 V144 5.499813973294685e-11
C9_144 V9 V144 -4.626710372370925e-21

R10_10 V10 0 -2864.0119840095977
L10_10 V10 0 8.570579482689701e-13
C10_10 V10 0 1.4226797424496013e-19

R10_11 V10 V11 -384887.7651601429
L10_11 V10 V11 1.5245497867914786e-11
C10_11 V10 V11 -1.1413602985186877e-21

R10_12 V10 V12 39768662.46362014
L10_12 V10 V12 2.254854767571768e-10
C10_12 V10 V12 1.412026495510377e-21

R10_13 V10 V13 281760.1773006562
L10_13 V10 V13 1.3059010453851194e-10
C10_13 V10 V13 -3.8170720543564896e-22

R10_14 V10 V14 -3224596.4016652727
L10_14 V10 V14 -1.476005112842666e-11
C10_14 V10 V14 1.7197452424610912e-21

R10_15 V10 V15 639432.6597924015
L10_15 V10 V15 -3.913985421041202e-11
C10_15 V10 V15 7.995595987176766e-22

R10_16 V10 V16 -2705403.9265726595
L10_16 V10 V16 -3.965017541301197e-11
C10_16 V10 V16 5.297384242873338e-22

R10_17 V10 V17 109554.19234948784
L10_17 V10 V17 -2.5772448272749885e-11
C10_17 V10 V17 2.120516676242135e-21

R10_18 V10 V18 -3129956.760082247
L10_18 V10 V18 -4.8420159491950225e-11
C10_18 V10 V18 7.153258847410566e-22

R10_19 V10 V19 168612.90329646782
L10_19 V10 V19 6.657367595823048e-11
C10_19 V10 V19 7.1045604896882035e-22

R10_20 V10 V20 -252550.8769384456
L10_20 V10 V20 3.854047606854667e-11
C10_20 V10 V20 -3.6404582816183416e-21

R10_21 V10 V21 -112807.9576350794
L10_21 V10 V21 -4.309183072821974e-11
C10_21 V10 V21 -5.267891960363455e-21

R10_22 V10 V22 -5092202.565788108
L10_22 V10 V22 -3.8050074867454044e-12
C10_22 V10 V22 -2.2120400738426045e-22

R10_23 V10 V23 400960.65421115403
L10_23 V10 V23 3.0278076441198595e-11
C10_23 V10 V23 1.834335890635341e-21

R10_24 V10 V24 653003.7289221239
L10_24 V10 V24 -6.03602876182998e-10
C10_24 V10 V24 1.976920060344062e-21

R10_25 V10 V25 105827.28973846501
L10_25 V10 V25 6.571329668860323e-11
C10_25 V10 V25 -1.173421662820187e-21

R10_26 V10 V26 2901375.625296263
L10_26 V10 V26 -7.022139326875593e-12
C10_26 V10 V26 -3.636389895764507e-21

R10_27 V10 V27 -362815.4602968141
L10_27 V10 V27 -2.478680322541943e-11
C10_27 V10 V27 -3.0061655291036884e-22

R10_28 V10 V28 -238320.78812792985
L10_28 V10 V28 -1.8636460491789653e-11
C10_28 V10 V28 1.4135403550641267e-22

R10_29 V10 V29 1957622.3126764758
L10_29 V10 V29 5.541528441417577e-11
C10_29 V10 V29 9.650608632717255e-21

R10_30 V10 V30 -1451486.6443750751
L10_30 V10 V30 -7.633946763060464e-12
C10_30 V10 V30 3.651929071169692e-21

R10_31 V10 V31 -1134287.61187697
L10_31 V10 V31 2.4049639508706172e-11
C10_31 V10 V31 -1.0478188272864614e-21

R10_32 V10 V32 148791.44998507705
L10_32 V10 V32 6.452602348010994e-10
C10_32 V10 V32 -3.70381612887786e-21

R10_33 V10 V33 79973.59866072868
L10_33 V10 V33 -3.3651871845582786e-11
C10_33 V10 V33 -8.740620548271178e-21

R10_34 V10 V34 -131189.90039541273
L10_34 V10 V34 -1.0057926443039232e-09
C10_34 V10 V34 -3.923431317854808e-22

R10_35 V10 V35 154911.50581757925
L10_35 V10 V35 -7.548566105945121e-11
C10_35 V10 V35 -8.493618079371853e-22

R10_36 V10 V36 -54340.88814328456
L10_36 V10 V36 -3.2021779108196665e-10
C10_36 V10 V36 2.0798949886937153e-21

R10_37 V10 V37 63914.51827095693
L10_37 V10 V37 2.2659804240097954e-11
C10_37 V10 V37 2.0731968440729668e-20

R10_38 V10 V38 103850.08293406009
L10_38 V10 V38 -1.6934953956436252e-11
C10_38 V10 V38 1.4833216156099232e-20

R10_39 V10 V39 119286.33453713273
L10_39 V10 V39 5.237545729421583e-11
C10_39 V10 V39 1.1628253457352036e-20

R10_40 V10 V40 4080015.7727708668
L10_40 V10 V40 1.0835682526875487e-10
C10_40 V10 V40 -1.971819850809978e-20

R10_41 V10 V41 51049.4157775511
L10_41 V10 V41 -5.995263199280628e-12
C10_41 V10 V41 -6.143865976129922e-20

R10_42 V10 V42 -41577.42069605865
L10_42 V10 V42 1.0696287970131289e-11
C10_42 V10 V42 -8.941607033466833e-20

R10_43 V10 V43 399342.5355786606
L10_43 V10 V43 -6.452345504902524e-11
C10_43 V10 V43 -4.332427401059939e-22

R10_44 V10 V44 -102578.14452618835
L10_44 V10 V44 1.71399599751709e-11
C10_44 V10 V44 3.1494026251363187e-20

R10_45 V10 V45 18431.41894299097
L10_45 V10 V45 3.5931431859127767e-09
C10_45 V10 V45 2.9945341862906384e-20

R10_46 V10 V46 16655.389230357705
L10_46 V10 V46 -1.9946346755425218e-10
C10_46 V10 V46 5.973892506939552e-20

R10_47 V10 V47 138400.97095244948
L10_47 V10 V47 -1.9960693138355833e-11
C10_47 V10 V47 -7.216412196271563e-21

R10_48 V10 V48 -29221.814298233567
L10_48 V10 V48 -3.0474838333187485e-11
C10_48 V10 V48 -9.615967089128354e-21

R10_49 V10 V49 -109046.71961936328
L10_49 V10 V49 4.808074669199282e-11
C10_49 V10 V49 -8.899859802266994e-21

R10_50 V10 V50 159093.21387800534
L10_50 V10 V50 1.8331292130342726e-11
C10_50 V10 V50 -1.7418126022987817e-20

R10_51 V10 V51 -298369.48986901244
L10_51 V10 V51 -1.3640984073045249e-11
C10_51 V10 V51 2.9366213533945126e-20

R10_52 V10 V52 3732208.3365697935
L10_52 V10 V52 1.6207615192320175e-11
C10_52 V10 V52 -3.038270665404621e-20

R10_53 V10 V53 -269673.54219872993
L10_53 V10 V53 -1.6318786585388878e-11
C10_53 V10 V53 -2.575450832915808e-20

R10_54 V10 V54 65130.69046699046
L10_54 V10 V54 -6.873877459041265e-11
C10_54 V10 V54 -1.7250329498095534e-20

R10_55 V10 V55 35704.28245343029
L10_55 V10 V55 3.4579607514092496e-11
C10_55 V10 V55 -6.507538522815771e-21

R10_56 V10 V56 21625.121375605642
L10_56 V10 V56 -1.825881700474626e-11
C10_56 V10 V56 7.989348624467857e-21

R10_57 V10 V57 4800.358432784308
L10_57 V10 V57 -1.0011377213001245e-11
C10_57 V10 V57 9.66755422934308e-21

R10_58 V10 V58 12273.516880523444
L10_58 V10 V58 3.5308355608215654e-11
C10_58 V10 V58 3.2627762284621572e-21

R10_59 V10 V59 64976.90113335742
L10_59 V10 V59 -3.34418919990321e-11
C10_59 V10 V59 5.258599385086768e-21

R10_60 V10 V60 -34974.83995090931
L10_60 V10 V60 1.0971990446014227e-10
C10_60 V10 V60 1.6537534709434591e-21

R10_61 V10 V61 -14066.989754755932
L10_61 V10 V61 -2.096476188982934e-11
C10_61 V10 V61 -2.7329137757986217e-20

R10_62 V10 V62 -10859.735557172025
L10_62 V10 V62 1.3170140374615813e-11
C10_62 V10 V62 -2.088306120174334e-20

R10_63 V10 V63 436220.88606331067
L10_63 V10 V63 -2.5361625682642124e-11
C10_63 V10 V63 1.359083453988668e-21

R10_64 V10 V64 93178.38721953056
L10_64 V10 V64 -1.0189818422323068e-11
C10_64 V10 V64 4.634401392101319e-21

R10_65 V10 V65 10346.426965431792
L10_65 V10 V65 1.3520230026427331e-11
C10_65 V10 V65 -8.50646293653064e-21

R10_66 V10 V66 10687.085916117652
L10_66 V10 V66 -4.331085656135321e-11
C10_66 V10 V66 -8.630267328595385e-21

R10_67 V10 V67 104929.90236616576
L10_67 V10 V67 -1.9372775504599282e-11
C10_67 V10 V67 1.973814769361505e-21

R10_68 V10 V68 -91321.70718266614
L10_68 V10 V68 3.19728032434921e-11
C10_68 V10 V68 1.1929115296631857e-21

R10_69 V10 V69 -66468.77162836364
L10_69 V10 V69 -1.225135712486891e-11
C10_69 V10 V69 7.083226314917303e-21

R10_70 V10 V70 -32542.98525189724
L10_70 V10 V70 -6.806389376119906e-12
C10_70 V10 V70 -1.0679708958519271e-20

R10_71 V10 V71 -161826.88698888934
L10_71 V10 V71 -2.207980982122426e-11
C10_71 V10 V71 3.448062146103808e-21

R10_72 V10 V72 -26312.46102818284
L10_72 V10 V72 -9.554187551864429e-12
C10_72 V10 V72 -4.089743254785398e-21

R10_73 V10 V73 -56851.78226837668
L10_73 V10 V73 -1.0300982397816209e-11
C10_73 V10 V73 -8.847833709762532e-21

R10_74 V10 V74 -48763.0055521088
L10_74 V10 V74 -7.943560161567002e-12
C10_74 V10 V74 1.665673243508371e-21

R10_75 V10 V75 48372.40181530972
L10_75 V10 V75 8.576978086067527e-12
C10_75 V10 V75 -1.9408085695173675e-22

R10_76 V10 V76 75059.88966617288
L10_76 V10 V76 -5.707091807675218e-12
C10_76 V10 V76 -1.190123717528801e-20

R10_77 V10 V77 96283.0483628089
L10_77 V10 V77 -3.6451257353069625e-10
C10_77 V10 V77 1.1931334155778879e-21

R10_78 V10 V78 -228232.41990307966
L10_78 V10 V78 -1.29084798302853e-11
C10_78 V10 V78 -7.05024639196336e-21

R10_79 V10 V79 -71094.286015542
L10_79 V10 V79 -3.853405828734678e-12
C10_79 V10 V79 -4.401309926608801e-21

R10_80 V10 V80 -151293.10465864177
L10_80 V10 V80 5.169453421184554e-12
C10_80 V10 V80 1.1976301594620183e-20

R10_81 V10 V81 -76069.28226791826
L10_81 V10 V81 -1.1973301136660054e-11
C10_81 V10 V81 -1.8380919266404618e-20

R10_82 V10 V82 105225.14800229497
L10_82 V10 V82 5.297047128146844e-12
C10_82 V10 V82 2.898131883107573e-20

R10_83 V10 V83 110655.65818202266
L10_83 V10 V83 4.439005321883503e-12
C10_83 V10 V83 2.6847276690528874e-20

R10_84 V10 V84 -949963.8543444021
L10_84 V10 V84 -7.070001172481813e-12
C10_84 V10 V84 4.505663169304895e-21

R10_85 V10 V85 -87289.14805351186
L10_85 V10 V85 -4.273009781697854e-12
C10_85 V10 V85 -6.506221805371e-21

R10_86 V10 V86 -115462.47651325913
L10_86 V10 V86 -1.3787684140198838e-11
C10_86 V10 V86 -7.807486312832663e-21

R10_87 V10 V87 -248214.71933760354
L10_87 V10 V87 -4.794301277936616e-12
C10_87 V10 V87 -2.0454448572733308e-20

R10_88 V10 V88 -114358.84338416425
L10_88 V10 V88 -1.588814404402438e-10
C10_88 V10 V88 -8.618679529651298e-21

R10_89 V10 V89 144809.38460617364
L10_89 V10 V89 2.0988666354722553e-11
C10_89 V10 V89 8.13296789958131e-21

R10_90 V10 V90 343652.31766028854
L10_90 V10 V90 4.034330950960717e-12
C10_90 V10 V90 -3.0897030413866953e-21

R10_91 V10 V91 132197.12967051362
L10_91 V10 V91 7.554369764524335e-12
C10_91 V10 V91 2.070847631864109e-20

R10_92 V10 V92 130031.8853513278
L10_92 V10 V92 6.614248139656585e-12
C10_92 V10 V92 2.6049886616978318e-20

R10_93 V10 V93 -28290.575485415327
L10_93 V10 V93 -1.155297115079739e-11
C10_93 V10 V93 -4.7432916044849575e-21

R10_94 V10 V94 -49573.01477349295
L10_94 V10 V94 -3.05543612118367e-11
C10_94 V10 V94 -1.76227376892078e-20

R10_95 V10 V95 -879314.8472579509
L10_95 V10 V95 1.1387047721530813e-11
C10_95 V10 V95 1.3979988201949994e-20

R10_96 V10 V96 100892.71429431508
L10_96 V10 V96 6.803464670689813e-12
C10_96 V10 V96 2.4504371679828243e-20

R10_97 V10 V97 1122756.3691839152
L10_97 V10 V97 1.1119042763401608e-11
C10_97 V10 V97 -1.1851480978037358e-20

R10_98 V10 V98 48219.88654738687
L10_98 V10 V98 5.570800184758335e-12
C10_98 V10 V98 1.5719110130499776e-20

R10_99 V10 V99 -176277.5798792557
L10_99 V10 V99 -7.610080088275774e-12
C10_99 V10 V99 -6.230778437726281e-21

R10_100 V10 V100 -1268144.3971433851
L10_100 V10 V100 -3.2373531643890594e-11
C10_100 V10 V100 -1.1534075128886919e-20

R10_101 V10 V101 -420019.73852406867
L10_101 V10 V101 9.407358168381955e-12
C10_101 V10 V101 1.5300663207217605e-20

R10_102 V10 V102 426557.0060853311
L10_102 V10 V102 1.835846788966042e-12
C10_102 V10 V102 5.444344158980558e-22

R10_103 V10 V103 354078.92201963713
L10_103 V10 V103 -3.380895285456712e-12
C10_103 V10 V103 2.6752817593078002e-21

R10_104 V10 V104 -498741.4536056545
L10_104 V10 V104 6.974678977308323e-11
C10_104 V10 V104 9.390779278235581e-21

R10_105 V10 V105 -236267.14833719068
L10_105 V10 V105 -3.7057231178854776e-12
C10_105 V10 V105 -2.1631320114727022e-20

R10_106 V10 V106 844077.789345879
L10_106 V10 V106 2.4839844653976454e-12
C10_106 V10 V106 3.309912718542582e-20

R10_107 V10 V107 179253.10522847273
L10_107 V10 V107 2.128993725503958e-12
C10_107 V10 V107 1.0885841963642457e-20

R10_108 V10 V108 57500.18003118639
L10_108 V10 V108 -2.4463830573146463e-12
C10_108 V10 V108 -1.548879247577023e-20

R10_109 V10 V109 84323.81448419235
L10_109 V10 V109 -6.060018340384505e-12
C10_109 V10 V109 1.1379171277289621e-20

R10_110 V10 V110 -210691.17672998158
L10_110 V10 V110 -5.102438876765503e-12
C10_110 V10 V110 -2.922705165953095e-20

R10_111 V10 V111 57006.888996654896
L10_111 V10 V111 -3.148878758746233e-12
C10_111 V10 V111 -1.5058594802844373e-20

R10_112 V10 V112 30303.826688850495
L10_112 V10 V112 2.6318795703637327e-12
C10_112 V10 V112 1.2657332164328225e-20

R10_113 V10 V113 60504.83394009447
L10_113 V10 V113 6.243164386625523e-12
C10_113 V10 V113 -9.90874507993822e-22

R10_114 V10 V114 110454.8247877658
L10_114 V10 V114 4.9751239687579325e-12
C10_114 V10 V114 2.1520735126016693e-20

R10_115 V10 V115 -428217.9855314069
L10_115 V10 V115 4.291733252643637e-12
C10_115 V10 V115 3.3341279002279734e-21

R10_116 V10 V116 -982574.8236792424
L10_116 V10 V116 -4.261897579068423e-12
C10_116 V10 V116 -6.4823002102568195e-21

R10_117 V10 V117 -163975.95174248345
L10_117 V10 V117 -8.55032350744844e-12
C10_117 V10 V117 3.0166846440899763e-21

R10_118 V10 V118 -243643.7540187898
L10_118 V10 V118 -5.9973853432709995e-12
C10_118 V10 V118 -1.1779040567284688e-20

R10_119 V10 V119 86629.41549111146
L10_119 V10 V119 -4.068246135899694e-12
C10_119 V10 V119 -2.3118970750482643e-20

R10_120 V10 V120 -30481.193725895166
L10_120 V10 V120 6.262539603593745e-12
C10_120 V10 V120 -1.0319121660259972e-20

R10_121 V10 V121 19380.98712602712
L10_121 V10 V121 1.8597580156739525e-11
C10_121 V10 V121 1.6675729815059852e-21

R10_122 V10 V122 16296.445288136865
L10_122 V10 V122 3.895134065515365e-12
C10_122 V10 V122 1.7822247000443694e-23

R10_123 V10 V123 76576.84208269109
L10_123 V10 V123 2.471735870448585e-11
C10_123 V10 V123 -2.1275052662284403e-21

R10_124 V10 V124 103167.33119650299
L10_124 V10 V124 -1.616322010529098e-11
C10_124 V10 V124 -1.1560111184107206e-20

R10_125 V10 V125 -16455.376505462507
L10_125 V10 V125 5.569792944522932e-11
C10_125 V10 V125 -2.8778499260288367e-21

R10_126 V10 V126 -33207.00620433593
L10_126 V10 V126 -2.919939335371818e-12
C10_126 V10 V126 -2.4727844167401603e-21

R10_127 V10 V127 375456.29445282347
L10_127 V10 V127 3.223764884477963e-12
C10_127 V10 V127 -1.751912021231684e-21

R10_128 V10 V128 -148568.00300431476
L10_128 V10 V128 3.376560820213964e-11
C10_128 V10 V128 -5.047154170081695e-22

R10_129 V10 V129 86193.40486178648
L10_129 V10 V129 9.618667139298061e-12
C10_129 V10 V129 -1.3908534994797014e-22

R10_130 V10 V130 -67536.44903049877
L10_130 V10 V130 -4.82689849471338e-12
C10_130 V10 V130 -3.818628498433927e-21

R10_131 V10 V131 -43318.07505794757
L10_131 V10 V131 3.3529301713556133e-11
C10_131 V10 V131 8.931425075119496e-22

R10_132 V10 V132 -114867.53067566747
L10_132 V10 V132 -1.252423454790351e-11
C10_132 V10 V132 3.435356170187216e-22

R10_133 V10 V133 -92821.08726315509
L10_133 V10 V133 1.0507682073806806e-11
C10_133 V10 V133 1.0404546518475644e-20

R10_134 V10 V134 -99459.68321820816
L10_134 V10 V134 -3.824280923740316e-11
C10_134 V10 V134 -2.5635191775396234e-21

R10_135 V10 V135 136858.4449288383
L10_135 V10 V135 5.783553510353327e-12
C10_135 V10 V135 -4.43503101610682e-21

R10_136 V10 V136 -174518.42714869572
L10_136 V10 V136 2.550223509955227e-10
C10_136 V10 V136 -3.712025661163601e-21

R10_137 V10 V137 -26149.272961001112
L10_137 V10 V137 -2.70050589714882e-11
C10_137 V10 V137 -1.0611915889279993e-20

R10_138 V10 V138 -25136.17775365937
L10_138 V10 V138 -3.188947769120741e-12
C10_138 V10 V138 -5.820737311904773e-22

R10_139 V10 V139 534084.0070235914
L10_139 V10 V139 2.3485609868573986e-12
C10_139 V10 V139 4.958900678129445e-21

R10_140 V10 V140 -193829.22863992126
L10_140 V10 V140 -5.7615589327832806e-12
C10_140 V10 V140 1.7719074250043137e-22

R10_141 V10 V141 -229461.32500311124
L10_141 V10 V141 -1.1196195867268892e-11
C10_141 V10 V141 4.875646324659387e-22

R10_142 V10 V142 -120559.79137991642
L10_142 V10 V142 -5.806002747233695e-12
C10_142 V10 V142 -2.8202768656732797e-21

R10_143 V10 V143 2138542.6218293
L10_143 V10 V143 -8.734544198012701e-12
C10_143 V10 V143 2.0858395943316153e-22

R10_144 V10 V144 63972.63491859698
L10_144 V10 V144 1.1855235121238154e-11
C10_144 V10 V144 -1.903862078616758e-21

R11_11 V11 0 -2631.598343745641
L11_11 V11 0 -7.820357118156757e-13
C11_11 V11 0 4.0600673963072685e-19

R11_12 V11 V12 2342941.37581182
L11_12 V11 V12 -3.5777224177601576e-11
C11_12 V11 V12 2.1830458778215145e-21

R11_13 V11 V13 174995.0479199129
L11_13 V11 V13 5.004489510763604e-11
C11_13 V11 V13 2.058156278463753e-21

R11_14 V11 V14 7498187.855672675
L11_14 V11 V14 -2.6697731234241053e-10
C11_14 V11 V14 -1.5335232250238969e-22

R11_15 V11 V15 719984.6403698231
L11_15 V11 V15 -6.891749153623002e-11
C11_15 V11 V15 2.848020495319674e-21

R11_16 V11 V16 5204029.040569117
L11_16 V11 V16 5.578821843609041e-09
C11_16 V11 V16 3.7612351356193257e-22

R11_17 V11 V17 69563.59502139267
L11_17 V11 V17 1.3718420241499925e-10
C11_17 V11 V17 5.5785638588802636e-21

R11_18 V11 V18 1448155.8461824446
L11_18 V11 V18 4.6709120632497247e-11
C11_18 V11 V18 -1.2682947424653418e-21

R11_19 V11 V19 132664.59974373647
L11_19 V11 V19 -2.346105738521341e-10
C11_19 V11 V19 2.6024910821738365e-21

R11_20 V11 V20 -156805.27689014707
L11_20 V11 V20 4.8592346937815264e-11
C11_20 V11 V20 -3.913832346172696e-21

R11_21 V11 V21 -61986.865892063935
L11_21 V11 V21 -1.600269296642491e-11
C11_21 V11 V21 -1.0515379919495031e-20

R11_22 V11 V22 382501.8684780216
L11_22 V11 V22 4.385721530051828e-12
C11_22 V11 V22 1.994224987691038e-21

R11_23 V11 V23 436020.9616295861
L11_23 V11 V23 -1.0595285931707948e-11
C11_23 V11 V23 1.8996860338220203e-21

R11_24 V11 V24 606731.5398289929
L11_24 V11 V24 -1.6492086455932294e-11
C11_24 V11 V24 2.304964256832224e-21

R11_25 V11 V25 62350.982030265346
L11_25 V11 V25 -5.921110671752208e-11
C11_25 V11 V25 -3.826490462463887e-21

R11_26 V11 V26 -821182.5761632555
L11_26 V11 V26 7.332049459832317e-12
C11_26 V11 V26 -1.8974866131790147e-22

R11_27 V11 V27 -889711.6344289327
L11_27 V11 V27 6.384439699459733e-11
C11_27 V11 V27 -1.9518949461577043e-21

R11_28 V11 V28 -265507.7026174821
L11_28 V11 V28 -9.26842589390592e-11
C11_28 V11 V28 -1.0040977788939193e-24

R11_29 V11 V29 367867.32903998945
L11_29 V11 V29 -1.5441640236407386e-11
C11_29 V11 V29 2.6586877350976315e-20

R11_30 V11 V30 6291147.811701299
L11_30 V11 V30 8.001083116365211e-12
C11_30 V11 V30 2.8870491016041844e-21

R11_31 V11 V31 4257645.528525344
L11_31 V11 V31 -1.4520065340918383e-11
C11_31 V11 V31 7.515757872985596e-21

R11_32 V11 V32 136523.33659787374
L11_32 V11 V32 -2.221456721764255e-11
C11_32 V11 V32 -8.895733285129956e-22

R11_33 V11 V33 73830.95473212043
L11_33 V11 V33 1.851330006866921e-11
C11_33 V11 V33 -2.007015126787631e-20

R11_34 V11 V34 -101198.7672787906
L11_34 V11 V34 -3.4314351587693466e-11
C11_34 V11 V34 8.897144963435775e-21

R11_35 V11 V35 125065.09504169815
L11_35 V11 V35 1.868552091532407e-11
C11_35 V11 V35 -1.0353974443120841e-20

R11_36 V11 V36 -44713.81664763122
L11_36 V11 V36 2.2902295680065515e-10
C11_36 V11 V36 2.50064999566894e-21

R11_37 V11 V37 24086.21489749268
L11_37 V11 V37 -2.380047441882036e-11
C11_37 V11 V37 6.280394484789107e-20

R11_38 V11 V38 360806.6564711728
L11_38 V11 V38 1.323252962828015e-11
C11_38 V11 V38 -2.1985672372018753e-21

R11_39 V11 V39 34240.632586452506
L11_39 V11 V39 -2.8476115978110593e-11
C11_39 V11 V39 5.302844480641223e-20

R11_40 V11 V40 248815.22443812454
L11_40 V11 V40 -5.781974693296386e-11
C11_40 V11 V40 -1.5918733119574092e-20

R11_41 V11 V41 -30313.582762939168
L11_41 V11 V41 6.8795875596169754e-12
C11_41 V11 V41 -1.9229665464091897e-19

R11_42 V11 V42 -27022.11642329327
L11_42 V11 V42 -1.0280812389401161e-11
C11_42 V11 V42 -1.2239269245551775e-19

R11_43 V11 V43 -31049.668353185683
L11_43 V11 V43 1.9313345592368058e-11
C11_43 V11 V43 -8.36306977278012e-20

R11_44 V11 V44 -60886.046187508255
L11_44 V11 V44 2.3550954181821992e-11
C11_44 V11 V44 2.7674451112606514e-20

R11_45 V11 V45 8750.142537001406
L11_45 V11 V45 -1.0515982959544384e-11
C11_45 V11 V45 1.2739114157986214e-19

R11_46 V11 V46 14541.76001742204
L11_46 V11 V46 1.3726985295566078e-11
C11_46 V11 V46 5.491302874918186e-20

R11_47 V11 V47 31914.66497719252
L11_47 V11 V47 1.6134776873034663e-11
C11_47 V11 V47 3.0467068867910314e-20

R11_48 V11 V48 -27447.88625603375
L11_48 V11 V48 5.867819190664902e-11
C11_48 V11 V48 1.655185158534905e-22

R11_49 V11 V49 -45144.378807140616
L11_49 V11 V49 2.384931099909236e-11
C11_49 V11 V49 -3.339509986048905e-20

R11_50 V11 V50 95092.63188205422
L11_50 V11 V50 4.331706768864807e-11
C11_50 V11 V50 -2.742041465552374e-20

R11_51 V11 V51 -56376.78438138721
L11_51 V11 V51 1.898413565244848e-11
C11_51 V11 V51 1.6092162634648087e-20

R11_52 V11 V52 -62245.230780432226
L11_52 V11 V52 1.1288401889014008e-11
C11_52 V11 V52 -8.42006409172946e-20

R11_53 V11 V53 -143896.4686324027
L11_53 V11 V53 6.557248765992269e-12
C11_53 V11 V53 -5.412311423895533e-20

R11_54 V11 V54 33987.79290814862
L11_54 V11 V54 6.243580244834511e-11
C11_54 V11 V54 -4.885180702105553e-21

R11_55 V11 V55 37789.3244128809
L11_55 V11 V55 2.711520446510525e-11
C11_55 V11 V55 -2.970283486126712e-20

R11_56 V11 V56 21047.304058960002
L11_56 V11 V56 8.294639635280923e-12
C11_56 V11 V56 -4.9623390988053575e-21

R11_57 V11 V57 3559.97837155317
L11_57 V11 V57 2.129852706251592e-11
C11_57 V11 V57 2.0142123148391914e-20

R11_58 V11 V58 11115.36652310624
L11_58 V11 V58 -9.40849111947903e-12
C11_58 V11 V58 1.0410841582316464e-20

R11_59 V11 V59 43606.36351554915
L11_59 V11 V59 1.9118718286727268e-11
C11_59 V11 V59 1.4219868644951198e-20

R11_60 V11 V60 -30310.27389962387
L11_60 V11 V60 9.487190325159195e-12
C11_60 V11 V60 2.8710662857500413e-21

R11_61 V11 V61 -9347.746007708263
L11_61 V11 V61 1.138037303176593e-11
C11_61 V11 V61 -6.329255526192631e-20

R11_62 V11 V62 -7821.078717641581
L11_62 V11 V62 -1.396358421350458e-10
C11_62 V11 V62 -5.277551963869449e-20

R11_63 V11 V63 -47151.345490150314
L11_63 V11 V63 3.9956919362302307e-10
C11_63 V11 V63 -4.0431183911523916e-21

R11_64 V11 V64 88029.59998986457
L11_64 V11 V64 1.3497902924201815e-11
C11_64 V11 V64 2.7598032230687627e-21

R11_65 V11 V65 7478.89618641235
L11_65 V11 V65 7.389722158055856e-12
C11_65 V11 V65 -1.9622896093653196e-20

R11_66 V11 V66 7160.55741611303
L11_66 V11 V66 5.917275649745848e-12
C11_66 V11 V66 -1.8969310540441357e-20

R11_67 V11 V67 102598.96843904664
L11_67 V11 V67 1.4019722310596562e-11
C11_67 V11 V67 -9.938387304217306e-21

R11_68 V11 V68 -57292.79718916389
L11_68 V11 V68 2.4039762279720983e-11
C11_68 V11 V68 -4.0957549750575626e-21

R11_69 V11 V69 -50544.03165176252
L11_69 V11 V69 -3.272273405215971e-11
C11_69 V11 V69 5.121521046447325e-21

R11_70 V11 V70 -20461.34734124138
L11_70 V11 V70 -3.808510225338133e-11
C11_70 V11 V70 -9.541432123823838e-21

R11_71 V11 V71 -96163.94607480949
L11_71 V11 V71 -1.427264057345675e-10
C11_71 V11 V71 -3.0822530242948266e-21

R11_72 V11 V72 -16204.485656650966
L11_72 V11 V72 -9.421901131024495e-12
C11_72 V11 V72 1.2974755570197917e-21

R11_73 V11 V73 -32095.30417611427
L11_73 V11 V73 -4.884167812383833e-11
C11_73 V11 V73 -9.568899221647948e-21

R11_74 V11 V74 -36088.06419814913
L11_74 V11 V74 2.1017337405457563e-11
C11_74 V11 V74 1.1621972224466334e-20

R11_75 V11 V75 35449.41504062462
L11_75 V11 V75 -7.683211050980272e-11
C11_75 V11 V75 -3.60236833341968e-21

R11_76 V11 V76 39945.45592325415
L11_76 V11 V76 5.46487456711723e-12
C11_76 V11 V76 -1.220491133881073e-20

R11_77 V11 V77 57953.70299593626
L11_77 V11 V77 1.2376524791706114e-11
C11_77 V11 V77 1.208904761099139e-21

R11_78 V11 V78 -1843944.9980088514
L11_78 V11 V78 2.3676069423991597e-11
C11_78 V11 V78 -8.290733412947379e-21

R11_79 V11 V79 -54614.89014567599
L11_79 V11 V79 5.830457398640628e-12
C11_79 V11 V79 -3.806838789996178e-21

R11_80 V11 V80 -65319.38170695126
L11_80 V11 V80 -9.423715719525677e-12
C11_80 V11 V80 6.933534768025728e-21

R11_81 V11 V81 -55078.170991770894
L11_81 V11 V81 -7.578248941390803e-12
C11_81 V11 V81 -1.8092532939489722e-20

R11_82 V11 V82 162463.42673295815
L11_82 V11 V82 1.1783575572458065e-11
C11_82 V11 V82 9.620828076100813e-21

R11_83 V11 V83 196848.43928563528
L11_83 V11 V83 -2.50420269678655e-11
C11_83 V11 V83 1.7690067015781507e-20

R11_84 V11 V84 -192686.05317320503
L11_84 V11 V84 1.4748588550540836e-11
C11_84 V11 V84 6.714260948118167e-21

R11_85 V11 V85 -61703.14423955668
L11_85 V11 V85 1.6065844288359395e-11
C11_85 V11 V85 -8.751879430583194e-22

R11_86 V11 V86 -94350.3916907839
L11_86 V11 V86 -2.188862041820979e-11
C11_86 V11 V86 -2.628108428171055e-21

R11_87 V11 V87 2456641.511413836
L11_87 V11 V87 1.764020210618909e-11
C11_87 V11 V87 -9.827607846761516e-21

R11_88 V11 V88 -120699.38453103005
L11_88 V11 V88 -3.258507658739509e-11
C11_88 V11 V88 -1.1472629212053972e-20

R11_89 V11 V89 321634.6961862927
L11_89 V11 V89 1.6884115147182606e-11
C11_89 V11 V89 -4.770241237736632e-21

R11_90 V11 V90 187862.10190130008
L11_90 V11 V90 -4.544262886595155e-12
C11_90 V11 V90 -2.752201900087181e-21

R11_91 V11 V91 303449.67926730384
L11_91 V11 V91 2.6648786946186706e-11
C11_91 V11 V91 1.2978427037338279e-20

R11_92 V11 V92 202581.47422693315
L11_92 V11 V92 1.695291071769965e-11
C11_92 V11 V92 2.1372323444984533e-20

R11_93 V11 V93 -20833.221726118572
L11_93 V11 V93 3.922063573802976e-11
C11_93 V11 V93 -7.010038952391918e-21

R11_94 V11 V94 -34656.1013009758
L11_94 V11 V94 -1.2260715386035617e-11
C11_94 V11 V94 -7.998698506774131e-21

R11_95 V11 V95 -332479.59305187874
L11_95 V11 V95 5.838033515190293e-11
C11_95 V11 V95 6.4202853641205985e-21

R11_96 V11 V96 87133.16361988932
L11_96 V11 V96 2.9388418298262536e-11
C11_96 V11 V96 2.2969416020587364e-20

R11_97 V11 V97 256469.90400008467
L11_97 V11 V97 -5.469822572385762e-12
C11_97 V11 V97 -1.1519921981236544e-20

R11_98 V11 V98 41699.203104817294
L11_98 V11 V98 -3.0357448428563373e-11
C11_98 V11 V98 6.228210082448305e-21

R11_99 V11 V99 -63468.11030820014
L11_99 V11 V99 1.0044516291238175e-11
C11_99 V11 V99 -9.081906159890657e-22

R11_100 V11 V100 -1454848.7363247979
L11_100 V11 V100 -2.0592474524563426e-11
C11_100 V11 V100 -9.104546778951276e-21

R11_101 V11 V101 -69653.42250305683
L11_101 V11 V101 2.022425693024236e-11
C11_101 V11 V101 2.079413796380666e-21

R11_102 V11 V102 -5369357.72748584
L11_102 V11 V102 -2.449544412337275e-12
C11_102 V11 V102 -8.23488349756504e-21

R11_103 V11 V103 341231.86107130756
L11_103 V11 V103 4.09772838332267e-12
C11_103 V11 V103 -4.881485823748273e-21

R11_104 V11 V104 -202884.3796098752
L11_104 V11 V104 2.481283339829504e-11
C11_104 V11 V104 1.4959144234513666e-20

R11_105 V11 V105 1232852.861361585
L11_105 V11 V105 1.0364560745349826e-11
C11_105 V11 V105 -1.2053511531043e-20

R11_106 V11 V106 -105911.4326341707
L11_106 V11 V106 -8.109118326487113e-12
C11_106 V11 V106 1.9315002379944786e-20

R11_107 V11 V107 692747.5421098626
L11_107 V11 V107 -2.8784157031131578e-12
C11_107 V11 V107 2.6004274012919757e-22

R11_108 V11 V108 29816.95945219926
L11_108 V11 V108 4.3814306843573206e-12
C11_108 V11 V108 3.681415817504503e-21

R11_109 V11 V109 62790.85135301472
L11_109 V11 V109 5.832312812924972e-12
C11_109 V11 V109 2.1111690076058333e-20

R11_110 V11 V110 65381.2259914948
L11_110 V11 V110 -3.496859961425751e-11
C11_110 V11 V110 -1.1932901727405102e-20

R11_111 V11 V111 73620.94132497073
L11_111 V11 V111 5.196996133481653e-12
C11_111 V11 V111 -6.091630015662647e-21

R11_112 V11 V112 22381.076721673082
L11_112 V11 V112 -4.5593674060515765e-12
C11_112 V11 V112 -3.4449159763690884e-22

R11_113 V11 V113 39070.5153160165
L11_113 V11 V113 -9.074321422284925e-12
C11_113 V11 V113 -5.403398019666774e-21

R11_114 V11 V114 104961.35737361362
L11_114 V11 V114 -1.349472044147577e-11
C11_114 V11 V114 8.663513594029084e-21

R11_115 V11 V115 362897.1800353507
L11_115 V11 V115 -5.5206901070867835e-12
C11_115 V11 V115 3.4475172714019546e-21

R11_116 V11 V116 -223079.24315438236
L11_116 V11 V116 9.700190584451943e-12
C11_116 V11 V116 -1.1811343494394608e-21

R11_117 V11 V117 759365.5763437347
L11_117 V11 V117 1.6954942115330707e-11
C11_117 V11 V117 7.237460373081223e-21

R11_118 V11 V118 -202705.87090133372
L11_118 V11 V118 1.590909445560431e-11
C11_118 V11 V118 -3.2780303838545737e-21

R11_119 V11 V119 81731.693540309
L11_119 V11 V119 1.3574795622112479e-11
C11_119 V11 V119 -1.41385334344085e-20

R11_120 V11 V120 -233594.28560507813
L11_120 V11 V120 -5.667200224010251e-12
C11_120 V11 V120 -6.88841169507512e-21

R11_121 V11 V121 15012.441003211694
L11_121 V11 V121 -3.753616029839205e-11
C11_121 V11 V121 1.9024673272479366e-21

R11_122 V11 V122 7986.53417308301
L11_122 V11 V122 -4.077761161664985e-12
C11_122 V11 V122 3.27421990673312e-21

R11_123 V11 V123 39894.02245426048
L11_123 V11 V123 -1.496908674121646e-11
C11_123 V11 V123 -4.722480485857287e-22

R11_124 V11 V124 93787.72720744826
L11_124 V11 V124 4.767758599391338e-11
C11_124 V11 V124 -9.051068608838688e-21

R11_125 V11 V125 -15179.089815727659
L11_125 V11 V125 -1.8445622587471692e-11
C11_125 V11 V125 1.1230811972151749e-21

R11_126 V11 V126 -9942.066436362922
L11_126 V11 V126 3.093181828077965e-12
C11_126 V11 V126 3.141492342669608e-21

R11_127 V11 V127 19704.459412518518
L11_127 V11 V127 -3.7511261363008815e-12
C11_127 V11 V127 -1.9859013740434808e-21

R11_128 V11 V128 -189136.6670490562
L11_128 V11 V128 -7.361706941905581e-11
C11_128 V11 V128 -9.151091714047713e-22

R11_129 V11 V129 31231.137811329478
L11_129 V11 V129 -8.78097713596876e-12
C11_129 V11 V129 -2.8138369684884535e-21

R11_130 V11 V130 -34044.14722713249
L11_130 V11 V130 5.254229950429454e-12
C11_130 V11 V130 -3.7014363865988384e-22

R11_131 V11 V131 -22637.7958221696
L11_131 V11 V131 9.619399875906482e-11
C11_131 V11 V131 -1.7425398363536143e-22

R11_132 V11 V132 -44153.36604956152
L11_132 V11 V132 1.5185554010246426e-11
C11_132 V11 V132 -1.033471449052253e-21

R11_133 V11 V133 -60011.20102653261
L11_133 V11 V133 -7.232669005459516e-11
C11_133 V11 V133 8.942747053905238e-21

R11_134 V11 V134 -55048.328437816046
L11_134 V11 V134 3.036607979804996e-11
C11_134 V11 V134 -4.813665639397689e-21

R11_135 V11 V135 24262.09493863244
L11_135 V11 V135 -6.2119131917227645e-12
C11_135 V11 V135 9.601546142297931e-22

R11_136 V11 V136 -144546.49080901756
L11_136 V11 V136 -7.800078353114687e-11
C11_136 V11 V136 -1.1836153295003575e-21

R11_137 V11 V137 -22279.794198032312
L11_137 V11 V137 1.1328857851624422e-10
C11_137 V11 V137 -5.128812689735e-21

R11_138 V11 V138 -9782.023496602571
L11_138 V11 V138 3.2286228129871496e-12
C11_138 V11 V138 -6.0090834027571486e-21

R11_139 V11 V139 16049.666341415441
L11_139 V11 V139 -2.74453785104705e-12
C11_139 V11 V139 5.295685475465306e-21

R11_140 V11 V140 -53423.23900564074
L11_140 V11 V140 7.347452400022224e-12
C11_140 V11 V140 2.3290457829391093e-21

R11_141 V11 V141 -62036.93956163462
L11_141 V11 V141 1.3082660686948177e-11
C11_141 V11 V141 8.099666796203377e-22

R11_142 V11 V142 -43065.153114112734
L11_142 V11 V142 6.006338878013255e-12
C11_142 V11 V142 3.054722045684808e-21

R11_143 V11 V143 -49498.41353359759
L11_143 V11 V143 9.53844906443986e-12
C11_143 V11 V143 -8.047776166744293e-22

R11_144 V11 V144 37511.93723798704
L11_144 V11 V144 -1.3515484212736187e-11
C11_144 V11 V144 -2.8331652817516532e-21

R12_12 V12 0 -23640.607973659404
L12_12 V12 0 1.5021485576073963e-12
C12_12 V12 0 7.735594308056963e-22

R12_13 V12 V13 8621297.643732807
L12_13 V12 V13 1.0365601448414614e-11
C12_13 V12 V13 9.79717828524161e-22

R12_14 V12 V14 4779448.368190708
L12_14 V12 V14 -1.737460237239184e-11
C12_14 V12 V14 6.67676228163578e-22

R12_15 V12 V15 -1218976.186558653
L12_15 V12 V15 -1.180687723040122e-11
C12_15 V12 V15 -1.693769054236177e-21

R12_16 V12 V16 2270932.505000198
L12_16 V12 V16 -9.065533985774181e-12
C12_16 V12 V16 -8.233208154153766e-22

R12_17 V12 V17 -936021.569733467
L12_17 V12 V17 5.814527108199836e-11
C12_17 V12 V17 -1.750235710953841e-22

R12_18 V12 V18 -4054929.5527105923
L12_18 V12 V18 2.9970287302061905e-11
C12_18 V12 V18 1.2887822286657576e-22

R12_19 V12 V19 -417899.76829380996
L12_19 V12 V19 -4.3733828805118665e-11
C12_19 V12 V19 -4.01084141980503e-21

R12_20 V12 V20 160319.9045790304
L12_20 V12 V20 2.040905913398902e-11
C12_20 V12 V20 7.171340289749921e-21

R12_21 V12 V21 444071.0967369589
L12_21 V12 V21 1.716108946857322e-11
C12_21 V12 V21 1.6721024941655645e-21

R12_22 V12 V22 21902038.02821148
L12_22 V12 V22 1.011169584910406e-11
C12_22 V12 V22 1.9808199167338796e-22

R12_23 V12 V23 360616.9704614017
L12_23 V12 V23 4.605459557575331e-12
C12_23 V12 V23 2.586185594642888e-21

R12_24 V12 V24 -201003.48796686996
L12_24 V12 V24 -2.5691453714451578e-12
C12_24 V12 V24 -2.614355274067434e-22

R12_25 V12 V25 -589696.849666679
L12_25 V12 V25 3.254792354349582e-10
C12_25 V12 V25 1.0540189985555196e-22

R12_26 V12 V26 -4399052.282768463
L12_26 V12 V26 1.2446285649600594e-11
C12_26 V12 V26 4.312216237595408e-22

R12_27 V12 V27 -280142.41916067374
L12_27 V12 V27 1.1329361638691634e-11
C12_27 V12 V27 5.2833628362340666e-21

R12_28 V12 V28 246978.17841138912
L12_28 V12 V28 -5.222195991285966e-12
C12_28 V12 V28 -2.2618250694291193e-21

R12_29 V12 V29 -807419.0651069197
L12_29 V12 V29 2.4537780997777468e-11
C12_29 V12 V29 -5.161167052876381e-21

R12_30 V12 V30 960765.5833707284
L12_30 V12 V30 1.5975501637130797e-11
C12_30 V12 V30 -2.569569727434626e-21

R12_31 V12 V31 -1696301.9007101394
L12_31 V12 V31 9.039634634279272e-12
C12_31 V12 V31 -1.5458010853814422e-20

R12_32 V12 V32 -647754.2525292456
L12_32 V12 V32 -3.9830592375416944e-12
C12_32 V12 V32 7.639285899543515e-21

R12_33 V12 V33 -773835.5131563371
L12_33 V12 V33 -1.5311769169397508e-09
C12_33 V12 V33 4.604786242529977e-22

R12_34 V12 V34 2181915.7471370404
L12_34 V12 V34 6.427905509378844e-11
C12_34 V12 V34 -2.4348203340064504e-21

R12_35 V12 V35 -116358.33330136571
L12_35 V12 V35 -6.0674672756061584e-12
C12_35 V12 V35 1.3360546946973962e-20

R12_36 V12 V36 164011.67682859837
L12_36 V12 V36 1.1156836616017254e-11
C12_36 V12 V36 -7.268538558616846e-21

R12_37 V12 V37 -742238.5977883313
L12_37 V12 V37 1.2670875501688206e-11
C12_37 V12 V37 -1.6509004049856197e-20

R12_38 V12 V38 -145899.82693675178
L12_38 V12 V38 6.717861021889339e-11
C12_38 V12 V38 -4.038527908277357e-21

R12_39 V12 V39 -60326.0005605911
L12_39 V12 V39 8.86610051045467e-12
C12_39 V12 V39 -3.986409791976991e-20

R12_40 V12 V40 38553.18803740324
L12_40 V12 V40 -4.465289709027256e-12
C12_40 V12 V40 5.93819615003596e-20

R12_41 V12 V41 73875.71589884034
L12_41 V12 V41 -6.855870568530285e-09
C12_41 V12 V41 1.6783090184019693e-20

R12_42 V12 V42 41300.644741918535
L12_42 V12 V42 -8.049136359554988e-12
C12_42 V12 V42 4.83504966064972e-20

R12_43 V12 V43 72005.9497797636
L12_43 V12 V43 -1.4520892228395645e-11
C12_43 V12 V43 3.090724947497295e-20

R12_44 V12 V44 -24447.134109673814
L12_44 V12 V44 2.285811093618971e-12
C12_44 V12 V44 -1.1453301734769e-19

R12_45 V12 V45 -114558.99495401046
L12_45 V12 V45 1.336417922340338e-11
C12_45 V12 V45 -5.144485086953218e-20

R12_46 V12 V46 -191487.48411886048
L12_46 V12 V46 1.7815427935552892e-11
C12_46 V12 V46 1.5242934660611817e-20

R12_47 V12 V47 -385221.77775726817
L12_47 V12 V47 -2.6905086959679732e-11
C12_47 V12 V47 2.0793451889712228e-20

R12_48 V12 V48 31066.318186765773
L12_48 V12 V48 9.458402450475397e-12
C12_48 V12 V48 2.1689651993685192e-20

R12_49 V12 V49 32751.170053503254
L12_49 V12 V49 -3.360394265161059e-11
C12_49 V12 V49 2.5167965775685072e-20

R12_50 V12 V50 -32021.13726198126
L12_50 V12 V50 -3.1159813279117364e-11
C12_50 V12 V50 -1.7413388838952657e-20

R12_51 V12 V51 -278400.97856502415
L12_51 V12 V51 1.708785961420977e-11
C12_51 V12 V51 -1.4349224091723637e-20

R12_52 V12 V52 -206479.8218812349
L12_52 V12 V52 -1.0562575171983935e-10
C12_52 V12 V52 3.8513245884271646e-21

R12_53 V12 V53 108738.58980220916
L12_53 V12 V53 -1.5393696075096827e-10
C12_53 V12 V53 2.75434024202601e-20

R12_54 V12 V54 161652.9272039461
L12_54 V12 V54 -8.278584987978733e-11
C12_54 V12 V54 1.3531802306219841e-20

R12_55 V12 V55 50413.751140930835
L12_55 V12 V55 5.545759440957009e-10
C12_55 V12 V55 2.487027255268882e-20

R12_56 V12 V56 -45439.84420843517
L12_56 V12 V56 2.8961319437345526e-11
C12_56 V12 V56 -4.5225563501143355e-20

R12_57 V12 V57 -142736.15707235862
L12_57 V12 V57 -8.64739090585727e-12
C12_57 V12 V57 -4.146160163786037e-21

R12_58 V12 V58 -269161.1428513674
L12_58 V12 V58 -6.641259994819477e-12
C12_58 V12 V58 3.3397341789403665e-22

R12_59 V12 V59 -28585.868408460643
L12_59 V12 V59 -8.464031557690986e-12
C12_59 V12 V59 -7.37305677042631e-21

R12_60 V12 V60 29206.440932575355
L12_60 V12 V60 3.430886394455917e-12
C12_60 V12 V60 5.905025845171789e-21

R12_61 V12 V61 112116.67252406824
L12_61 V12 V61 -4.61389632221829e-11
C12_61 V12 V61 8.331289536382843e-21

R12_62 V12 V62 367053.9351905825
L12_62 V12 V62 1.5191336601148436e-10
C12_62 V12 V62 1.31896723714283e-20

R12_63 V12 V63 1613162.9074237633
L12_63 V12 V63 1.306053113522185e-11
C12_63 V12 V63 4.0906827359399425e-21

R12_64 V12 V64 -44934.725088399064
L12_64 V12 V64 -1.8396987815757027e-11
C12_64 V12 V64 -2.468076892277078e-20

R12_65 V12 V65 -970595.8221257352
L12_65 V12 V65 -1.1760630093107031e-11
C12_65 V12 V65 3.0347884154234383e-21

R12_66 V12 V66 -102103.48671142383
L12_66 V12 V66 -8.280012206835837e-12
C12_66 V12 V66 -7.011188162685253e-22

R12_67 V12 V67 -193331.360220296
L12_67 V12 V67 2.8509332033318156e-11
C12_67 V12 V67 1.2144081821083517e-21

R12_68 V12 V68 62658.16509074615
L12_68 V12 V68 1.1107050877956323e-11
C12_68 V12 V68 -9.833973534482188e-21

R12_69 V12 V69 313042.68107086536
L12_69 V12 V69 -1.3458914757563788e-11
C12_69 V12 V69 1.4782433544552011e-21

R12_70 V12 V70 -2215652.4144095643
L12_70 V12 V70 -1.9804653472480102e-11
C12_70 V12 V70 -1.025254847793386e-20

R12_71 V12 V71 325906.8874689599
L12_71 V12 V71 1.4894670521701563e-10
C12_71 V12 V71 -9.335634000065344e-24

R12_72 V12 V72 -321127.7526524816
L12_72 V12 V72 1.4193920213410327e-11
C12_72 V12 V72 -8.422521760405389e-21

R12_73 V12 V73 130980.63774912615
L12_73 V12 V73 -8.015460536621118e-12
C12_73 V12 V73 4.0852275763801936e-21

R12_74 V12 V74 211197.32755382775
L12_74 V12 V74 -2.6570143366823734e-11
C12_74 V12 V74 1.5622901732146566e-21

R12_75 V12 V75 -1112992.7885536705
L12_75 V12 V75 -4.778053648792196e-11
C12_75 V12 V75 2.2499889812546247e-21

R12_76 V12 V76 -423389.6618457762
L12_76 V12 V76 -2.0150615717943906e-11
C12_76 V12 V76 -8.530323757684733e-22

R12_77 V12 V77 500548.1057191185
L12_77 V12 V77 6.142747911250816e-12
C12_77 V12 V77 3.476385175903604e-22

R12_78 V12 V78 -164308.00291279698
L12_78 V12 V78 2.7463852250647476e-11
C12_78 V12 V78 -9.12466749349686e-21

R12_79 V12 V79 416041.8595679589
L12_79 V12 V79 -4.845597191865538e-11
C12_79 V12 V79 3.761311813148653e-21

R12_80 V12 V80 -1423000.223276659
L12_80 V12 V80 3.221180764078009e-12
C12_80 V12 V80 -1.1884550847266437e-21

R12_81 V12 V81 -479487.4892976567
L12_81 V12 V81 -1.350792736432294e-12
C12_81 V12 V81 -3.4198399075304575e-21

R12_82 V12 V82 88899.62272383535
L12_82 V12 V82 -7.343185603352285e-12
C12_82 V12 V82 3.850091481434998e-20

R12_83 V12 V83 99025.57380682114
L12_83 V12 V83 5.685492270689476e-12
C12_83 V12 V83 2.7021477017526214e-20

R12_84 V12 V84 1899905.259394827
L12_84 V12 V84 9.734701772521934e-12
C12_84 V12 V84 -1.7196473290852223e-22

R12_85 V12 V85 -735372.2249220574
L12_85 V12 V85 -2.0702963530558664e-11
C12_85 V12 V85 -6.84465710245755e-21

R12_86 V12 V86 -269385.13379593875
L12_86 V12 V86 1.4094565299518888e-11
C12_86 V12 V86 -1.2396186516554735e-20

R12_87 V12 V87 -182886.04697270412
L12_87 V12 V87 -6.104995608343937e-11
C12_87 V12 V87 -2.0287820333332176e-20

R12_88 V12 V88 -276636.0136021296
L12_88 V12 V88 -7.97422944820195e-12
C12_88 V12 V88 -7.168967673271193e-21

R12_89 V12 V89 311786.89406615135
L12_89 V12 V89 2.1632471009764068e-11
C12_89 V12 V89 1.0938295885783048e-20

R12_90 V12 V90 -1559886.634245631
L12_90 V12 V90 -1.459772103645854e-11
C12_90 V12 V90 -5.5671455143873276e-21

R12_91 V12 V91 81845.20432400708
L12_91 V12 V91 -2.833716683009814e-12
C12_91 V12 V91 3.0120836257569166e-20

R12_92 V12 V92 200896.4278579718
L12_92 V12 V92 1.8680035844477465e-12
C12_92 V12 V92 1.7651244859578142e-20

R12_93 V12 V93 -412448.7276331028
L12_93 V12 V93 -2.9440684957265244e-11
C12_93 V12 V93 -2.0554565347893583e-21

R12_94 V12 V94 -137259.83912307257
L12_94 V12 V94 -5.187215640459825e-12
C12_94 V12 V94 -1.3131842847900311e-20

R12_95 V12 V95 166310.12238228138
L12_95 V12 V95 -1.1577874412500875e-11
C12_95 V12 V95 1.9359212164247566e-20

R12_96 V12 V96 1271950.098692511
L12_96 V12 V96 1.3276959479080723e-12
C12_96 V12 V96 6.717477372424648e-21

R12_97 V12 V97 -336009.47777953173
L12_97 V12 V97 -4.842593631982076e-12
C12_97 V12 V97 -1.3697543808004477e-20

R12_98 V12 V98 114736.1346366097
L12_98 V12 V98 8.690626220734957e-12
C12_98 V12 V98 1.6542330805655243e-20

R12_99 V12 V99 -475277.6787789777
L12_99 V12 V99 -2.551558478711119e-11
C12_99 V12 V99 -1.742613528825442e-21

R12_100 V12 V100 -3173267.0742431236
L12_100 V12 V100 -3.9664097848936e-12
C12_100 V12 V100 -2.7300071672305894e-21

R12_101 V12 V101 200604.4496962927
L12_101 V12 V101 7.836528857798617e-12
C12_101 V12 V101 1.5905859114610245e-20

R12_102 V12 V102 219120.10543435282
L12_102 V12 V102 -7.577988757794324e-12
C12_102 V12 V102 4.266151940796367e-21

R12_103 V12 V103 187685.90679525744
L12_103 V12 V103 -4.9479320420986123e-11
C12_103 V12 V103 6.6421739864031424e-21

R12_104 V12 V104 -242532.2385661212
L12_104 V12 V104 1.843338258705744e-12
C12_104 V12 V104 -1.3342910615988486e-20

R12_105 V12 V105 -165099.12416407687
L12_105 V12 V105 -1.073201944612223e-11
C12_105 V12 V105 -1.2211765598334403e-20

R12_106 V12 V106 131548.0107184297
L12_106 V12 V106 -3.4168066375200187e-11
C12_106 V12 V106 2.865788046499334e-20

R12_107 V12 V107 3055433.902886941
L12_107 V12 V107 -1.774372383469152e-11
C12_107 V12 V107 3.410955105852601e-21

R12_108 V12 V108 514411.6452176943
L12_108 V12 V108 -5.18912047380536e-12
C12_108 V12 V108 -4.317511640073132e-21

R12_109 V12 V109 -344814.79755311494
L12_109 V12 V109 2.2910253609661664e-12
C12_109 V12 V109 -8.627818874116096e-21

R12_110 V12 V110 -189709.87426842947
L12_110 V12 V110 -2.005375952420471e-11
C12_110 V12 V110 -3.431127570151013e-20

R12_111 V12 V111 -1258975.4665198033
L12_111 V12 V111 -1.512496749266196e-11
C12_111 V12 V111 -1.0281778187743024e-20

R12_112 V12 V112 118068.02991854757
L12_112 V12 V112 4.0617046481637194e-11
C12_112 V12 V112 1.3922203337338746e-20

R12_113 V12 V113 205921.5720264015
L12_113 V12 V113 -4.594915379871749e-12
C12_113 V12 V113 1.8675727495046988e-21

R12_114 V12 V114 111548.3941364925
L12_114 V12 V114 3.198134240321762e-11
C12_114 V12 V114 2.6867689219697598e-20

R12_115 V12 V115 566232.2161078632
L12_115 V12 V115 -8.066353857872519e-11
C12_115 V12 V115 1.2398350068910457e-21

R12_116 V12 V116 -291749.4714712491
L12_116 V12 V116 -7.58786442170384e-12
C12_116 V12 V116 -7.154663873429224e-21

R12_117 V12 V117 -1913709.5221552434
L12_117 V12 V117 7.653468084812207e-12
C12_117 V12 V117 5.813271274139801e-22

R12_118 V12 V118 -164839.47341117437
L12_118 V12 V118 5.2348907530545326e-12
C12_118 V12 V118 -1.3525182575183805e-20

R12_119 V12 V119 -127890.5559269431
L12_119 V12 V119 -7.78830426612052e-12
C12_119 V12 V119 -2.749566610055661e-20

R12_120 V12 V120 193558.47876950027
L12_120 V12 V120 -4.5989952548013704e-12
C12_120 V12 V120 -6.014983052024954e-21

R12_121 V12 V121 162029.84479378504
L12_121 V12 V121 -1.1773310107049745e-11
C12_121 V12 V121 2.431019678459005e-21

R12_122 V12 V122 62869.492149679376
L12_122 V12 V122 -5.94353816829831e-12
C12_122 V12 V122 -2.453177868110426e-21

R12_123 V12 V123 152293.91147725517
L12_123 V12 V123 -2.1969922223078442e-11
C12_123 V12 V123 -5.437918256525024e-21

R12_124 V12 V124 201247.92342698816
L12_124 V12 V124 -7.886971803641032e-12
C12_124 V12 V124 -3.970905486937742e-21

R12_125 V12 V125 -248093.4899927246
L12_125 V12 V125 9.663975685028515e-11
C12_125 V12 V125 -3.3653298302991822e-21

R12_126 V12 V126 -65945.49097274199
L12_126 V12 V126 5.054397260454298e-12
C12_126 V12 V126 1.8071040877057884e-21

R12_127 V12 V127 91704.49898740402
L12_127 V12 V127 -6.068472560174111e-12
C12_127 V12 V127 -1.697704686187586e-21

R12_128 V12 V128 -656546.3862804536
L12_128 V12 V128 2.0560668017330402e-11
C12_128 V12 V128 5.076227617181673e-21

R12_129 V12 V129 90112.61565014199
L12_129 V12 V129 -8.781025450944899e-12
C12_129 V12 V129 -1.7058577605837516e-21

R12_130 V12 V130 -99940.52511324253
L12_130 V12 V130 7.487580635851458e-12
C12_130 V12 V130 8.727983361346219e-21

R12_131 V12 V131 -99436.20202499794
L12_131 V12 V131 9.485686434284375e-12
C12_131 V12 V131 5.4929783762823405e-21

R12_132 V12 V132 -206861.27755983346
L12_132 V12 V132 -8.986990114004893e-12
C12_132 V12 V132 -4.405054810527446e-22

R12_133 V12 V133 -5143736.317445722
L12_133 V12 V133 -5.3434477823704343e-11
C12_133 V12 V133 2.948986649518262e-21

R12_134 V12 V134 -280917.5483979294
L12_134 V12 V134 2.6179141420399397e-11
C12_134 V12 V134 -1.2123727732161226e-21

R12_135 V12 V135 131347.5535837114
L12_135 V12 V135 -1.062794475436946e-11
C12_135 V12 V135 2.171119283946528e-21

R12_136 V12 V136 -1088889.5390934777
L12_136 V12 V136 1.7221957804746251e-10
C12_136 V12 V136 -8.711605358200588e-21

R12_137 V12 V137 -2477782.510479055
L12_137 V12 V137 4.9481437014738254e-11
C12_137 V12 V137 -1.0143903113308187e-21

R12_138 V12 V138 -61302.16322258448
L12_138 V12 V138 7.502110107966421e-12
C12_138 V12 V138 -8.065834790683663e-21

R12_139 V12 V139 79660.3530469437
L12_139 V12 V139 -4.922432259842149e-12
C12_139 V12 V139 -3.9823398567844745e-21

R12_140 V12 V140 -124829.12464666054
L12_140 V12 V140 1.801252480854342e-11
C12_140 V12 V140 -1.9154101180969347e-21

R12_141 V12 V141 764175.200245821
L12_141 V12 V141 -9.398447106936045e-11
C12_141 V12 V141 -1.019089436357347e-20

R12_142 V12 V142 -81161.17158894667
L12_142 V12 V142 1.0143823025796358e-11
C12_142 V12 V142 -3.991151314102436e-21

R12_143 V12 V143 -178775.16994003253
L12_143 V12 V143 1.6830910851492016e-11
C12_143 V12 V143 1.263678255546368e-22

R12_144 V12 V144 202770.65300202405
L12_144 V12 V144 1.3071307273628396e-11
C12_144 V12 V144 9.888194926846249e-21

R13_13 V13 0 1042.4278463595967
L13_13 V13 0 -2.0061959773138538e-12
C13_13 V13 0 -2.19974093159774e-19

R13_14 V13 V14 -2371439.0905172452
L13_14 V13 V14 1.4052935353101109e-11
C13_14 V13 V14 2.7373957240534598e-21

R13_15 V13 V15 -304953.1535650052
L13_15 V13 V15 1.698631424853695e-11
C13_15 V13 V15 7.212036498793624e-22

R13_16 V13 V16 -826296.4409584542
L13_16 V13 V16 1.9469782181302605e-11
C13_16 V13 V16 4.41977600284143e-22

R13_17 V13 V17 -50605.74637200477
L13_17 V13 V17 8.369387103908425e-11
C13_17 V13 V17 -3.9858373338189007e-22

R13_18 V13 V18 1196861.0846230434
L13_18 V13 V18 -5.563097144857263e-11
C13_18 V13 V18 4.286268439677703e-22

R13_19 V13 V19 -85337.13852423351
L13_19 V13 V19 -7.907448291709854e-10
C13_19 V13 V19 -1.0750948018666173e-21

R13_20 V13 V20 -1318501.8747013179
L13_20 V13 V20 -4.1380575097080016e-11
C13_20 V13 V20 -2.755690565659436e-21

R13_21 V13 V21 70697.04678889315
L13_21 V13 V21 -6.028640171072361e-11
C13_21 V13 V21 -2.1083742193750186e-21

R13_22 V13 V22 -436777.18834623386
L13_22 V13 V22 -4.725295879332319e-11
C13_22 V13 V22 -1.3090232253033526e-21

R13_23 V13 V23 -684424.4757020898
L13_23 V13 V23 1.4867613224843337e-11
C13_23 V13 V23 3.0493114093434745e-22

R13_24 V13 V24 614946.1006318149
L13_24 V13 V24 6.793119947293647e-12
C13_24 V13 V24 2.732480178144469e-22

R13_25 V13 V25 -60434204.08065577
L13_25 V13 V25 -4.178520392563759e-11
C13_25 V13 V25 8.728844582556945e-21

R13_26 V13 V26 187130.64726234213
L13_26 V13 V26 -2.7242966805506543e-11
C13_26 V13 V26 -5.06811391629035e-22

R13_27 V13 V27 229351.33588131107
L13_27 V13 V27 -3.329315880097286e-10
C13_27 V13 V27 2.3847108917299546e-21

R13_28 V13 V28 979770.6941692864
L13_28 V13 V28 1.1118618321311669e-11
C13_28 V13 V28 1.4325857676096642e-21

R13_29 V13 V29 -47443.20392118497
L13_29 V13 V29 -4.0557458481763766e-11
C13_29 V13 V29 -1.0331729363863926e-20

R13_30 V13 V30 -187541.7824800828
L13_30 V13 V30 -4.2803932399579164e-11
C13_30 V13 V30 -2.0404854338495617e-21

R13_31 V13 V31 -783894.2278052863
L13_31 V13 V31 3.303022395791694e-11
C13_31 V13 V31 -6.767216538305732e-21

R13_32 V13 V32 -643853.7925590903
L13_32 V13 V32 1.0261141909367504e-11
C13_32 V13 V32 -6.320092578170997e-21

R13_33 V13 V33 -26135.432550514703
L13_33 V13 V33 5.4701923898455245e-11
C13_33 V13 V33 -1.2434002679077128e-21

R13_34 V13 V34 45441.85735790488
L13_34 V13 V34 4.980136308971512e-10
C13_34 V13 V34 1.2795211857565835e-23

R13_35 V13 V35 -40416.52032314203
L13_35 V13 V35 -6.919256708609068e-10
C13_35 V13 V35 5.856482150685382e-21

R13_36 V13 V36 129835.49450333454
L13_36 V13 V36 -3.671368715842811e-11
C13_36 V13 V36 3.8980031853608375e-21

R13_37 V13 V37 -213398.11988863302
L13_37 V13 V37 -2.71111311824504e-11
C13_37 V13 V37 -2.2752193666365886e-20

R13_38 V13 V38 263685.80153209413
L13_38 V13 V38 -4.5458801823858975e-11
C13_38 V13 V38 9.047168142085753e-21

R13_39 V13 V39 202869.7271108869
L13_39 V13 V39 -7.832346490507256e-11
C13_39 V13 V39 -2.1984241601284752e-20

R13_40 V13 V40 -62562.976134059834
L13_40 V13 V40 1.3813156364024946e-11
C13_40 V13 V40 -2.539033159363065e-20

R13_41 V13 V41 -11358.848932605606
L13_41 V13 V41 7.85626793601081e-12
C13_41 V13 V41 7.343556100821959e-20

R13_42 V13 V42 -23319.01201771564
L13_42 V13 V42 9.987166488988304e-12
C13_42 V13 V42 2.93217712522822e-20

R13_43 V13 V43 -82671.56354593758
L13_43 V13 V43 2.759728615336016e-11
C13_43 V13 V43 3.8123912789197727e-20

R13_44 V13 V44 55806.225977955466
L13_44 V13 V44 -7.898549494792072e-12
C13_44 V13 V44 2.904536078637661e-20

R13_45 V13 V45 -9879.598054771604
L13_45 V13 V45 2.0176422580026233e-11
C13_45 V13 V45 -8.390800793245623e-20

R13_46 V13 V46 -14092.638741818982
L13_46 V13 V46 -1.0303747641860303e-11
C13_46 V13 V46 1.276932782342513e-20

R13_47 V13 V47 -14568.351314673642
L13_47 V13 V47 -4.8107904176543757e-11
C13_47 V13 V47 -6.7030430490550254e-21

R13_48 V13 V48 179104.89213885448
L13_48 V13 V48 -2.983051627407492e-11
C13_48 V13 V48 -6.162337791545876e-21

R13_49 V13 V49 19554.272984900093
L13_49 V13 V49 2.870750587038308e-10
C13_49 V13 V49 2.0259762859806303e-20

R13_50 V13 V50 -26403.849032149214
L13_50 V13 V50 -3.995226885331717e-11
C13_50 V13 V50 3.2275855026517403e-21

R13_51 V13 V51 36933.988652277956
L13_51 V13 V51 -3.301110631742266e-11
C13_51 V13 V51 -2.874007115860123e-21

R13_52 V13 V52 37044.21718249889
L13_52 V13 V52 -3.4532563606190377e-11
C13_52 V13 V52 3.7810633236999997e-20

R13_53 V13 V53 -95330.43936718882
L13_53 V13 V53 -1.0023514327087627e-10
C13_53 V13 V53 8.801589304877944e-21

R13_54 V13 V54 -20064.858913434786
L13_54 V13 V54 4.87077199125997e-11
C13_54 V13 V54 -3.3272889843360232e-21

R13_55 V13 V55 -25630.37430949695
L13_55 V13 V55 -7.37444046881634e-11
C13_55 V13 V55 1.8721373563416468e-20

R13_56 V13 V56 -59458.34421162808
L13_56 V13 V56 1.9806079627546924e-10
C13_56 V13 V56 3.415604424911938e-20

R13_57 V13 V57 -2116.1426511748296
L13_57 V13 V57 7.364647463301195e-12
C13_57 V13 V57 -3.3633698353079267e-21

R13_58 V13 V58 -10946.619572766087
L13_58 V13 V58 1.0387253580159566e-11
C13_58 V13 V58 -2.7502549412613464e-21

R13_59 V13 V59 -23744.63975864747
L13_59 V13 V59 -5.667591985618775e-11
C13_59 V13 V59 -5.2369238838529535e-21

R13_60 V13 V60 -11310.435623756359
L13_60 V13 V60 -9.469703367062397e-12
C13_60 V13 V60 -2.3710189141009956e-21

R13_61 V13 V61 6375.395015719673
L13_61 V13 V61 -2.54198928570233e-10
C13_61 V13 V61 1.7541367205960942e-20

R13_62 V13 V62 7214.555217031338
L13_62 V13 V62 -2.4800183130158705e-11
C13_62 V13 V62 1.2384108564441892e-20

R13_63 V13 V63 34142.076458282005
L13_63 V13 V63 -1.0130878462514231e-10
C13_63 V13 V63 1.324257370715676e-20

R13_64 V13 V64 430889.3999384211
L13_64 V13 V64 4.1932815487445697e-11
C13_64 V13 V64 1.2287609853059497e-20

R13_65 V13 V65 -5445.889858224515
L13_65 V13 V65 -3.7718815879749105e-11
C13_65 V13 V65 3.137027600878612e-21

R13_66 V13 V66 -6560.049259202621
L13_66 V13 V66 3.1709545773530914e-11
C13_66 V13 V66 3.891956691023795e-21

R13_67 V13 V67 -22299.366764157832
L13_67 V13 V67 -3.789971438112707e-11
C13_67 V13 V67 7.571907486262926e-21

R13_68 V13 V68 -58570.10724488564
L13_68 V13 V68 -2.3951921883275416e-11
C13_68 V13 V68 8.22001425304038e-21

R13_69 V13 V69 40409.58992562811
L13_69 V13 V69 3.248370057056837e-11
C13_69 V13 V69 -3.522432472956792e-21

R13_70 V13 V70 24602.941393497156
L13_70 V13 V70 7.817495962410033e-12
C13_70 V13 V70 2.411389426855025e-21

R13_71 V13 V71 38503.14690323344
L13_71 V13 V71 2.7168744334193162e-11
C13_71 V13 V71 1.636675916376024e-21

R13_72 V13 V72 22389.437662956083
L13_72 V13 V72 1.1936701471650537e-11
C13_72 V13 V72 2.0374617427973498e-21

R13_73 V13 V73 2691591.357466151
L13_73 V13 V73 1.2766974374737474e-11
C13_73 V13 V73 4.883690922727747e-22

R13_74 V13 V74 38778.650509547435
L13_74 V13 V74 1.98432346937036e-10
C13_74 V13 V74 2.1752053064101756e-21

R13_75 V13 V75 -38245.21917566469
L13_75 V13 V75 -1.9692468363766118e-11
C13_75 V13 V75 6.913728156459703e-21

R13_76 V13 V76 -42452.138951717556
L13_76 V13 V76 4.991164766013704e-11
C13_76 V13 V76 1.2706327520317075e-21

R13_77 V13 V77 -99391.66740449994
L13_77 V13 V77 -1.2713915521604221e-11
C13_77 V13 V77 1.6418567718493636e-21

R13_78 V13 V78 -824638.3336542344
L13_78 V13 V78 3.313125392233313e-11
C13_78 V13 V78 -6.949448357593159e-21

R13_79 V13 V79 70707.79232728384
L13_79 V13 V79 2.845139957308681e-11
C13_79 V13 V79 3.964450440995773e-21

R13_80 V13 V80 75385.47832838191
L13_80 V13 V80 -9.581020759648975e-12
C13_80 V13 V80 -3.757300659924229e-21

R13_81 V13 V81 239890.67711188114
L13_81 V13 V81 3.5022930321960377e-12
C13_81 V13 V81 -2.3581876828741596e-21

R13_82 V13 V82 144615.23533758163
L13_82 V13 V82 -5.255440999469751e-12
C13_82 V13 V82 1.4503368644415013e-20

R13_83 V13 V83 143916.01014511258
L13_83 V13 V83 -4.797971625339439e-12
C13_83 V13 V83 1.087593322406086e-20

R13_84 V13 V84 -261826.48344645454
L13_84 V13 V84 -3.459164946822477e-11
C13_84 V13 V84 5.4170593887054825e-21

R13_85 V13 V85 133173.77324659206
L13_85 V13 V85 1.1128206718160104e-11
C13_85 V13 V85 -1.2833959941535539e-21

R13_86 V13 V86 -2850090.1869310024
L13_86 V13 V86 1.2940092557439337e-11
C13_86 V13 V86 -6.081796418931326e-21

R13_87 V13 V87 -262889.8279161112
L13_87 V13 V87 8.986549963876074e-12
C13_87 V13 V87 -5.150307093910866e-21

R13_88 V13 V88 160077.05349007424
L13_88 V13 V88 1.394517308817637e-11
C13_88 V13 V88 -3.563585477520424e-21

R13_89 V13 V89 -183809.13725283556
L13_89 V13 V89 -2.259566284031913e-11
C13_89 V13 V89 6.826258456759144e-22

R13_90 V13 V90 431709.6319109203
L13_90 V13 V90 2.691598378650053e-11
C13_90 V13 V90 -3.999154943078029e-21

R13_91 V13 V91 113395.5572181983
L13_91 V13 V91 -1.0033139877653678e-11
C13_91 V13 V91 1.5528155028868976e-20

R13_92 V13 V92 338027.5366183259
L13_92 V13 V92 -3.694802244903019e-12
C13_92 V13 V92 3.3066063104982146e-21

R13_93 V13 V93 20698.84916897339
L13_93 V13 V93 2.3304526351540973e-11
C13_93 V13 V93 -2.7225331820623696e-21

R13_94 V13 V94 80258.4356691187
L13_94 V13 V94 8.308171865090503e-12
C13_94 V13 V94 -7.67563137322607e-21

R13_95 V13 V95 84743.95915789506
L13_95 V13 V95 -1.1604680931110166e-11
C13_95 V13 V95 7.552271128479969e-21

R13_96 V13 V96 -319609.3656889543
L13_96 V13 V96 -3.5585708906163367e-12
C13_96 V13 V96 2.5272449317310634e-21

R13_97 V13 V97 -1789785.2730459075
L13_97 V13 V97 5.964548306900125e-12
C13_97 V13 V97 -6.62111582274533e-21

R13_98 V13 V98 -191812.16050322264
L13_98 V13 V98 -1.0354669824689189e-11
C13_98 V13 V98 3.876664508681646e-21

R13_99 V13 V99 1005997.2351094894
L13_99 V13 V99 4.671795588082681e-11
C13_99 V13 V99 -8.745675725269105e-22

R13_100 V13 V100 -215098.26456621906
L13_100 V13 V100 8.540347287844737e-12
C13_100 V13 V100 -2.9657048585755623e-21

R13_101 V13 V101 86205.39621538634
L13_101 V13 V101 -9.047213419695551e-12
C13_101 V13 V101 5.745494828378135e-21

R13_102 V13 V102 117950.96098522167
L13_102 V13 V102 2.0562286120229022e-10
C13_102 V13 V102 -4.43779970183203e-21

R13_103 V13 V103 268706.6455663418
L13_103 V13 V103 5.6963370229703115e-11
C13_103 V13 V103 4.56749292627835e-21

R13_104 V13 V104 339116.04825227347
L13_104 V13 V104 -7.109404295937129e-12
C13_104 V13 V104 8.005369453042147e-22

R13_105 V13 V105 -83902.359802154
L13_105 V13 V105 6.967364889112644e-12
C13_105 V13 V105 -1.1338092692350918e-20

R13_106 V13 V106 132469.43460559545
L13_106 V13 V106 -4.280273302700856e-12
C13_106 V13 V106 1.5554618206128833e-20

R13_107 V13 V107 -165428.77136855322
L13_107 V13 V107 -3.6254846627812536e-11
C13_107 V13 V107 -1.3483496636325557e-21

R13_108 V13 V108 -66179.95474236953
L13_108 V13 V108 8.541688813300065e-12
C13_108 V13 V108 1.6663255642352414e-21

R13_109 V13 V109 -106010.48914157659
L13_109 V13 V109 -8.39445465509932e-12
C13_109 V13 V109 3.1905503965864655e-21

R13_110 V13 V110 199982.76202635225
L13_110 V13 V110 5.038346114929516e-12
C13_110 V13 V110 -1.5993108911924666e-20

R13_111 V13 V111 -31683.406441970485
L13_111 V13 V111 9.891331143268404e-12
C13_111 V13 V111 -2.361462049337065e-21

R13_112 V13 V112 -37345.674799827444
L13_112 V13 V112 -1.8496813678400476e-11
C13_112 V13 V112 -2.1387274899561643e-21

R13_113 V13 V113 -61316.23973277627
L13_113 V13 V113 2.4543294164254584e-11
C13_113 V13 V113 2.5913717815019617e-21

R13_114 V13 V114 97062.09754336931
L13_114 V13 V114 -9.473689724207914e-12
C13_114 V13 V114 7.023334800999528e-21

R13_115 V13 V115 77916.25259254071
L13_115 V13 V115 -3.549222885960399e-11
C13_115 V13 V115 -3.9400984409053785e-21

R13_116 V13 V116 -598366.3720169317
L13_116 V13 V116 1.2016326104169257e-11
C13_116 V13 V116 1.1895133458663964e-21

R13_117 V13 V117 53569.52226669981
L13_117 V13 V117 -5.558277760088073e-11
C13_117 V13 V117 -1.1910366654900572e-21

R13_118 V13 V118 -173401.81238446597
L13_118 V13 V118 2.979282576920469e-11
C13_118 V13 V118 -8.379623921663362e-21

R13_119 V13 V119 -26018.299718966286
L13_119 V13 V119 5.9239268887392914e-12
C13_119 V13 V119 -4.769410519118096e-21

R13_120 V13 V120 14938.814152660407
L13_120 V13 V120 1.5558984314314985e-11
C13_120 V13 V120 1.1277541702129089e-21

R13_121 V13 V121 -16951.29311901696
L13_121 V13 V121 2.475565434961767e-11
C13_121 V13 V121 3.092036757999954e-21

R13_122 V13 V122 -32419.100627163378
L13_122 V13 V122 1.0909051754248477e-11
C13_122 V13 V122 4.2581305647422817e-23

R13_123 V13 V123 218530.09769386522
L13_123 V13 V123 1.9584485402880543e-11
C13_123 V13 V123 -6.948066563019824e-22

R13_124 V13 V124 -180822.253657508
L13_124 V13 V124 1.3310246161754235e-11
C13_124 V13 V124 -5.061523596605581e-22

R13_125 V13 V125 11701.213216563017
L13_125 V13 V125 -3.1645814089446674e-11
C13_125 V13 V125 -1.6966262251668982e-21

R13_126 V13 V126 -70348.00772193963
L13_126 V13 V126 -1.1414518155963634e-11
C13_126 V13 V126 -5.6230153663185e-23

R13_127 V13 V127 27106.858931908395
L13_127 V13 V127 3.263513975583385e-11
C13_127 V13 V127 4.241932335127323e-22

R13_128 V13 V128 134261.96035845598
L13_128 V13 V128 -3.00762711112693e-11
C13_128 V13 V128 -3.983037336577631e-21

R13_129 V13 V129 51755.19555365276
L13_129 V13 V129 2.0330952580054187e-11
C13_129 V13 V129 -7.329344077312519e-22

R13_130 V13 V130 -129372.06263777021
L13_130 V13 V130 -1.4641827428395093e-11
C13_130 V13 V130 -3.474536617460898e-21

R13_131 V13 V131 8901416.25239967
L13_131 V13 V131 -1.4676056452713945e-11
C13_131 V13 V131 -1.230802315321181e-21

R13_132 V13 V132 -276410.2172844068
L13_132 V13 V132 5.55585691574507e-11
C13_132 V13 V132 2.6683801192380534e-22

R13_133 V13 V133 92780.46075169004
L13_133 V13 V133 -1.0158295281993905e-11
C13_133 V13 V133 5.0904958689971174e-21

R13_134 V13 V134 -239539.14570273834
L13_134 V13 V134 -2.8200957415305023e-11
C13_134 V13 V134 -1.0107875869939438e-21

R13_135 V13 V135 59516.55520992197
L13_135 V13 V135 3.328645327999899e-11
C13_135 V13 V135 -2.3946142608735e-22

R13_136 V13 V136 162292.92530043196
L13_136 V13 V136 1.373441247685546e-10
C13_136 V13 V136 3.438779686402748e-21

R13_137 V13 V137 19401.217766720678
L13_137 V13 V137 1.5267818925737468e-10
C13_137 V13 V137 -1.885952951995313e-21

R13_138 V13 V138 -112272.61829263628
L13_138 V13 V138 -1.1150421933197628e-11
C13_138 V13 V138 3.6626376958650615e-21

R13_139 V13 V139 18497.460027691966
L13_139 V13 V139 2.275554576458741e-11
C13_139 V13 V139 1.8807289977571575e-21

R13_140 V13 V140 -109141.4999724465
L13_140 V13 V140 -5.401140827453698e-11
C13_140 V13 V140 2.1240103992999237e-21

R13_141 V13 V141 96437.16820552692
L13_141 V13 V141 1.7355931653236743e-10
C13_141 V13 V141 3.656272879008319e-21

R13_142 V13 V142 -42629.86330585466
L13_142 V13 V142 -1.901131132923307e-11
C13_142 V13 V142 -1.5684454743325992e-21

R13_143 V13 V143 -43168.02318134071
L13_143 V13 V143 -4.195977077815144e-11
C13_143 V13 V143 -8.006880013324054e-22

R13_144 V13 V144 -58279.54381286166
L13_144 V13 V144 -3.4277377629409833e-11
C13_144 V13 V144 -3.62328225795415e-21

R14_14 V14 0 2140.0223646212385
L14_14 V14 0 2.715739497386021e-12
C14_14 V14 0 1.2340677559950553e-19

R14_15 V14 V15 -9456443.108346565
L14_15 V14 V15 -9.724605083315092e-12
C14_15 V14 V15 -1.5999489143776852e-21

R14_16 V14 V16 -3194059.5698334286
L14_16 V14 V16 -1.2229279665697211e-11
C14_16 V14 V16 -1.4001717539895533e-21

R14_17 V14 V17 -376016.25345085777
L14_17 V14 V17 -1.3908793136168947e-11
C14_17 V14 V17 2.184425373460149e-22

R14_18 V14 V18 -83377704.46438342
L14_18 V14 V18 1.2529495266514333e-10
C14_18 V14 V18 -6.675694737772034e-22

R14_19 V14 V19 312767.05142770114
L14_19 V14 V19 -2.9903572768421827e-10
C14_19 V14 V19 5.12952374584745e-21

R14_20 V14 V20 312181.81695895246
L14_20 V14 V20 2.9051013114554856e-11
C14_20 V14 V20 3.609684067240819e-21

R14_21 V14 V21 -13956295.430017013
L14_21 V14 V21 -1.2710143326521473e-11
C14_21 V14 V21 -1.672131291242699e-21

R14_22 V14 V22 972746.5990670123
L14_22 V14 V22 -7.638387917727937e-12
C14_22 V14 V22 1.2361528750001829e-21

R14_23 V14 V23 -203456.89609971253
L14_23 V14 V23 -4.519635106557979e-12
C14_23 V14 V23 -1.3372667350897425e-21

R14_24 V14 V24 -340689.2525733435
L14_24 V14 V24 -7.257180556618503e-12
C14_24 V14 V24 -7.629064912186239e-22

R14_25 V14 V25 548933.9171370984
L14_25 V14 V25 4.360750166103308e-11
C14_25 V14 V25 3.143550475268768e-21

R14_26 V14 V26 -582416.4682287095
L14_26 V14 V26 -3.325073132640786e-11
C14_26 V14 V26 5.341735961956923e-21

R14_27 V14 V27 175570.8308750066
L14_27 V14 V27 -1.9101307228977238e-11
C14_27 V14 V27 -3.885381906444778e-21

R14_28 V14 V28 201100.5104756584
L14_28 V14 V28 -7.172625430299889e-12
C14_28 V14 V28 2.433973871375664e-22

R14_29 V14 V29 -255768.81777231372
L14_29 V14 V29 8.396756632319341e-10
C14_29 V14 V29 3.6661918077904836e-21

R14_30 V14 V30 332356.6837908759
L14_30 V14 V30 -2.2986478448826167e-11
C14_30 V14 V30 -1.6290655991778168e-22

R14_31 V14 V31 633066.1423362662
L14_31 V14 V31 -1.0758049617421936e-11
C14_31 V14 V31 1.4046074858268342e-20

R14_32 V14 V32 -178167.9301887796
L14_32 V14 V32 -1.0441119000122644e-11
C14_32 V14 V32 6.23268496225817e-21

R14_33 V14 V33 -160475.41593300237
L14_33 V14 V33 -5.0657165116531034e-11
C14_33 V14 V33 -5.748960630748709e-22

R14_34 V14 V34 -1340281.0544221755
L14_34 V14 V34 -4.403066813372271e-11
C14_34 V14 V34 -1.4490551928681588e-22

R14_35 V14 V35 141005.40814026745
L14_35 V14 V35 1.1020961239009066e-11
C14_35 V14 V35 -1.801510308594669e-20

R14_36 V14 V36 105716.87689175308
L14_36 V14 V36 1.1746475679614374e-10
C14_36 V14 V36 -2.8832092750699885e-21

R14_37 V14 V37 -213860.33123492077
L14_37 V14 V37 -1.2478272959665137e-11
C14_37 V14 V37 1.1416102926489373e-20

R14_38 V14 V38 -699308.5566248987
L14_38 V14 V38 -2.1213783214949734e-09
C14_38 V14 V38 -1.356606696121811e-20

R14_39 V14 V39 61248.0482223097
L14_39 V14 V39 -7.669208744229242e-12
C14_39 V14 V39 3.6882572828758674e-20

R14_40 V14 V40 78843.25089517042
L14_40 V14 V40 -1.494914093028644e-11
C14_40 V14 V40 3.254369784855657e-20

R14_41 V14 V41 -21208.52741529971
L14_41 V14 V41 1.0850883572134046e-11
C14_41 V14 V41 -1.2909635758714755e-20

R14_42 V14 V42 -27302.41973637427
L14_42 V14 V42 4.609976490577247e-12
C14_42 V14 V42 -6.51497923107848e-21

R14_43 V14 V43 -94832.83410789167
L14_43 V14 V43 1.0087165987916143e-11
C14_43 V14 V43 -4.628094546624315e-20

R14_44 V14 V44 -209930.01327215208
L14_44 V14 V44 9.43106044422268e-12
C14_44 V14 V44 -2.563496771455656e-20

R14_45 V14 V45 -143804.8268627772
L14_45 V14 V45 -3.4710121860779855e-12
C14_45 V14 V45 9.435155197799668e-20

R14_46 V14 V46 -18709.32533658267
L14_46 V14 V46 5.980861024321842e-12
C14_46 V14 V46 -7.657518730365721e-20

R14_47 V14 V47 28585.72265393003
L14_47 V14 V47 2.0015610873907546e-11
C14_47 V14 V47 -9.192029041853188e-21

R14_48 V14 V48 60785.73362478999
L14_48 V14 V48 -7.42810414147665e-11
C14_48 V14 V48 5.765211081717507e-21

R14_49 V14 V49 -30563.018663384548
L14_49 V14 V49 -5.5237216431329e-11
C14_49 V14 V49 -2.8533583310331096e-20

R14_50 V14 V50 34425.3253991182
L14_50 V14 V50 7.46022783777466e-12
C14_50 V14 V50 1.8968805513819067e-20

R14_51 V14 V51 106687.64386967619
L14_51 V14 V51 -1.9521527598175705e-11
C14_51 V14 V51 4.753059167192747e-21

R14_52 V14 V52 -138609.670072677
L14_52 V14 V52 8.427762211620242e-12
C14_52 V14 V52 -1.9460527556391028e-20

R14_53 V14 V53 45136.091993517264
L14_53 V14 V53 -2.435634846185648e-11
C14_53 V14 V53 1.2161498693941426e-20

R14_54 V14 V54 -152981.87857759045
L14_54 V14 V54 -3.210896328849473e-11
C14_54 V14 V54 5.5729081064747406e-21

R14_55 V14 V55 -21276.904685668385
L14_55 V14 V55 9.31710910178856e-12
C14_55 V14 V55 -2.772074365591629e-20

R14_56 V14 V56 -34266.9843092602
L14_56 V14 V56 -4.222018541288455e-11
C14_56 V14 V56 -3.133545751056567e-20

R14_57 V14 V57 -7721.981163531482
L14_57 V14 V57 6.757627486532424e-12
C14_57 V14 V57 -2.882083771226675e-22

R14_58 V14 V58 -7879.378882739065
L14_58 V14 V58 -2.3555542248208153e-11
C14_58 V14 V58 4.9381375673798214e-21

R14_59 V14 V59 25280.202433091945
L14_59 V14 V59 1.4961877994933352e-11
C14_59 V14 V59 9.556537035385751e-21

R14_60 V14 V60 48314.24487834056
L14_60 V14 V60 7.167447693112227e-12
C14_60 V14 V60 2.218428511535778e-21

R14_61 V14 V61 29284.038371697192
L14_61 V14 V61 -8.715624629626123e-12
C14_61 V14 V61 8.65619295023331e-22

R14_62 V14 V62 14212.23553208831
L14_62 V14 V62 1.846940494250932e-11
C14_62 V14 V62 -7.674446933857008e-21

R14_63 V14 V63 -25756.040798333797
L14_63 V14 V63 2.050713705080331e-11
C14_63 V14 V63 -8.56902460069274e-21

R14_64 V14 V64 -121740.1092695961
L14_64 V14 V64 -9.474033451171681e-12
C14_64 V14 V64 -3.367745182805476e-21

R14_65 V14 V65 -20526.860496225134
L14_65 V14 V65 8.17382298997213e-12
C14_65 V14 V65 -1.1905385280505228e-21

R14_66 V14 V66 -16540.265672523168
L14_66 V14 V66 -6.438908842790001e-12
C14_66 V14 V66 -2.5215920841772523e-21

R14_67 V14 V67 39784.233998103744
L14_67 V14 V67 3.11755610030768e-11
C14_67 V14 V67 -6.845369180711847e-21

R14_68 V14 V68 530704.7821753242
L14_68 V14 V68 1.0754045405326167e-11
C14_68 V14 V68 -5.9317313176229846e-21

R14_69 V14 V69 391198.4256618308
L14_69 V14 V69 -2.682027027679373e-11
C14_69 V14 V69 1.1662870127058192e-20

R14_70 V14 V70 64326.67706596935
L14_70 V14 V70 -3.962531839000742e-12
C14_70 V14 V70 1.4915505004548794e-20

R14_71 V14 V71 -42473.68135422847
L14_71 V14 V71 -2.3280225614480734e-11
C14_71 V14 V71 5.335970297461743e-21

R14_72 V14 V72 42714.66773063689
L14_72 V14 V72 -6.9370933422682126e-12
C14_72 V14 V72 4.953422105899413e-21

R14_73 V14 V73 106195.02668116103
L14_73 V14 V73 -1.2194872927287123e-11
C14_73 V14 V73 6.703567755834853e-21

R14_74 V14 V74 113679.72072673833
L14_74 V14 V74 -4.8769282718385556e-11
C14_74 V14 V74 -7.93542293988912e-21

R14_75 V14 V75 -72907.83570071882
L14_75 V14 V75 7.45286609309344e-12
C14_75 V14 V75 -1.9911583016621767e-20

R14_76 V14 V76 -190422.94806576843
L14_76 V14 V76 -5.1367550356938915e-12
C14_76 V14 V76 6.929886197162131e-21

R14_77 V14 V77 -184047.35710794595
L14_77 V14 V77 1.3268683751613861e-11
C14_77 V14 V77 -6.5551227301072824e-21

R14_78 V14 V78 85330.42669758161
L14_78 V14 V78 -6.193854699158868e-12
C14_78 V14 V78 2.3737144095935394e-20

R14_79 V14 V79 315317.56915431423
L14_79 V14 V79 -6.5866025173358365e-12
C14_79 V14 V79 3.9343308938399956e-21

R14_80 V14 V80 2211615.235322388
L14_80 V14 V80 4.109116634331318e-12
C14_80 V14 V80 -1.1045735368906266e-20

R14_81 V14 V81 169302.81513357963
L14_81 V14 V81 -3.203880637132555e-12
C14_81 V14 V81 1.4896971647234967e-20

R14_82 V14 V82 -71973.28646928332
L14_82 V14 V82 1.7250742067631852e-12
C14_82 V14 V82 -5.412328171657121e-20

R14_83 V14 V83 -44630.048805059356
L14_83 V14 V83 1.9228104376555756e-12
C14_83 V14 V83 -4.266628047865272e-20

R14_84 V14 V84 490436.97825027985
L14_84 V14 V84 -1.7995584131179807e-11
C14_84 V14 V84 7.367433281580324e-22

R14_85 V14 V85 109257.71109342856
L14_85 V14 V85 -3.4684397877249834e-12
C14_85 V14 V85 2.1495424069958045e-20

R14_86 V14 V86 72400.61231764819
L14_86 V14 V86 -3.9309374386333586e-12
C14_86 V14 V86 2.0418867478775497e-20

R14_87 V14 V87 109468.19018798969
L14_87 V14 V87 -2.453918209031785e-12
C14_87 V14 V87 2.819117091715811e-20

R14_88 V14 V88 100281.66087096436
L14_88 V14 V88 -6.698515223251851e-12
C14_88 V14 V88 1.1000759224047624e-20

R14_89 V14 V89 -167787.65066386285
L14_89 V14 V89 5.073815952523997e-12
C14_89 V14 V89 -2.0277007598526457e-20

R14_90 V14 V90 -82956.36288136791
L14_90 V14 V90 1.1279572741237092e-11
C14_90 V14 V90 -6.630517747432392e-21

R14_91 V14 V91 -50745.05173351256
L14_91 V14 V91 2.101237432558368e-12
C14_91 V14 V91 -4.8739491044467663e-20

R14_92 V14 V92 -86841.5898223096
L14_92 V14 V92 2.2128908299915293e-12
C14_92 V14 V92 -2.7738763978108797e-20

R14_93 V14 V93 49483.24744532353
L14_93 V14 V93 -8.461027023569123e-12
C14_93 V14 V93 5.041168335389605e-21

R14_94 V14 V94 31084.828240101462
L14_94 V14 V94 -4.121807635000396e-12
C14_94 V14 V94 2.477034353125862e-20

R14_95 V14 V95 -76610.95734027485
L14_95 V14 V95 3.675630154698491e-12
C14_95 V14 V95 -2.853462264414405e-20

R14_96 V14 V96 -134121.86193785715
L14_96 V14 V96 2.918711870204996e-12
C14_96 V14 V96 -2.0891220348041013e-20

R14_97 V14 V97 -227749.73964636648
L14_97 V14 V97 -6.122567278741262e-12
C14_97 V14 V97 1.4241467315059673e-20

R14_98 V14 V98 -34412.02670916928
L14_98 V14 V98 2.6785363121966867e-12
C14_98 V14 V98 -2.473584135728998e-20

R14_99 V14 V99 42317.022201328036
L14_99 V14 V99 -1.008647942938609e-11
C14_99 V14 V99 5.513984019280124e-21

R14_100 V14 V100 288534.12289555836
L14_100 V14 V100 -5.867004642607832e-12
C14_100 V14 V100 8.680346019284501e-21

R14_101 V14 V101 -5888849.691043046
L14_101 V14 V101 2.6871657651965326e-12
C14_101 V14 V101 -3.16163845573176e-20

R14_102 V14 V102 -56855.6399884491
L14_102 V14 V102 2.377138920066388e-12
C14_102 V14 V102 -2.5128804565323097e-20

R14_103 V14 V103 -593018.0063155364
L14_103 V14 V103 -6.8638643211738315e-12
C14_103 V14 V103 6.723956287997949e-21

R14_104 V14 V104 200120.51721677222
L14_104 V14 V104 1.7713992639240644e-11
C14_104 V14 V104 -7.91745124358124e-21

R14_105 V14 V105 85584.83650688593
L14_105 V14 V105 -2.1505167806025688e-12
C14_105 V14 V105 3.9530822861975e-20

R14_106 V14 V106 -114235.59031565161
L14_106 V14 V106 1.3585513320552521e-12
C14_106 V14 V106 -6.475977410207187e-20

R14_107 V14 V107 -273842.4337961047
L14_107 V14 V107 2.9211637106790743e-12
C14_107 V14 V107 -2.0726261363007447e-20

R14_108 V14 V108 -68432.9213827049
L14_108 V14 V108 -2.263081900128324e-12
C14_108 V14 V108 2.3824148289539424e-20

R14_109 V14 V109 -162729.96930012116
L14_109 V14 V109 -6.484194528974268e-11
C14_109 V14 V109 -1.8071789538418626e-23

R14_110 V14 V110 -74477.46779729321
L14_110 V14 V110 -1.6871681730579923e-12
C14_110 V14 V110 6.243632167276357e-20

R14_111 V14 V111 60278.43787270118
L14_111 V14 V111 -3.1577109825530605e-12
C14_111 V14 V111 1.8967588796533638e-20

R14_112 V14 V112 -20795.070899595983
L14_112 V14 V112 2.1342353432051492e-12
C14_112 V14 V112 -2.185973340000018e-20

R14_113 V14 V113 -38455.19225927863
L14_113 V14 V113 6.686602478439132e-12
C14_113 V14 V113 -1.3384323492214596e-20

R14_114 V14 V114 -48901.31054009504
L14_114 V14 V114 2.65818156853158e-12
C14_114 V14 V114 -3.2609537219374054e-20

R14_115 V14 V115 -63564.549734633765
L14_115 V14 V115 5.625748750201271e-12
C14_115 V14 V115 -8.611471595558665e-21

R14_116 V14 V116 62417.562887412096
L14_116 V14 V116 -3.3560333813304444e-12
C14_116 V14 V116 1.6666806222329152e-20

R14_117 V14 V117 -154283.41928845897
L14_117 V14 V117 -7.672217680359975e-12
C14_117 V14 V117 1.5385992989399855e-20

R14_118 V14 V118 64231.00938882463
L14_118 V14 V118 -3.2942307093604124e-12
C14_118 V14 V118 2.7523438880005376e-20

R14_119 V14 V119 57033.691262916254
L14_119 V14 V119 -2.2514708061268637e-12
C14_119 V14 V119 3.288195526052928e-20

R14_120 V14 V120 -17657.704993805804
L14_120 V14 V120 -1.8902769683566923e-11
C14_120 V14 V120 6.161955456762839e-21

R14_121 V14 V121 -27360.70603664111
L14_121 V14 V121 9.078108191246806e-12
C14_121 V14 V121 -8.686027446764892e-21

R14_122 V14 V122 -7383.879729327963
L14_122 V14 V122 7.087805705989097e-12
C14_122 V14 V122 -9.06713747906186e-22

R14_123 V14 V123 -37548.59396167637
L14_123 V14 V123 -2.6440616541683326e-11
C14_123 V14 V123 4.534242326606915e-21

R14_124 V14 V124 3746443.136513094
L14_124 V14 V124 -8.491015684512896e-12
C14_124 V14 V124 8.475300872376318e-21

R14_125 V14 V125 65382.516013486405
L14_125 V14 V125 -8.84166931713311e-12
C14_125 V14 V125 5.919882620887182e-21

R14_126 V14 V126 6727.645039301962
L14_126 V14 V126 -8.606471038857867e-12
C14_126 V14 V126 -3.779295066691291e-21

R14_127 V14 V127 -9901.60671652684
L14_127 V14 V127 6.124612658639151e-12
C14_127 V14 V127 2.0312967016514217e-21

R14_128 V14 V128 -354284.86612622923
L14_128 V14 V128 1.4215742322595663e-11
C14_128 V14 V128 7.839671715059779e-21

R14_129 V14 V129 -23705.22693098725
L14_129 V14 V129 7.065130833175469e-11
C14_129 V14 V129 7.67583210159209e-21

R14_130 V14 V130 26566.63349716529
L14_130 V14 V130 -2.229384259794275e-11
C14_130 V14 V130 1.1871463651185441e-20

R14_131 V14 V131 22543.00315826894
L14_131 V14 V131 1.0808492895123972e-11
C14_131 V14 V131 -5.4739798759755675e-21

R14_132 V14 V132 35093.39547162318
L14_132 V14 V132 -2.506048163516199e-11
C14_132 V14 V132 2.8227643446393626e-21

R14_133 V14 V133 114755.75727304508
L14_133 V14 V133 4.242572584073614e-12
C14_133 V14 V133 -1.6797320960582694e-20

R14_134 V14 V134 45163.195273399215
L14_134 V14 V134 -4.973312061323487e-11
C14_134 V14 V134 1.5734181599618058e-21

R14_135 V14 V135 -13936.602776512851
L14_135 V14 V135 1.553079618545369e-11
C14_135 V14 V135 1.264261013893714e-21

R14_136 V14 V136 291568.1928447369
L14_136 V14 V136 -3.540733080039542e-11
C14_136 V14 V136 -4.99765642420499e-21

R14_137 V14 V137 59964.8296530753
L14_137 V14 V137 -7.893179588710298e-12
C14_137 V14 V137 8.266454888629799e-21

R14_138 V14 V138 7497.571454748392
L14_138 V14 V138 -1.0890661674868193e-11
C14_138 V14 V138 1.642504883005439e-21

R14_139 V14 V139 -7597.375433225062
L14_139 V14 V139 4.660372122712758e-12
C14_139 V14 V139 -5.1878862051269796e-21

R14_140 V14 V140 26675.416328254327
L14_140 V14 V140 -7.93052084737261e-12
C14_140 V14 V140 -1.3988118128947116e-21

R14_141 V14 V141 33708.0573980239
L14_141 V14 V141 -1.3289739873588736e-11
C14_141 V14 V141 -7.365514924431129e-22

R14_142 V14 V142 25044.745070873734
L14_142 V14 V142 -1.6802613725776414e-11
C14_142 V14 V142 6.767033801533971e-21

R14_143 V14 V143 24081.520091007296
L14_143 V14 V143 -8.791044484398638e-11
C14_143 V14 V143 3.2641553802564835e-21

R14_144 V14 V144 -38604.108146152605
L14_144 V14 V144 9.658057006954162e-12
C14_144 V14 V144 -5.197672368120803e-22

R15_15 V15 0 6877.1483144401955
L15_15 V15 0 2.048323035719436e-12
C15_15 V15 0 -3.963372609776708e-20

R15_16 V15 V16 1801109.499652636
L15_16 V15 V16 -1.610325306409354e-11
C15_16 V15 V16 -6.050635905298295e-22

R15_17 V15 V17 -100639.38234339314
L15_17 V15 V17 -3.8381181131093307e-11
C15_17 V15 V17 -9.734677048941862e-22

R15_18 V15 V18 454778.3550982397
L15_18 V15 V18 9.882583280645252e-11
C15_18 V15 V18 1.4319925944902821e-21

R15_19 V15 V19 -121203.5415420341
L15_19 V15 V19 1.631228107133048e-10
C15_19 V15 V19 2.515436113915703e-21

R15_20 V15 V20 188482.47050815137
L15_20 V15 V20 3.9421630320551237e-11
C15_20 V15 V20 3.0669285651912222e-21

R15_21 V15 V21 115620.91814619975
L15_21 V15 V21 -1.0772503030005033e-10
C15_21 V15 V21 3.213887787389535e-22

R15_22 V15 V22 -407774.20714750537
L15_22 V15 V22 -7.370556415126168e-11
C15_22 V15 V22 8.518515771895548e-22

R15_23 V15 V23 -2661722.850607697
L15_23 V15 V23 -9.071790656100708e-12
C15_23 V15 V23 -1.5287409398398107e-21

R15_24 V15 V24 -585017.439280914
L15_24 V15 V24 -6.903206734443321e-12
C15_24 V15 V24 -6.469083017969223e-22

R15_25 V15 V25 -333377.5529935249
L15_25 V15 V25 6.774503974920731e-11
C15_25 V15 V25 5.629913727698169e-21

R15_26 V15 V26 206493.72537913424
L15_26 V15 V26 5.226547301000308e-11
C15_26 V15 V26 2.9144315866066807e-22

R15_27 V15 V27 1054960.0614218607
L15_27 V15 V27 -6.170231009542506e-11
C15_27 V15 V27 8.009853884828881e-22

R15_28 V15 V28 400851.1246413139
L15_28 V15 V28 -9.612744748031159e-12
C15_28 V15 V28 -1.9251135695931036e-22

R15_29 V15 V29 -130124.71971019276
L15_29 V15 V29 2.9692911800016896e-11
C15_29 V15 V29 -8.538762655566504e-21

R15_30 V15 V30 -110804.50570136584
L15_30 V15 V30 7.660614124841655e-11
C15_30 V15 V30 -1.9817573038413852e-21

R15_31 V15 V31 -199591.1401913198
L15_31 V15 V31 -2.9769393646365525e-11
C15_31 V15 V31 3.2538975588505343e-21

R15_32 V15 V32 -992392.4494303131
L15_32 V15 V32 -1.0642593151435834e-11
C15_32 V15 V32 2.5440510725928e-21

R15_33 V15 V33 -43019.98590043547
L15_33 V15 V33 -5.449338186862624e-11
C15_33 V15 V33 5.05570336540942e-21

R15_34 V15 V34 59156.584980505344
L15_34 V15 V34 -1.8946838077263003e-10
C15_34 V15 V34 -2.9224751228568188e-21

R15_35 V15 V35 -50507.421957049984
L15_35 V15 V35 5.5074523103859076e-11
C15_35 V15 V35 -3.754250497748586e-21

R15_36 V15 V36 115542.07064297626
L15_36 V15 V36 4.751185881629643e-11
C15_36 V15 V36 -2.658161594918923e-21

R15_37 V15 V37 -274845.7603958385
L15_37 V15 V37 -3.7038282696002097e-11
C15_37 V15 V37 -1.8976332663517376e-20

R15_38 V15 V38 381357.77526959596
L15_38 V15 V38 4.386782948292606e-11
C15_38 V15 V38 -1.2888204241031118e-23

R15_39 V15 V39 134952.30645556666
L15_39 V15 V39 -2.4890130625191732e-11
C15_39 V15 V39 -6.858853553275678e-21

R15_40 V15 V40 92417.59940091088
L15_40 V15 V40 -1.385301437101384e-11
C15_40 V15 V40 2.606555924987065e-20

R15_41 V15 V41 -28905.137185836047
L15_41 V15 V41 2.0426553244595834e-10
C15_41 V15 V41 6.310049877907413e-20

R15_42 V15 V42 89766.22148664217
L15_42 V15 V42 2.49901225821539e-10
C15_42 V15 V42 3.011266060759194e-20

R15_43 V15 V43 -33636.591808398436
L15_43 V15 V43 2.3884715176698316e-11
C15_43 V15 V43 3.329626322398369e-20

R15_44 V15 V44 -81957.36157075052
L15_44 V15 V44 8.121732386103393e-12
C15_44 V15 V44 -2.737768517807152e-20

R15_45 V15 V45 -22849.585542088716
L15_45 V15 V45 -7.982304746581783e-12
C15_45 V15 V45 -1.1741597052256223e-20

R15_46 V15 V46 -24065.268204419644
L15_46 V15 V46 8.587036196063998e-12
C15_46 V15 V46 -4.062058586414181e-20

R15_47 V15 V47 -10796.54331553677
L15_47 V15 V47 4.36647623498652e-11
C15_47 V15 V47 -3.101189233189555e-20

R15_48 V15 V48 -459734.8864814765
L15_48 V15 V48 4.988112509490548e-11
C15_48 V15 V48 -3.1422289110986853e-21

R15_49 V15 V49 32744.254983491137
L15_49 V15 V49 -3.599708857656543e-11
C15_49 V15 V49 -6.914388247929259e-22

R15_50 V15 V50 -98282.2254526404
L15_50 V15 V50 1.713103446182184e-11
C15_50 V15 V50 1.599388217059798e-20

R15_51 V15 V51 85976.98672447956
L15_51 V15 V51 -2.4760044662478555e-11
C15_51 V15 V51 2.3148357466142136e-21

R15_52 V15 V52 40998.55069244029
L15_52 V15 V52 7.129943315890504e-11
C15_52 V15 V52 1.9809052536546783e-20

R15_53 V15 V53 -159335.0457188085
L15_53 V15 V53 -2.5498227716899442e-11
C15_53 V15 V53 2.1313617753909526e-20

R15_54 V15 V54 -41784.87554896622
L15_54 V15 V54 -3.861029127147246e-11
C15_54 V15 V54 -1.443104482572589e-21

R15_55 V15 V55 -101487.11051111876
L15_55 V15 V55 2.1613319814568506e-11
C15_55 V15 V55 -9.55175333418503e-22

R15_56 V15 V56 -30313.542751295023
L15_56 V15 V56 -5.469294812705151e-11
C15_56 V15 V56 -2.4989230339055163e-20

R15_57 V15 V57 -3922.9516762164503
L15_57 V15 V57 6.962545786973293e-11
C15_57 V15 V57 -3.661991514995118e-21

R15_58 V15 V58 10179.356409845874
L15_58 V15 V58 -8.405200149241196e-12
C15_58 V15 V58 -5.5256560626418486e-21

R15_59 V15 V59 -38848.783733617965
L15_59 V15 V59 6.932783661310009e-11
C15_59 V15 V59 -4.2343479847869455e-21

R15_60 V15 V60 -44781.008266458935
L15_60 V15 V60 8.53900762554958e-12
C15_60 V15 V60 4.597113279340276e-22

R15_61 V15 V61 11680.368756677495
L15_61 V15 V61 -1.6916058538622673e-11
C15_61 V15 V61 1.4413712700701884e-20

R15_62 V15 V62 17418.362240071776
L15_62 V15 V62 3.5413025993465124e-11
C15_62 V15 V62 1.9526770327929426e-20

R15_63 V15 V63 12968.343782625732
L15_63 V15 V63 9.219810525113449e-11
C15_63 V15 V63 -1.2094954643849616e-20

R15_64 V15 V64 -471977.16373018967
L15_64 V15 V64 -1.7665619445413728e-11
C15_64 V15 V64 -1.3406702151725552e-20

R15_65 V15 V65 -11729.028009204938
L15_65 V15 V65 -2.7251009683022927e-10
C15_65 V15 V65 6.191306639723286e-21

R15_66 V15 V66 -24989.412335144516
L15_66 V15 V66 -1.0398645769355426e-11
C15_66 V15 V66 4.395448837580131e-22

R15_67 V15 V67 -11915.192866054105
L15_67 V15 V67 -1.8923978279076008e-11
C15_67 V15 V67 2.737462202101143e-22

R15_68 V15 V68 -143533.99203758204
L15_68 V15 V68 2.5499636619065705e-11
C15_68 V15 V68 -3.935605211444257e-21

R15_69 V15 V69 -71494.39874020175
L15_69 V15 V69 -2.655329419724321e-11
C15_69 V15 V69 3.871732503438722e-21

R15_70 V15 V70 30837.851791290184
L15_70 V15 V70 -1.2002336974864289e-11
C15_70 V15 V70 -4.385641546512741e-22

R15_71 V15 V71 16316.345349284
L15_71 V15 V71 7.675774277831223e-12
C15_71 V15 V71 2.6616711736186282e-21

R15_72 V15 V72 2167418.7699205913
L15_72 V15 V72 -1.2263562219444537e-11
C15_72 V15 V72 -8.509386695235167e-22

R15_73 V15 V73 -82806.57491773092
L15_73 V15 V73 -1.0125286844839986e-11
C15_73 V15 V73 4.877297204994358e-21

R15_74 V15 V74 -167834.57011975022
L15_74 V15 V74 5.41370714468583e-10
C15_74 V15 V74 -9.131835201574557e-21

R15_75 V15 V75 -72543.47125201364
L15_75 V15 V75 2.57534771885568e-11
C15_75 V15 V75 -3.3545491104154086e-21

R15_76 V15 V76 -70913.52700252313
L15_76 V15 V76 -1.3523825215161395e-11
C15_76 V15 V76 -2.1270397604416872e-21

R15_77 V15 V77 -296196.41804596345
L15_77 V15 V77 1.4094792483172055e-11
C15_77 V15 V77 -2.6435584478825358e-21

R15_78 V15 V78 -563869.3263387379
L15_78 V15 V78 -1.3051331886381844e-11
C15_78 V15 V78 1.0025769408416357e-20

R15_79 V15 V79 470645.62219029426
L15_79 V15 V79 -2.9249951537543243e-11
C15_79 V15 V79 -1.2073068825148548e-20

R15_80 V15 V80 99826.22117812686
L15_80 V15 V80 6.836452417727848e-12
C15_80 V15 V80 8.869723924707e-21

R15_81 V15 V81 230052.0267810271
L15_81 V15 V81 -3.629600405132966e-12
C15_81 V15 V81 7.930485052089381e-21

R15_82 V15 V82 -130613.02992645005
L15_82 V15 V82 3.823171943995798e-12
C15_82 V15 V82 -1.4270831901701385e-20

R15_83 V15 V83 89947.86523849687
L15_83 V15 V83 3.0863926498691423e-12
C15_83 V15 V83 -6.237532134316275e-21

R15_84 V15 V84 -67894.43281363639
L15_84 V15 V84 1.0158289267552783e-10
C15_84 V15 V84 -7.792956608318889e-21

R15_85 V15 V85 -3165696.8279124917
L15_85 V15 V85 -8.20365560282321e-12
C15_85 V15 V85 -2.187454936602378e-21

R15_86 V15 V86 -106389.39735503879
L15_86 V15 V86 -6.9263308172180905e-12
C15_86 V15 V86 5.038016261805601e-21

R15_87 V15 V87 -210831.05691376762
L15_87 V15 V87 -5.515314003841884e-12
C15_87 V15 V87 5.199710482214539e-22

R15_88 V15 V88 552465.633348399
L15_88 V15 V88 -9.69486278405248e-12
C15_88 V15 V88 5.740584099946728e-21

R15_89 V15 V89 -150962.0643877711
L15_89 V15 V89 1.0406655105854166e-11
C15_89 V15 V89 -3.218751537260804e-21

R15_90 V15 V90 41405.27417252859
L15_90 V15 V90 -7.26280052996313e-11
C15_90 V15 V90 1.1803456953178076e-20

R15_91 V15 V91 310533.9810418967
L15_91 V15 V91 5.038434648079072e-12
C15_91 V15 V91 -1.432616684306973e-20

R15_92 V15 V92 -2189512.308609516
L15_92 V15 V92 3.156676647912494e-12
C15_92 V15 V92 -4.668116139663407e-21

R15_93 V15 V93 40614.023553588384
L15_93 V15 V93 -2.1557712442011374e-11
C15_93 V15 V93 5.992690386400673e-23

R15_94 V15 V94 -93299.01807190965
L15_94 V15 V94 -5.736959125747263e-12
C15_94 V15 V94 1.1513074255913628e-20

R15_95 V15 V95 83947.85666009085
L15_95 V15 V95 7.583771350555265e-12
C15_95 V15 V95 -7.178877474349069e-21

R15_96 V15 V96 -1138296.028508259
L15_96 V15 V96 3.496812470400636e-12
C15_96 V15 V96 -4.994177930063775e-21

R15_97 V15 V97 62998.02522293064
L15_97 V15 V97 -6.063306288881173e-12
C15_97 V15 V97 1.2812689546381187e-20

R15_98 V15 V98 62033.72480471747
L15_98 V15 V98 5.302821099925015e-12
C15_98 V15 V98 -1.1647544708691339e-21

R15_99 V15 V99 -34773.82936473609
L15_99 V15 V99 -3.303581099684311e-11
C15_99 V15 V99 -1.2757473813033218e-21

R15_100 V15 V100 -259297.21513508013
L15_100 V15 V100 -7.614162615036902e-12
C15_100 V15 V100 5.060405905812529e-21

R15_101 V15 V101 -353125.76430977025
L15_101 V15 V101 5.028064789267058e-12
C15_101 V15 V101 -6.639545733169116e-21

R15_102 V15 V102 33301.55433194516
L15_102 V15 V102 1.1589991800474872e-11
C15_102 V15 V102 2.2776614083379072e-20

R15_103 V15 V103 -160796.94154618657
L15_103 V15 V103 -5.99940905271071e-11
C15_103 V15 V103 -1.5302266349505722e-20

R15_104 V15 V104 -150800.41526601388
L15_104 V15 V104 8.769397037563921e-12
C15_104 V15 V104 -6.08195975731707e-21

R15_105 V15 V105 -166888.32227921204
L15_105 V15 V105 -4.611626802483025e-12
C15_105 V15 V105 6.603446312476342e-21

R15_106 V15 V106 -97273.4263698626
L15_106 V15 V106 2.958945582571862e-12
C15_106 V15 V106 -6.6283195043349405e-21

R15_107 V15 V107 -349440.9350107926
L15_107 V15 V107 1.115229988227242e-11
C15_107 V15 V107 2.0807526504771337e-20

R15_108 V15 V108 119613.18225391408
L15_108 V15 V108 -5.529551629140718e-12
C15_108 V15 V108 -1.630082532305107e-20

R15_109 V15 V109 -109972.53019379104
L15_109 V15 V109 1.023026215594322e-11
C15_109 V15 V109 -1.481365131536394e-20

R15_110 V15 V110 19907.4819032914
L15_110 V15 V110 -3.3140290718568325e-12
C15_110 V15 V110 1.1201166109368612e-20

R15_111 V15 V111 -19727.330565441996
L15_111 V15 V111 -7.942580737403418e-12
C15_111 V15 V111 -6.121258460133808e-21

R15_112 V15 V112 37582.39174703648
L15_112 V15 V112 5.910515825130894e-12
C15_112 V15 V112 1.1498414721463732e-20

R15_113 V15 V113 50805.159228572666
L15_113 V15 V113 1.195675943849993e-10
C15_113 V15 V113 2.0469023538845395e-21

R15_114 V15 V114 71524.38565400825
L15_114 V15 V114 5.813495268676073e-12
C15_114 V15 V114 -3.971573664756138e-21

R15_115 V15 V115 31461.85455185623
L15_115 V15 V115 1.6748360060176223e-11
C15_115 V15 V115 1.2040438873508464e-20

R15_116 V15 V116 -50608.67541159647
L15_116 V15 V116 -7.550160759146845e-12
C15_116 V15 V116 -8.217213300264529e-21

R15_117 V15 V117 33151.89892524715
L15_117 V15 V117 -4.05009712962812e-11
C15_117 V15 V117 -4.2245852589613725e-21

R15_118 V15 V118 -70161.41938899124
L15_118 V15 V118 -9.80030591341782e-12
C15_118 V15 V118 2.6360854034583967e-21

R15_119 V15 V119 -24461.768506787823
L15_119 V15 V119 -4.464710858555695e-12
C15_119 V15 V119 1.8274522005086763e-21

R15_120 V15 V120 6743.58400720024
L15_120 V15 V120 -1.0692109175188519e-11
C15_120 V15 V120 -2.11429442677445e-21

R15_121 V15 V121 -56295.655388201965
L15_121 V15 V121 3.489665385187475e-11
C15_121 V15 V121 -2.4649553786505263e-21

R15_122 V15 V122 6791.172978824413
L15_122 V15 V122 -3.358186007318257e-11
C15_122 V15 V122 -3.0341391430603555e-21

R15_123 V15 V123 30743.087619364283
L15_123 V15 V123 -2.4286130206298185e-11
C15_123 V15 V123 8.09452683894136e-22

R15_124 V15 V124 -86541.74040179326
L15_124 V15 V124 -1.3287828783857e-11
C15_124 V15 V124 1.3900396435353194e-21

R15_125 V15 V125 14316.757817904772
L15_125 V15 V125 -1.9050663034098352e-11
C15_125 V15 V125 -1.83162530645692e-21

R15_126 V15 V126 -4644.4123135993705
L15_126 V15 V126 1.6701436520661892e-11
C15_126 V15 V126 3.246752324854746e-22

R15_127 V15 V127 5650.362465610847
L15_127 V15 V127 -1.0684478893024776e-10
C15_127 V15 V127 1.3765818027740684e-21

R15_128 V15 V128 57001.96992874588
L15_128 V15 V128 2.3023848170311603e-11
C15_128 V15 V128 5.644541099511044e-21

R15_129 V15 V129 15115.27912927328
L15_129 V15 V129 -3.5286801022861834e-11
C15_129 V15 V129 4.8401724130325135e-21

R15_130 V15 V130 -24242.179333361553
L15_130 V15 V130 2.0974679578596427e-11
C15_130 V15 V130 7.634670289981988e-23

R15_131 V15 V131 -20553.933490157848
L15_131 V15 V131 1.3452044635801177e-11
C15_131 V15 V131 4.561474264006029e-21

R15_132 V15 V132 -23663.888238319883
L15_132 V15 V132 -5.485551855417673e-11
C15_132 V15 V132 1.3287102593903302e-21

R15_133 V15 V133 -207748.66362580637
L15_133 V15 V133 8.69425578662799e-12
C15_133 V15 V133 -3.5038423727942515e-21

R15_134 V15 V134 -32437.155718173795
L15_134 V15 V134 1.3313648631126524e-10
C15_134 V15 V134 1.6246396899244422e-21

R15_135 V15 V135 8707.864027570318
L15_135 V15 V135 -3.340854711755201e-11
C15_135 V15 V135 -2.794593582558535e-21

R15_136 V15 V136 167220.03888238774
L15_136 V15 V136 -6.429032075142172e-11
C15_136 V15 V136 -5.2891491774980754e-21

R15_137 V15 V137 31317.098145052976
L15_137 V15 V137 -2.2319713340528877e-11
C15_137 V15 V137 1.5298124178402947e-21

R15_138 V15 V138 -5551.963550610495
L15_138 V15 V138 1.6465041745891424e-11
C15_138 V15 V138 -5.046602061316736e-22

R15_139 V15 V139 4313.033460811168
L15_139 V15 V139 -9.105130996946347e-11
C15_139 V15 V139 -5.168915963976154e-22

R15_140 V15 V140 -18242.877559274482
L15_140 V15 V140 -4.928036042625744e-11
C15_140 V15 V140 -4.7193369105677086e-21

R15_141 V15 V141 -29470.475409266626
L15_141 V15 V141 -4.1535900820087853e-11
C15_141 V15 V141 -3.4142783941409695e-21

R15_142 V15 V142 -16530.456591665352
L15_142 V15 V142 3.578328021667037e-11
C15_142 V15 V142 2.2482236160732285e-22

R15_143 V15 V143 -13072.036414463688
L15_143 V15 V143 3.4463322133189573e-11
C15_143 V15 V143 4.27028831499385e-22

R15_144 V15 V144 63395.08687643072
L15_144 V15 V144 1.9967541711641717e-11
C15_144 V15 V144 4.671875105295509e-21

R16_16 V16 0 2614.0455561163267
L16_16 V16 0 2.8661444492459008e-12
C16_16 V16 0 -5.0536662008114167e-20

R16_17 V16 V17 -306533.26886005467
L16_17 V16 V17 -4.298390506693427e-11
C16_17 V16 V17 -8.528776233208277e-22

R16_18 V16 V18 3589021.5358439
L16_18 V16 V18 1.0331311946364563e-10
C16_18 V16 V18 -3.6866132256702235e-22

R16_19 V16 V19 422391.2167989607
L16_19 V16 V19 -1.0854124479144052e-10
C16_19 V16 V19 2.6439642086622454e-22

R16_20 V16 V20 -138622.05977994128
L16_20 V16 V20 2.66884726218773e-11
C16_20 V16 V20 2.616031833901306e-21

R16_21 V16 V21 532315.5938489676
L16_21 V16 V21 -1.7977889875482448e-10
C16_21 V16 V21 1.2021307174274958e-21

R16_22 V16 V22 -8386366.386964154
L16_22 V16 V22 -2.5584633757504077e-11
C16_22 V16 V22 -3.065999697983342e-22

R16_23 V16 V23 -278076.1990672358
L16_23 V16 V23 -5.485457606919079e-11
C16_23 V16 V23 3.2894350699691583e-22

R16_24 V16 V24 -368204.46161944885
L16_24 V16 V24 -6.4732984055992225e-12
C16_24 V16 V24 -3.474196888324639e-22

R16_25 V16 V25 13642280.624077715
L16_25 V16 V25 9.696047254151579e-11
C16_25 V16 V25 1.4229810738817616e-21

R16_26 V16 V26 -2417472.3133141375
L16_26 V16 V26 8.565187762597563e-10
C16_26 V16 V26 2.235717757775199e-21

R16_27 V16 V27 217219.75173484726
L16_27 V16 V27 2.7624942021340454e-10
C16_27 V16 V27 -1.49990882848146e-21

R16_28 V16 V28 211718.30865506188
L16_28 V16 V28 -9.144250349081178e-12
C16_28 V16 V28 8.564016313573782e-22

R16_29 V16 V29 -270553.9455441337
L16_29 V16 V29 5.108622643335154e-11
C16_29 V16 V29 -3.1974393377890172e-21

R16_30 V16 V30 1760610.527530904
L16_30 V16 V30 -1.958608815107416e-10
C16_30 V16 V30 -5.056275959013372e-22

R16_31 V16 V31 466020.91359188285
L16_31 V16 V31 -1.3977451721172305e-10
C16_31 V16 V31 -2.893539591628953e-22

R16_32 V16 V32 -503673.3474435813
L16_32 V16 V32 -1.0489691092647499e-11
C16_32 V16 V32 1.7289040520117177e-21

R16_33 V16 V33 1889864.144078723
L16_33 V16 V33 -5.589418111376252e-11
C16_33 V16 V33 2.0165187484011187e-21

R16_34 V16 V34 -669096.3117018279
L16_34 V16 V34 -2.7591838117107985e-10
C16_34 V16 V34 -1.5986016515619442e-21

R16_35 V16 V35 97297.17252062575
L16_35 V16 V35 -7.017338552649535e-11
C16_35 V16 V35 -1.5708302202251954e-21

R16_36 V16 V36 -84262.75901063893
L16_36 V16 V36 4.1766966470566075e-11
C16_36 V16 V36 -9.636116959517941e-22

R16_37 V16 V37 -71694.2966089482
L16_37 V16 V37 -1.5411058379534065e-10
C16_37 V16 V37 -6.814939244750224e-21

R16_38 V16 V38 545387.3970101626
L16_38 V16 V38 -2.7955489292310284e-10
C16_38 V16 V38 -4.377624296601123e-21

R16_39 V16 V39 -478085.61147495575
L16_39 V16 V39 -5.1624619637714237e-11
C16_39 V16 V39 -1.0043179177279327e-22

R16_40 V16 V40 128278.78437310169
L16_40 V16 V40 -1.3735953609629059e-11
C16_40 V16 V40 1.2802531630665702e-20

R16_41 V16 V41 -94947.09449500474
L16_41 V16 V41 4.5355919663553374e-11
C16_41 V16 V41 2.5717127022440657e-20

R16_42 V16 V42 -118645.26018174141
L16_42 V16 V42 2.070365358616076e-11
C16_42 V16 V42 2.1249186233279284e-20

R16_43 V16 V43 125969.90349890696
L16_43 V16 V43 6.193079160619171e-11
C16_43 V16 V43 -4.5907300439614365e-21

R16_44 V16 V44 -36223.95807625031
L16_44 V16 V44 6.594072055132444e-12
C16_44 V16 V44 -1.4276109184122225e-20

R16_45 V16 V45 -49761.873169448656
L16_45 V16 V45 -1.1791166057425056e-11
C16_45 V16 V45 9.745907361487291e-22

R16_46 V16 V46 -47241.60350478082
L16_46 V16 V46 1.2695448661023133e-11
C16_46 V16 V46 -2.811018187338678e-20

R16_47 V16 V47 52728.2161266165
L16_47 V16 V47 9.109422872270159e-11
C16_47 V16 V47 5.036758311820448e-22

R16_48 V16 V48 -43713.40256083282
L16_48 V16 V48 7.268860706088256e-11
C16_48 V16 V48 3.1187221474116478e-21

R16_49 V16 V49 -51503.586523252205
L16_49 V16 V49 -5.475333054608247e-11
C16_49 V16 V49 6.993843194054122e-22

R16_50 V16 V50 50272.33691389282
L16_50 V16 V50 2.701007652955928e-11
C16_50 V16 V50 6.547041713493962e-21

R16_51 V16 V51 -330966.395996642
L16_51 V16 V51 5.560287204657675e-09
C16_51 V16 V51 -3.1385893493044058e-21

R16_52 V16 V52 105065.159678434
L16_52 V16 V52 2.8630953507400106e-11
C16_52 V16 V52 7.599610148182613e-21

R16_53 V16 V53 501978.51165868156
L16_53 V16 V53 -2.6635823876467918e-11
C16_53 V16 V53 1.3008544627350253e-20

R16_54 V16 V54 -139968.03745705166
L16_54 V16 V54 -5.015920282595846e-11
C16_54 V16 V54 3.84116261476239e-21

R16_55 V16 V55 -44934.593010266806
L16_55 V16 V55 2.8412623206866085e-11
C16_55 V16 V55 -2.0003076135957656e-21

R16_56 V16 V56 84732.69780839817
L16_56 V16 V56 6.78652250396118e-11
C16_56 V16 V56 -5.24160861935179e-21

R16_57 V16 V57 -13765.61941203629
L16_57 V16 V57 4.893363227303323e-11
C16_57 V16 V57 -3.2301774737397556e-21

R16_58 V16 V58 -13787.561386351748
L16_58 V16 V58 -1.9849931184841402e-11
C16_58 V16 V58 1.5158753006138988e-21

R16_59 V16 V59 32151.83087798225
L16_59 V16 V59 -1.1600658532952709e-09
C16_59 V16 V59 1.7044856133670956e-21

R16_60 V16 V60 -12391.856557390032
L16_60 V16 V60 7.70460519752002e-12
C16_60 V16 V60 1.2105890720669663e-21

R16_61 V16 V61 36350.48894568533
L16_61 V16 V61 -1.722385560165461e-11
C16_61 V16 V61 1.1205251912994231e-20

R16_62 V16 V62 29494.17845180955
L16_62 V16 V62 4.206329342512287e-11
C16_62 V16 V62 5.088787652296667e-21

R16_63 V16 V63 -45533.17687105166
L16_63 V16 V63 2.1113004549795224e-11
C16_63 V16 V63 4.7957436632855515e-21

R16_64 V16 V64 -39640685.243909754
L16_64 V16 V64 -1.48381098333975e-11
C16_64 V16 V64 4.034839628909289e-21

R16_65 V16 V65 -28098.72323214919
L16_65 V16 V65 1.2386244330139204e-10
C16_65 V16 V65 3.04785852368977e-21

R16_66 V16 V66 -21481.12592835967
L16_66 V16 V66 -7.973198151137684e-12
C16_66 V16 V66 8.817055214145504e-22

R16_67 V16 V67 68334.6538263136
L16_67 V16 V67 3.8829459018048933e-11
C16_67 V16 V67 3.046060706309602e-22

R16_68 V16 V68 -35946.24072342287
L16_68 V16 V68 1.4229931408613688e-11
C16_68 V16 V68 -1.3066515237822968e-21

R16_69 V16 V69 80971.24825831655
L16_69 V16 V69 -2.9233602757488944e-11
C16_69 V16 V69 5.4436225286288085e-21

R16_70 V16 V70 108573.01092508517
L16_70 V16 V70 -9.658988574548006e-12
C16_70 V16 V70 3.7317914487731036e-21

R16_71 V16 V71 -112283.43981279687
L16_71 V16 V71 -4.0348683163305186e-11
C16_71 V16 V71 2.897872826534933e-21

R16_72 V16 V72 42686.37961640685
L16_72 V16 V72 -5.3984249137070065e-11
C16_72 V16 V72 -7.049893746390805e-22

R16_73 V16 V73 1908051.3543177214
L16_73 V16 V73 -1.8988880762249875e-11
C16_73 V16 V73 4.0198881763848684e-21

R16_74 V16 V74 124965.02749219502
L16_74 V16 V74 -5.980083503809383e-11
C16_74 V16 V74 -2.261060362752234e-21

R16_75 V16 V75 -132611.84912537358
L16_75 V16 V75 2.282972420835811e-11
C16_75 V16 V75 -5.451862660136467e-21

R16_76 V16 V76 -260788.91891078744
L16_76 V16 V76 -9.206523206800597e-12
C16_76 V16 V76 4.848128747782447e-21

R16_77 V16 V77 -1271370.4610140526
L16_77 V16 V77 1.481312906719408e-11
C16_77 V16 V77 -2.2186521225557153e-21

R16_78 V16 V78 371399.9888350588
L16_78 V16 V78 -1.7573129574231994e-11
C16_78 V16 V78 4.598168599138376e-21

R16_79 V16 V79 173635.0255945
L16_79 V16 V79 -1.3800213710551155e-11
C16_79 V16 V79 7.231337126470443e-21

R16_80 V16 V80 615751.9845685336
L16_80 V16 V80 5.3707417277792566e-12
C16_80 V16 V80 -7.596951363420338e-21

R16_81 V16 V81 1514333.250482467
L16_81 V16 V81 -3.16686999925657e-12
C16_81 V16 V81 3.6366720650333026e-21

R16_82 V16 V82 -345702.1559880429
L16_82 V16 V82 5.5869703802404915e-12
C16_82 V16 V82 -4.22479215838597e-21

R16_83 V16 V83 -201082.58442336743
L16_83 V16 V83 3.9857176565924126e-12
C16_83 V16 V83 -7.11980484576535e-21

R16_84 V16 V84 184824.8807638031
L16_84 V16 V84 9.736381763911946e-11
C16_84 V16 V84 2.174308108797127e-21

R16_85 V16 V85 189971.07323301325
L16_85 V16 V85 -8.03171895236749e-12
C16_85 V16 V85 7.340304740741867e-21

R16_86 V16 V86 373173.53962649056
L16_86 V16 V86 -1.3658792381560443e-11
C16_86 V16 V86 2.1946706847737195e-21

R16_87 V16 V87 530337.5182399122
L16_87 V16 V87 -6.071742975510033e-12
C16_87 V16 V87 3.777761487757736e-21

R16_88 V16 V88 267517.47847922205
L16_88 V16 V88 -1.102179577284004e-11
C16_88 V16 V88 6.800120600056725e-22

R16_89 V16 V89 -1623762.9623822558
L16_89 V16 V89 1.2256015555932268e-11
C16_89 V16 V89 -2.4942795028511233e-21

R16_90 V16 V90 -115455.31903992099
L16_90 V16 V90 3.652350536422674e-11
C16_90 V16 V90 -8.996467368672738e-21

R16_91 V16 V91 -512224.0212395451
L16_91 V16 V91 1.1901083777776277e-11
C16_91 V16 V91 -4.254504472722676e-21

R16_92 V16 V92 -332474.6958982454
L16_92 V16 V92 3.154163720083555e-12
C16_92 V16 V92 -4.426876956107112e-21

R16_93 V16 V93 88200.4081015831
L16_93 V16 V93 -1.7190869104595963e-11
C16_93 V16 V93 1.9663366916892836e-21

R16_94 V16 V94 80001.84547913603
L16_94 V16 V94 -7.0989371605050415e-12
C16_94 V16 V94 2.0727196191450786e-21

R16_95 V16 V95 -347530.73026057053
L16_95 V16 V95 1.274636568771192e-11
C16_95 V16 V95 -2.8868378700601593e-21

R16_96 V16 V96 -4899631.254052135
L16_96 V16 V96 2.94984632792244e-12
C16_96 V16 V96 -6.080798500078355e-21

R16_97 V16 V97 -213672.18705630937
L16_97 V16 V97 -9.329688387044873e-12
C16_97 V16 V97 -2.428534755620621e-21

R16_98 V16 V98 -85211.28321573237
L16_98 V16 V98 5.684112391305322e-12
C16_98 V16 V98 -4.2522818533428086e-21

R16_99 V16 V99 84763.63189584867
L16_99 V16 V99 -1.786447446235971e-11
C16_99 V16 V99 1.962173888023838e-21

R16_100 V16 V100 507140.1106326309
L16_100 V16 V100 -7.56320220518168e-12
C16_100 V16 V100 -1.4906229385161132e-22

R16_101 V16 V101 315896.50746420224
L16_101 V16 V101 5.8095391107185646e-12
C16_101 V16 V101 -4.318036966206822e-21

R16_102 V16 V102 -112529.28119605134
L16_102 V16 V102 6.6259211804642234e-12
C16_102 V16 V102 -1.6368937056491596e-20

R16_103 V16 V103 226042.33276973703
L16_103 V16 V103 -1.3125184643490418e-11
C16_103 V16 V103 1.1185368056198092e-20

R16_104 V16 V104 1255100.634338248
L16_104 V16 V104 6.009841293086859e-12
C16_104 V16 V104 -6.798819501840831e-21

R16_105 V16 V105 326510.677230906
L16_105 V16 V105 -4.71408683894003e-12
C16_105 V16 V105 9.330478438621153e-21

R16_106 V16 V106 499029.2916553091
L16_106 V16 V106 3.5314900409596203e-12
C16_106 V16 V106 -1.4257699689478196e-20

R16_107 V16 V107 -258313.0637184416
L16_107 V16 V107 7.226332344617325e-12
C16_107 V16 V107 -1.450430905520762e-20

R16_108 V16 V108 -208163.79278021873
L16_108 V16 V108 -4.2945878978727194e-12
C16_108 V16 V108 1.1104693689160314e-20

R16_109 V16 V109 -169537.29547787787
L16_109 V16 V109 1.0278623088804478e-11
C16_109 V16 V109 1.6506246013704764e-21

R16_110 V16 V110 -81949.74751893498
L16_110 V16 V110 -4.206281978725858e-12
C16_110 V16 V110 1.0685860446211937e-20

R16_111 V16 V111 100713.69721850712
L16_111 V16 V111 -6.612438481638615e-12
C16_111 V16 V111 6.667706926729854e-21

R16_112 V16 V112 -40714.03790124886
L16_112 V16 V112 4.995093456352467e-12
C16_112 V16 V112 -6.765800555806106e-21

R16_113 V16 V113 -86781.34116144197
L16_113 V16 V113 1.5652009317737801e-10
C16_113 V16 V113 -5.7526475214168835e-21

R16_114 V16 V114 -4867674.774439133
L16_114 V16 V114 6.322695307124173e-12
C16_114 V16 V114 -3.1051902102821893e-21

R16_115 V16 V115 -120654.21692335566
L16_115 V16 V115 1.3263451468765463e-11
C16_115 V16 V115 -7.545283603421306e-21

R16_116 V16 V116 113903.71418576934
L16_116 V16 V116 -6.581630762880248e-12
C16_116 V16 V116 7.059041626694576e-21

R16_117 V16 V117 -287791.8338060558
L16_117 V16 V117 -5.211341705493679e-11
C16_117 V16 V117 7.719547698016337e-21

R16_118 V16 V118 219365.90763745023
L16_118 V16 V118 -1.4572811684790548e-11
C16_118 V16 V118 5.220526982458068e-21

R16_119 V16 V119 497565.01161002455
L16_119 V16 V119 -4.774367038137767e-12
C16_119 V16 V119 3.469952756371529e-21

R16_120 V16 V120 -34257.35995312768
L16_120 V16 V120 -1.598297111530644e-11
C16_120 V16 V120 1.293424200167727e-21

R16_121 V16 V121 -53052.03627986469
L16_121 V16 V121 4.6109869352098157e-11
C16_121 V16 V121 -1.9717559546313433e-21

R16_122 V16 V122 -14846.776916124316
L16_122 V16 V122 4.531601742502148e-11
C16_122 V16 V122 -5.779345413572672e-22

R16_123 V16 V123 -171168.1171331788
L16_123 V16 V123 -4.248555624377394e-11
C16_123 V16 V123 1.0013049303558001e-22

R16_124 V16 V124 175142.30463808659
L16_124 V16 V124 -1.3822848991747543e-11
C16_124 V16 V124 2.0456467685645057e-21

R16_125 V16 V125 110635.77248726605
L16_125 V16 V125 -2.8718991276825367e-11
C16_125 V16 V125 1.5146347034010525e-21

R16_126 V16 V126 13159.212510864641
L16_126 V16 V126 -8.80421869315142e-11
C16_126 V16 V126 -1.4602188775788149e-21

R16_127 V16 V127 -18847.71431102903
L16_127 V16 V127 2.7736532901579357e-11
C16_127 V16 V127 -6.433690587823296e-23

R16_128 V16 V128 -301213.45929254004
L16_128 V16 V128 2.986925568997517e-11
C16_128 V16 V128 3.6092004389248966e-21

R16_129 V16 V129 -80871.71701311211
L16_129 V16 V129 -5.973269241364477e-11
C16_129 V16 V129 2.0019233656641144e-21

R16_130 V16 V130 131258.71336018003
L16_130 V16 V130 3.48695611560118e-10
C16_130 V16 V130 7.3978017521128e-21

R16_131 V16 V131 80657.28294688404
L16_131 V16 V131 1.5891682334038758e-11
C16_131 V16 V131 -2.39440839657578e-21

R16_132 V16 V132 80074.048270885
L16_132 V16 V132 -2.0987693219275883e-11
C16_132 V16 V132 1.6140410219887188e-21

R16_133 V16 V133 198681.2120001316
L16_133 V16 V133 1.1533336028704916e-11
C16_133 V16 V133 -3.805445371773146e-21

R16_134 V16 V134 101120.8597591152
L16_134 V16 V134 1.3169352560892857e-09
C16_134 V16 V134 -1.2894647580050835e-22

R16_135 V16 V135 -27599.509990234037
L16_135 V16 V135 9.068323748216007e-11
C16_135 V16 V135 1.7324370199473275e-21

R16_136 V16 V136 584981.3096052577
L16_136 V16 V136 -1.0856954209713037e-10
C16_136 V16 V136 -3.7768875129395985e-21

R16_137 V16 V137 96881.06846475886
L16_137 V16 V137 -2.377300035844041e-11
C16_137 V16 V137 1.1571672962429403e-21

R16_138 V16 V138 16123.584895418415
L16_138 V16 V138 -5.847149408274656e-11
C16_138 V16 V138 -6.072180861943939e-22

R16_139 V16 V139 -14592.350427111014
L16_139 V16 V139 1.9508639927689654e-11
C16_139 V16 V139 -3.33534125707156e-21

R16_140 V16 V140 59289.966805686556
L16_140 V16 V140 -2.1599046895617116e-11
C16_140 V16 V140 -5.181969296120573e-22

R16_141 V16 V141 51071.248197149354
L16_141 V16 V141 -2.939860121171831e-11
C16_141 V16 V141 -2.1557135882795902e-21

R16_142 V16 V142 89751.13075455154
L16_142 V16 V142 -1.1228569247791169e-10
C16_142 V16 V142 1.3004869055995848e-21

R16_143 V16 V143 52858.13899290527
L16_143 V16 V143 1.5922807055136643e-10
C16_143 V16 V143 1.5906880965626861e-21

R16_144 V16 V144 -83153.34368381382
L16_144 V16 V144 1.51458913617699e-11
C16_144 V16 V144 1.3706868861231027e-21

R17_17 V17 0 313.7235474937221
L17_17 V17 0 -9.656080081481408e-13
C17_17 V17 0 -2.9219120956714713e-19

R17_18 V17 V18 423288.77430436265
L17_18 V17 V18 -8.166121110922177e-11
C17_18 V17 V18 1.004817090114282e-21

R17_19 V17 V19 -33270.66546738268
L17_19 V17 V19 -5.269214270683375e-11
C17_19 V17 V19 4.06242234030263e-21

R17_20 V17 V20 203671.20573500026
L17_20 V17 V20 9.017309542938649e-11
C17_20 V17 V20 -7.237551055113562e-22

R17_21 V17 V21 24950.992453404
L17_21 V17 V21 -6.990350695527097e-12
C17_21 V17 V21 -1.0914381500890043e-20

R17_22 V17 V22 -210380.3011423485
L17_22 V17 V22 -1.1847122471392417e-11
C17_22 V17 V22 5.386589002180889e-22

R17_23 V17 V23 -109874.52412033924
L17_23 V17 V23 -1.47163679741597e-11
C17_23 V17 V23 -5.599487441954029e-22

R17_24 V17 V24 -868894.5970249383
L17_24 V17 V24 2.2892575730858506e-10
C17_24 V17 V24 3.8875607927415985e-22

R17_25 V17 V25 140407.22476092965
L17_25 V17 V25 -2.2869512451395944e-11
C17_25 V17 V25 3.0585088622140576e-20

R17_26 V17 V26 63010.07015893743
L17_26 V17 V26 -2.5294209444696502e-11
C17_26 V17 V26 5.694357958904901e-21

R17_27 V17 V27 51884.04233089696
L17_27 V17 V27 -2.9573673709584974e-11
C17_27 V17 V27 3.851622982248275e-21

R17_28 V17 V28 100232.20281754764
L17_28 V17 V28 -2.5264892517410144e-11
C17_28 V17 V28 3.0561681451133702e-21

R17_29 V17 V29 -14049.956102720904
L17_29 V17 V29 -1.7721780166578602e-11
C17_29 V17 V29 -2.1637059228716453e-20

R17_30 V17 V30 -63782.03721437432
L17_30 V17 V30 -2.5064415391435625e-11
C17_30 V17 V30 -9.214245170626653e-21

R17_31 V17 V31 -150742.11680202885
L17_31 V17 V31 -4.524606349758196e-11
C17_31 V17 V31 -2.1304346752569005e-21

R17_32 V17 V32 -106139.13655297413
L17_32 V17 V32 -4.9594495094703264e-09
C17_32 V17 V32 -6.3918724093612164e-21

R17_33 V17 V33 -8613.759343988173
L17_33 V17 V33 2.5259916991094298e-11
C17_33 V17 V33 -1.0661153202754517e-20

R17_34 V17 V34 15578.485794576776
L17_34 V17 V34 -4.05895902295155e-11
C17_34 V17 V34 3.542375925336976e-21

R17_35 V17 V35 -15657.11765388192
L17_35 V17 V35 1.5971000113667272e-11
C17_35 V17 V35 -7.543498656646766e-21

R17_36 V17 V36 32577.905390015163
L17_36 V17 V36 -5.287783515084648e-11
C17_36 V17 V36 4.6466869263161085e-21

R17_37 V17 V37 -183940.31778965954
L17_37 V17 V37 -5.225068598643196e-12
C17_37 V17 V37 -4.229452282184339e-20

R17_38 V17 V38 283685.38144885836
L17_38 V17 V38 -4.2757708243409383e-11
C17_38 V17 V38 5.986788042526573e-22

R17_39 V17 V39 22233.852547400784
L17_39 V17 V39 -5.67921989458976e-12
C17_39 V17 V39 -1.4044300315825913e-20

R17_40 V17 V40 -89288.88464812683
L17_40 V17 V40 -1.3158595767316353e-10
C17_40 V17 V40 -2.3031175949574365e-21

R17_41 V17 V41 -3028.282243555327
L17_41 V17 V41 1.9273256879496756e-12
C17_41 V17 V41 1.4999464336830534e-19

R17_42 V17 V42 -6669.035695651582
L17_42 V17 V42 2.0886202906081548e-12
C17_42 V17 V42 8.598911409348751e-20

R17_43 V17 V43 -15035.5410122656
L17_43 V17 V43 4.60602347341987e-12
C17_43 V17 V43 4.584582783102362e-20

R17_44 V17 V44 58630.39617982806
L17_44 V17 V44 5.6325745544960766e-11
C17_44 V17 V44 4.916344977864845e-21

R17_45 V17 V45 -3580.594375576005
L17_45 V17 V45 -3.7847550005382285e-12
C17_45 V17 V45 -1.0577908848439431e-19

R17_46 V17 V46 -3855.231401494678
L17_46 V17 V46 5.2164497411718664e-11
C17_46 V17 V46 -6.143533488880592e-20

R17_47 V17 V47 -5767.005528929073
L17_47 V17 V47 4.935677865313733e-11
C17_47 V17 V47 -2.4101909975233024e-20

R17_48 V17 V48 33531.130709242316
L17_48 V17 V48 -1.844431806582806e-11
C17_48 V17 V48 -5.301571134233831e-21

R17_49 V17 V49 8756.502270967483
L17_49 V17 V49 -5.625709044273312e-11
C17_49 V17 V49 1.8442165716300574e-20

R17_50 V17 V50 -13771.053633679778
L17_50 V17 V50 9.106530257104974e-12
C17_50 V17 V50 2.6156798818443556e-20

R17_51 V17 V51 11217.626409435421
L17_51 V17 V51 -8.645694682272137e-12
C17_51 V17 V51 -1.2973184425714738e-20

R17_52 V17 V52 12393.319135716303
L17_52 V17 V52 9.500385835607717e-12
C17_52 V17 V52 6.514569934131264e-20

R17_53 V17 V53 7451042.485728563
L17_53 V17 V53 -2.8569735537033138e-11
C17_53 V17 V53 3.448254469236449e-20

R17_54 V17 V54 -7098.137449730232
L17_54 V17 V54 5.865393462313197e-11
C17_54 V17 V54 4.140618335505414e-21

R17_55 V17 V55 -6324.407385933704
L17_55 V17 V55 8.222688981900417e-12
C17_55 V17 V55 1.4963349987931256e-20

R17_56 V17 V56 -10877.54211853688
L17_56 V17 V56 2.638910150424976e-11
C17_56 V17 V56 2.0626903661414724e-20

R17_57 V17 V57 -680.7471054170351
L17_57 V17 V57 1.867667522445381e-12
C17_57 V17 V57 -2.238032351940135e-21

R17_58 V17 V58 -2974.9374937632274
L17_58 V17 V58 9.890455032463201e-12
C17_58 V17 V58 -4.496262583701182e-21

R17_59 V17 V59 -13868.791098713746
L17_59 V17 V59 9.460564833341472e-11
C17_59 V17 V59 -5.297266544189147e-21

R17_60 V17 V60 -4509.43784702542
L17_60 V17 V60 1.2857070189735307e-11
C17_60 V17 V60 -1.8200230757396857e-21

R17_61 V17 V61 2128.949659245185
L17_61 V17 V61 -6.923942488037013e-12
C17_61 V17 V61 3.0691618279450575e-20

R17_62 V17 V62 2180.888529478419
L17_62 V17 V62 -2.6838076260706897e-11
C17_62 V17 V62 2.5088530247546794e-20

R17_63 V17 V63 22628.222670474
L17_63 V17 V63 1.3345481646215336e-11
C17_63 V17 V63 1.0360015171109575e-20

R17_64 V17 V64 -74119.72078917279
L17_64 V17 V64 -1.3070369219814819e-11
C17_64 V17 V64 7.94369436712024e-21

R17_65 V17 V65 -1849.971056328686
L17_65 V17 V65 1.0295842361539548e-11
C17_65 V17 V65 4.6157362254090115e-21

R17_66 V17 V66 -2148.92092033897
L17_66 V17 V66 -9.056762107751026e-12
C17_66 V17 V66 -2.9664037862017e-21

R17_67 V17 V67 -9983.675213342463
L17_67 V17 V67 -1.2717989976432923e-10
C17_67 V17 V67 5.112345764370642e-21

R17_68 V17 V68 -23436.71404310732
L17_68 V17 V68 1.528929347293113e-11
C17_68 V17 V68 7.715739653267194e-21

R17_69 V17 V69 16166.954275317104
L17_69 V17 V69 -7.38225839718588e-11
C17_69 V17 V69 6.524631979103525e-21

R17_70 V17 V70 9216.296880468251
L17_70 V17 V70 -4.989065165127016e-11
C17_70 V17 V70 1.1199454013464503e-20

R17_71 V17 V71 51419.826478497154
L17_71 V17 V71 1.4259476902473919e-11
C17_71 V17 V71 9.155561306214142e-21

R17_72 V17 V72 7529.635754761659
L17_72 V17 V72 4.9609485988982605e-11
C17_72 V17 V72 8.760065640350201e-21

R17_73 V17 V73 100546.56075081299
L17_73 V17 V73 3.0345193142073764e-11
C17_73 V17 V73 9.635936051853429e-21

R17_74 V17 V74 13038.58948977033
L17_74 V17 V74 -3.0571806911097155e-10
C17_74 V17 V74 -7.815827165762964e-22

R17_75 V17 V75 -12225.016484529255
L17_75 V17 V75 3.770483771357623e-11
C17_75 V17 V75 -2.7653928404578357e-21

R17_76 V17 V76 -15399.503697908289
L17_76 V17 V76 -6.546020195773418e-12
C17_76 V17 V76 1.6111397065915798e-21

R17_77 V17 V77 -39339.301215786436
L17_77 V17 V77 -5.093734432066725e-10
C17_77 V17 V77 -2.3311856692931918e-21

R17_78 V17 V78 82671.22314356585
L17_78 V17 V78 -9.44513481524927e-12
C17_78 V17 V78 2.941279515219588e-21

R17_79 V17 V79 30528.59068635611
L17_79 V17 V79 -2.0546302556346e-11
C17_79 V17 V79 -1.2326135109228046e-22

R17_80 V17 V80 28294.540543520983
L17_80 V17 V80 6.705365715964396e-12
C17_80 V17 V80 -6.731350982300897e-21

R17_81 V17 V81 113670.77731620432
L17_81 V17 V81 -2.4606639151742982e-11
C17_81 V17 V81 4.600346344487776e-21

R17_82 V17 V82 67894.4132257714
L17_82 V17 V82 4.132944018186531e-12
C17_82 V17 V82 -5.70807328234045e-21

R17_83 V17 V83 -161264.17479998656
L17_83 V17 V83 4.518176671919388e-12
C17_83 V17 V83 5.294702244998036e-21

R17_84 V17 V84 -89887.33537914508
L17_84 V17 V84 -1.3837931610804251e-11
C17_84 V17 V84 1.167705176176128e-20

R17_85 V17 V85 44185.112083101034
L17_85 V17 V85 -7.202749525522111e-12
C17_85 V17 V85 9.790409503167291e-21

R17_86 V17 V86 73887.98376449493
L17_86 V17 V86 -7.7780383440555e-12
C17_86 V17 V86 7.739926342514204e-22

R17_87 V17 V87 -182384.5713553726
L17_87 V17 V87 -4.2966815547367855e-12
C17_87 V17 V87 7.544216148368646e-22

R17_88 V17 V88 40723.23268130712
L17_88 V17 V88 -1.2605040888206753e-11
C17_88 V17 V88 -2.8446634584210984e-21

R17_89 V17 V89 -51599.6993976312
L17_89 V17 V89 5.472638219272518e-12
C17_89 V17 V89 -2.04320188964012e-20

R17_90 V17 V90 -459941.0966354601
L17_90 V17 V90 9.9772456144137e-12
C17_90 V17 V90 -5.392668346908686e-21

R17_91 V17 V91 145041.29544053116
L17_91 V17 V91 4.178301073869706e-12
C17_91 V17 V91 2.6925640863693047e-21

R17_92 V17 V92 -4619869.743190538
L17_92 V17 V92 6.423354758840595e-12
C17_92 V17 V92 -2.8785980982706595e-21

R17_93 V17 V93 7001.342638087944
L17_93 V17 V93 -2.0716326563753718e-11
C17_93 V17 V93 -8.87499353631643e-21

R17_94 V17 V94 15972.37066558798
L17_94 V17 V94 -7.82939514647511e-12
C17_94 V17 V94 4.591153756375535e-21

R17_95 V17 V95 53723.575874808026
L17_95 V17 V95 9.157892074243696e-12
C17_95 V17 V95 -2.19837524239187e-21

R17_96 V17 V96 -79205.200577682
L17_96 V17 V96 1.5164365813828355e-11
C17_96 V17 V96 -2.652042673126333e-21

R17_97 V17 V97 -728000.7317091181
L17_97 V17 V97 1.8725751756841473e-11
C17_97 V17 V97 -2.4201069691441438e-21

R17_98 V17 V98 -32168.124163636683
L17_98 V17 V98 3.6085950265580554e-12
C17_98 V17 V98 -4.197195732815723e-21

R17_99 V17 V99 40629.437800363085
L17_99 V17 V99 -1.9488782860902634e-11
C17_99 V17 V99 8.275643703012793e-22

R17_100 V17 V100 -102405.28738677554
L17_100 V17 V100 -2.0427159504533754e-11
C17_100 V17 V100 -2.203155285644279e-22

R17_101 V17 V101 31552.297076878494
L17_101 V17 V101 3.660592036440114e-12
C17_101 V17 V101 -1.5341086767943756e-20

R17_102 V17 V102 55414.789815639146
L17_102 V17 V102 2.915596857584907e-12
C17_102 V17 V102 -1.1132716807087845e-20

R17_103 V17 V103 235745.994599861
L17_103 V17 V103 -1.629821526931794e-11
C17_103 V17 V103 -1.1268561113734439e-21

R17_104 V17 V104 93425.41456914377
L17_104 V17 V104 -2.7331429389519633e-11
C17_104 V17 V104 -6.4414360525301475e-21

R17_105 V17 V105 -38524.768048055426
L17_105 V17 V105 -4.1378460689858415e-12
C17_105 V17 V105 -5.146698210232102e-22

R17_106 V17 V106 74970.48055829741
L17_106 V17 V106 3.2414647454765625e-12
C17_106 V17 V106 -4.860878272989249e-22

R17_107 V17 V107 -118369.77202063658
L17_107 V17 V107 4.62164469624042e-12
C17_107 V17 V107 2.5729375611324414e-21

R17_108 V17 V108 -18555.278901843885
L17_108 V17 V108 -3.735870403029681e-12
C17_108 V17 V108 9.67877656121464e-21

R17_109 V17 V109 -30673.881108582333
L17_109 V17 V109 -1.464658415690472e-11
C17_109 V17 V109 1.837128148245312e-21

R17_110 V17 V110 -549040.909371656
L17_110 V17 V110 -3.261674116389218e-12
C17_110 V17 V110 4.175258927477727e-21

R17_111 V17 V111 -14359.333786709929
L17_111 V17 V111 -9.338474776708877e-12
C17_111 V17 V111 -2.4499848953089846e-21

R17_112 V17 V112 -9553.396451499773
L17_112 V17 V112 2.5538075398364756e-12
C17_112 V17 V112 -1.0334739256861695e-20

R17_113 V17 V113 -16335.523730270032
L17_113 V17 V113 6.173107111685914e-12
C17_113 V17 V113 -4.159442642291841e-21

R17_114 V17 V114 85376.92911518893
L17_114 V17 V114 4.89067068665724e-12
C17_114 V17 V114 -2.015190325832392e-21

R17_115 V17 V115 37847.76456168166
L17_115 V17 V115 1.132761551498856e-11
C17_115 V17 V115 -1.459894515284696e-21

R17_116 V17 V116 151199.28466378883
L17_116 V17 V116 -4.992488671340801e-12
C17_116 V17 V116 3.786995549757052e-21

R17_117 V17 V117 23864.024163039787
L17_117 V17 V117 -7.303482414354935e-12
C17_117 V17 V117 8.41876404153506e-21

R17_118 V17 V118 -167745.14463845504
L17_118 V17 V118 -4.771099322094919e-12
C17_118 V17 V118 -3.308062811999955e-21

R17_119 V17 V119 -11400.492131384626
L17_119 V17 V119 -5.553237103512201e-12
C17_119 V17 V119 1.2071404922230343e-21

R17_120 V17 V120 8286.805914958984
L17_120 V17 V120 -1.5480702331807e-11
C17_120 V17 V120 1.883834875229466e-21

R17_121 V17 V121 -5551.493244529748
L17_121 V17 V121 5.019987879148139e-12
C17_121 V17 V121 8.198368954481304e-22

R17_122 V17 V122 -5173.976527340854
L17_122 V17 V122 4.081999018374428e-12
C17_122 V17 V122 -3.1010408045946353e-21

R17_123 V17 V123 -108918.94697302554
L17_123 V17 V123 2.8450179419111222e-11
C17_123 V17 V123 8.198698875353447e-22

R17_124 V17 V124 -81714.08723630967
L17_124 V17 V124 -9.112876868217928e-11
C17_124 V17 V124 1.915438279117869e-21

R17_125 V17 V125 4336.006099282172
L17_125 V17 V125 -4.038560815882683e-12
C17_125 V17 V125 -3.080756898235883e-21

R17_126 V17 V126 10630.938258422853
L17_126 V17 V126 -6.041011131682124e-12
C17_126 V17 V126 -6.928882996486891e-22

R17_127 V17 V127 103338.63224537513
L17_127 V17 V127 8.648430313526296e-12
C17_127 V17 V127 3.235845136895373e-21

R17_128 V17 V128 56293.64134139015
L17_128 V17 V128 4.2884324361313435e-11
C17_128 V17 V128 2.4599915972450923e-21

R17_129 V17 V129 52580.700876396135
L17_129 V17 V129 1.924252719812048e-11
C17_129 V17 V129 8.365083736133232e-21

R17_130 V17 V130 99197.1700213972
L17_130 V17 V130 -1.0302865653503893e-11
C17_130 V17 V130 3.550046037828619e-21

R17_131 V17 V131 25626.40267202736
L17_131 V17 V131 -1.388678875561101e-10
C17_131 V17 V131 -1.7378798940356033e-21

R17_132 V17 V132 79770.34203118825
L17_132 V17 V132 -3.5879890770183284e-11
C17_132 V17 V132 3.1649052181400254e-21

R17_133 V17 V133 28252.818959205248
L17_133 V17 V133 2.310511854855296e-11
C17_133 V17 V133 1.0843367422615423e-21

R17_134 V17 V134 246892.56766115493
L17_134 V17 V134 -1.1277966573184972e-11
C17_134 V17 V134 -2.977066733685378e-21

R17_135 V17 V135 -47583.02528638032
L17_135 V17 V135 1.7570533157015512e-11
C17_135 V17 V135 -8.738321161190957e-22

R17_136 V17 V136 49587.132378216396
L17_136 V17 V136 -4.715147161232758e-11
C17_136 V17 V136 -2.6195222584450446e-21

R17_137 V17 V137 6769.736688499277
L17_137 V17 V137 -7.587948148445451e-12
C17_137 V17 V137 2.6189035444357324e-21

R17_138 V17 V138 11314.304790959606
L17_138 V17 V138 -6.0047210964384245e-12
C17_138 V17 V138 5.2126633720623585e-21

R17_139 V17 V139 34468.43604096414
L17_139 V17 V139 6.201580614260915e-12
C17_139 V17 V139 1.3414007535535932e-21

R17_140 V17 V140 140117.76544351384
L17_140 V17 V140 -7.443807290826523e-12
C17_140 V17 V140 8.105309954039674e-22

R17_141 V17 V141 17402.127272870643
L17_141 V17 V141 -1.664149090327652e-11
C17_141 V17 V141 3.2470102487647626e-21

R17_142 V17 V142 -32320.674381277935
L17_142 V17 V142 -1.0182063651228098e-11
C17_142 V17 V142 3.1839991299552223e-21

R17_143 V17 V143 -39470.64756059163
L17_143 V17 V143 -6.251185217486423e-11
C17_143 V17 V143 -1.5447602109079024e-21

R17_144 V17 V144 -14652.259490643703
L17_144 V17 V144 1.5020542214623018e-11
C17_144 V17 V144 -3.745665298283605e-21

R18_18 V18 0 3403.334502992464
L18_18 V18 0 -2.51873838756897e-11
C18_18 V18 0 3.873699819702937e-20

R18_19 V18 V19 -457510.3345824112
L18_19 V18 V19 -2.9333035364180727e-10
C18_19 V18 V19 -1.6435671369130343e-22

R18_20 V18 V20 645509.1078697874
L18_20 V18 V20 -1.1018539255837913e-10
C18_20 V18 V20 -5.797833223090144e-22

R18_21 V18 V21 -323650.6480801855
L18_21 V18 V21 -4.65761636812535e-11
C18_21 V18 V21 -1.4660239511336588e-21

R18_22 V18 V22 492199.2364371336
L18_22 V18 V22 -1.1744712729332742e-11
C18_22 V18 V22 -6.744819228705454e-22

R18_23 V18 V23 2406720.481617666
L18_23 V18 V23 2.8170445276647253e-11
C18_23 V18 V23 -1.0184474015139345e-23

R18_24 V18 V24 54844752.78711068
L18_24 V18 V24 1.8812913179071922e-11
C18_24 V18 V24 1.4715462902482758e-22

R18_25 V18 V25 256081.66163249925
L18_25 V18 V25 -3.481343438339489e-10
C18_25 V18 V25 -6.433799732862658e-22

R18_26 V18 V26 -216675.73521380746
L18_26 V18 V26 -2.003240790830509e-11
C18_26 V18 V26 2.33912439383604e-21

R18_27 V18 V27 2953838.191558858
L18_27 V18 V27 -1.0820092208304985e-10
C18_27 V18 V27 1.407675130479663e-21

R18_28 V18 V28 2567188.4428402525
L18_28 V18 V28 5.038489798887628e-11
C18_28 V18 V28 -1.3218009264634036e-22

R18_29 V18 V29 -960892.6066002077
L18_29 V18 V29 -4.5880386856413354e-11
C18_29 V18 V29 5.15039202615942e-21

R18_30 V18 V30 116427.37564713367
L18_30 V18 V30 -1.891227435121066e-11
C18_30 V18 V30 4.17052830541844e-22

R18_31 V18 V31 483265.8749787429
L18_31 V18 V31 4.648368310198734e-11
C18_31 V18 V31 1.601876962081201e-21

R18_32 V18 V32 -423873.91715304425
L18_32 V18 V32 3.273265521039467e-11
C18_32 V18 V32 8.275471556548732e-22

R18_33 V18 V33 418887.60931569786
L18_33 V18 V33 1.9570924132017146e-10
C18_33 V18 V33 -3.7643113906566806e-21

R18_34 V18 V34 -159154.6250579401
L18_34 V18 V34 4.880274289946583e-10
C18_34 V18 V34 2.8193643006449373e-21

R18_35 V18 V35 -633693.7510650881
L18_35 V18 V35 -2.3268677543301076e-10
C18_35 V18 V35 -2.6640160185786683e-21

R18_36 V18 V36 114768.57042813639
L18_36 V18 V36 -1.1253246049266325e-10
C18_36 V18 V36 5.229965601701731e-23

R18_37 V18 V37 87809.36701135094
L18_37 V18 V37 -3.4284732618477455e-10
C18_37 V18 V37 1.2342756645137562e-20

R18_38 V18 V38 -112290.86456176972
L18_38 V18 V38 -2.5706973138614453e-11
C18_38 V18 V38 -4.888827541623566e-21

R18_39 V18 V39 -314819.36648965644
L18_39 V18 V39 -3.137834693537234e-10
C18_39 V18 V39 9.906310920920485e-21

R18_40 V18 V40 -143476.6543604893
L18_40 V18 V40 5.213995702485534e-11
C18_40 V18 V40 3.9190132230101874e-22

R18_41 V18 V41 -254301.3476784938
L18_41 V18 V41 2.993189825751071e-11
C18_41 V18 V41 -3.544948582522892e-20

R18_42 V18 V42 -43440.4452014271
L18_42 V18 V42 7.585284471064238e-12
C18_42 V18 V42 -1.1466325146326354e-20

R18_43 V18 V43 52429.41937938214
L18_43 V18 V43 -1.1227963627855495e-10
C18_43 V18 V43 -3.5000879166082215e-20

R18_44 V18 V44 46438.392700568395
L18_44 V18 V44 -3.792538470112751e-11
C18_44 V18 V44 -9.217185791490322e-21

R18_45 V18 V45 44821.06228585728
L18_45 V18 V45 8.49276341636674e-11
C18_45 V18 V45 2.4005265394142968e-20

R18_46 V18 V46 -57815.05193213263
L18_46 V18 V46 -1.8119397428577852e-11
C18_46 V18 V46 4.152069905601865e-21

R18_47 V18 V47 17477.927776322245
L18_47 V18 V47 -4.257520519931075e-11
C18_47 V18 V47 2.5863984401817156e-20

R18_48 V18 V48 23657.66143949375
L18_48 V18 V48 -5.161085642049686e-11
C18_48 V18 V48 9.812458441497993e-21

R18_49 V18 V49 170156.6911059131
L18_49 V18 V49 6.931189070547966e-11
C18_49 V18 V49 -2.8117821496410028e-21

R18_50 V18 V50 -41853.155980226315
L18_50 V18 V50 4.2260002422019934e-10
C18_50 V18 V50 -6.462290664219902e-21

R18_51 V18 V51 363684.6502419504
L18_51 V18 V51 -6.42784013054755e-10
C18_51 V18 V51 -3.923083772930145e-21

R18_52 V18 V52 -38235.98771844772
L18_52 V18 V52 3.2647662029810206e-11
C18_52 V18 V52 -1.546672422195872e-20

R18_53 V18 V53 70177.3248012793
L18_53 V18 V53 -8.598250829079037e-11
C18_53 V18 V53 -1.3343673540978389e-21

R18_54 V18 V54 198743.4999349416
L18_54 V18 V54 9.608110496106833e-11
C18_54 V18 V54 7.89590930245029e-21

R18_55 V18 V55 -160707.294411392
L18_55 V18 V55 8.48982508032904e-11
C18_55 V18 V55 1.0290648561542869e-21

R18_56 V18 V56 -148872.488785315
L18_56 V18 V56 -7.55636095755311e-11
C18_56 V18 V56 6.510417762000778e-21

R18_57 V18 V57 26437.512305027853
L18_57 V18 V57 1.8017829022390894e-11
C18_57 V18 V57 -2.99344047035689e-22

R18_58 V18 V58 -6392.6480183727035
L18_58 V18 V58 9.201307278115108e-12
C18_58 V18 V58 6.978190924939866e-21

R18_59 V18 V59 -34124.65898035364
L18_59 V18 V59 -4.890303697612049e-11
C18_59 V18 V59 4.018341056340263e-21

R18_60 V18 V60 20028.475050931924
L18_60 V18 V60 -2.907215383009164e-11
C18_60 V18 V60 1.6041162731935682e-21

R18_61 V18 V61 -75440.50154994518
L18_61 V18 V61 -5.848610005013466e-11
C18_61 V18 V61 -3.4159234996027934e-21

R18_62 V18 V62 124050.47219413653
L18_62 V18 V62 -2.2171165630161352e-10
C18_62 V18 V62 -1.543117079228705e-20

R18_63 V18 V63 -13494.918509123589
L18_63 V18 V63 4.893239166612429e-11
C18_63 V18 V63 1.1082282812518415e-20

R18_64 V18 V64 -71826.12352603814
L18_64 V18 V64 -6.313237873613095e-11
C18_64 V18 V64 6.422305078824974e-21

R18_65 V18 V65 1068794.7090372394
L18_65 V18 V65 2.6946057161069394e-11
C18_65 V18 V65 -7.097350725809843e-21

R18_66 V18 V66 -43281.778081501165
L18_66 V18 V66 -4.846371275107941e-11
C18_66 V18 V66 3.8358076113043464e-21

R18_67 V18 V67 15608.378341373007
L18_67 V18 V67 2.2572714703426023e-11
C18_67 V18 V67 5.195095980771961e-22

R18_68 V18 V68 40924.33447207422
L18_68 V18 V68 1.0807944835851779e-10
C18_68 V18 V68 -4.1009493457998677e-22

R18_69 V18 V69 30795.482522364444
L18_69 V18 V69 7.120905214464796e-11
C18_69 V18 V69 -2.164628793082001e-21

R18_70 V18 V70 -63912.78749554761
L18_70 V18 V70 -2.5661452378672127e-11
C18_70 V18 V70 1.2502962197441825e-20

R18_71 V18 V71 -18688.723885521184
L18_71 V18 V71 -7.81242106972385e-12
C18_71 V18 V71 3.1830666284558216e-22

R18_72 V18 V72 74685.86494873144
L18_72 V18 V72 3.280045831143699e-11
C18_72 V18 V72 5.679816812659363e-21

R18_73 V18 V73 47351.830369585914
L18_73 V18 V73 2.288020678024244e-11
C18_73 V18 V73 4.764140845269629e-22

R18_74 V18 V74 45059.405263327135
L18_74 V18 V74 -4.1669677479295444e-11
C18_74 V18 V74 3.1923397655376844e-21

R18_75 V18 V75 1134093.9440790378
L18_75 V18 V75 3.882488003004485e-11
C18_75 V18 V75 -6.91378910891507e-21

R18_76 V18 V76 207685.66596799958
L18_76 V18 V76 -1.7126372280126e-11
C18_76 V18 V76 7.417802718768415e-21

R18_77 V18 V77 -557587.4278529387
L18_77 V18 V77 -3.3065025562031246e-11
C18_77 V18 V77 -3.0320424310787367e-22

R18_78 V18 V78 134657.38948727495
L18_78 V18 V78 -6.87513688244535e-11
C18_78 V18 V78 5.002485024517126e-21

R18_79 V18 V79 199347.85303692592
L18_79 V18 V79 -1.4252015215865291e-11
C18_79 V18 V79 1.5599549728904858e-20

R18_80 V18 V80 -151753.10387894683
L18_80 V18 V80 4.1995670371718435e-11
C18_80 V18 V80 -1.5992103062625253e-20

R18_81 V18 V81 1503069.3101057706
L18_81 V18 V81 1.4161485067812706e-11
C18_81 V18 V81 -3.2524524323976854e-22

R18_82 V18 V82 -620566.52677641
L18_82 V18 V82 1.8618217697225797e-10
C18_82 V18 V82 -2.2490874710262598e-20

R18_83 V18 V83 -47703.71410099913
L18_83 V18 V83 -2.7923272448188387e-11
C18_83 V18 V83 -2.227988134183361e-20

R18_84 V18 V84 99072.00970929048
L18_84 V18 V84 -2.142511417273842e-11
C18_84 V18 V84 6.861765372241488e-21

R18_85 V18 V85 141393.22869589957
L18_85 V18 V85 -2.313639065517298e-11
C18_85 V18 V85 1.4196791853539667e-20

R18_86 V18 V86 55538.70011161017
L18_86 V18 V86 3.893059811741358e-11
C18_86 V18 V86 9.156916934608268e-21

R18_87 V18 V87 88674.18215236663
L18_87 V18 V87 -2.6456922306836017e-11
C18_87 V18 V87 1.8794511078587653e-20

R18_88 V18 V88 206783.34906330687
L18_88 V18 V88 5.8200340680963914e-11
C18_88 V18 V88 1.4655926475430685e-21

R18_89 V18 V89 944876.3542041574
L18_89 V18 V89 2.016785664393609e-10
C18_89 V18 V89 -8.796997204664575e-21

R18_90 V18 V90 -39829.01619001411
L18_90 V18 V90 1.1102281364166086e-11
C18_90 V18 V90 -1.4562936873853684e-20

R18_91 V18 V91 -65957.26622404183
L18_91 V18 V91 2.488716443761271e-10
C18_91 V18 V91 -2.155724130907389e-20

R18_92 V18 V92 -203000.37034622277
L18_92 V18 V92 -2.0619695320873642e-11
C18_92 V18 V92 -1.3571031664943838e-20

R18_93 V18 V93 2429727.5007927055
L18_93 V18 V93 -4.91747279371972e-11
C18_93 V18 V93 3.650278500273181e-21

R18_94 V18 V94 36142.76848831739
L18_94 V18 V94 2.3538843121741067e-11
C18_94 V18 V94 4.508028877745521e-21

R18_95 V18 V95 -63533.47878950379
L18_95 V18 V95 -2.05758448987855e-10
C18_95 V18 V95 -1.2284875924552105e-20

R18_96 V18 V96 -147533.14305302838
L18_96 V18 V96 -1.892295553309727e-11
C18_96 V18 V96 -7.167893508019294e-21

R18_97 V18 V97 -68586.90823620302
L18_97 V18 V97 1.0441207357503547e-11
C18_97 V18 V97 -2.6776882141626614e-21

R18_98 V18 V98 -34494.527241848824
L18_98 V18 V98 3.815004644693913e-11
C18_98 V18 V98 -1.4258599355938843e-20

R18_99 V18 V99 27739.077005237297
L18_99 V18 V99 -2.6132428133923227e-11
C18_99 V18 V99 4.621475287485263e-21

R18_100 V18 V100 262291.73098549695
L18_100 V18 V100 3.3151682814983484e-11
C18_100 V18 V100 1.4652983240591672e-21

R18_101 V18 V101 288686.61978293874
L18_101 V18 V101 3.0835657216837537e-10
C18_101 V18 V101 -1.2004496334194123e-20

R18_102 V18 V102 -32808.440312473846
L18_102 V18 V102 5.298637239301825e-12
C18_102 V18 V102 -3.563311912696834e-20

R18_103 V18 V103 147996.85130548087
L18_103 V18 V103 -1.0085311621280246e-11
C18_103 V18 V103 1.7286604614362172e-20

R18_104 V18 V104 99997.1893794589
L18_104 V18 V104 -2.358624757937239e-11
C18_104 V18 V104 2.555769918590008e-21

R18_105 V18 V105 108381.7097105585
L18_105 V18 V105 -2.257633691172357e-11
C18_105 V18 V105 1.860882019030406e-20

R18_106 V18 V106 1711473.3919189204
L18_106 V18 V106 1.9341644528154314e-11
C18_106 V18 V106 -3.612644893253553e-20

R18_107 V18 V107 -312616.9535446907
L18_107 V18 V107 7.208013071489174e-12
C18_107 V18 V107 -3.3168386988931564e-20

R18_108 V18 V108 -58229.08530198276
L18_108 V18 V108 -9.756773094599345e-12
C18_108 V18 V108 2.9688853359492986e-20

R18_109 V18 V109 208660.46371481364
L18_109 V18 V109 -1.0824887675788454e-11
C18_109 V18 V109 1.3238895500333346e-20

R18_110 V18 V110 -24210.0590166143
L18_110 V18 V110 4.6003170840961497e-10
C18_110 V18 V110 2.7545751022368715e-20

R18_111 V18 V111 22431.824747798673
L18_111 V18 V111 -1.4480243066332679e-11
C18_111 V18 V111 1.764094143046713e-20

R18_112 V18 V112 -20340.94517349854
L18_112 V18 V112 8.459699042412703e-12
C18_112 V18 V112 -2.4945667470673253e-20

R18_113 V18 V113 -28208.452984365147
L18_113 V18 V113 1.424663879500922e-11
C18_113 V18 V113 -9.854717843251005e-21

R18_114 V18 V114 -46178.278799248576
L18_114 V18 V114 2.907869171113161e-11
C18_114 V18 V114 -1.6730056889254404e-20

R18_115 V18 V115 -32652.248869452236
L18_115 V18 V115 1.6576666967704275e-11
C18_115 V18 V115 -1.8037293130225638e-20

R18_116 V18 V116 44943.18756717406
L18_116 V18 V116 -1.8822067833050148e-11
C18_116 V18 V116 1.651509614624851e-20

R18_117 V18 V117 -43058.126467055066
L18_117 V18 V117 -2.216414268856012e-11
C18_117 V18 V117 1.2512283798409479e-20

R18_118 V18 V118 48097.764801105426
L18_118 V18 V118 -2.2376320448566194e-11
C18_118 V18 V118 1.6289598418893568e-20

R18_119 V18 V119 28050.061875102154
L18_119 V18 V119 -4.69476339838101e-11
C18_119 V18 V119 2.0354021436209193e-20

R18_120 V18 V120 -7447.726899857528
L18_120 V18 V120 1.4257832987636431e-11
C18_120 V18 V120 6.5690668679730704e-21

R18_121 V18 V121 -72186.91964249017
L18_121 V18 V121 3.0065769783524785e-11
C18_121 V18 V121 -3.154673243639919e-21

R18_122 V18 V122 -5246.285520475178
L18_122 V18 V122 7.336739545648455e-12
C18_122 V18 V122 1.927544447294677e-21

R18_123 V18 V123 -26746.77148578486
L18_123 V18 V123 2.771594053057235e-11
C18_123 V18 V123 2.6749808229079426e-21

R18_124 V18 V124 78766.01105548283
L18_124 V18 V124 3.1427464278367776e-10
C18_124 V18 V124 4.781759895918946e-21

R18_125 V18 V125 -30228.825177222658
L18_125 V18 V125 -1.18579230057715e-10
C18_125 V18 V125 4.967860690783527e-21

R18_126 V18 V126 4114.703659144441
L18_126 V18 V126 -6.503386714215655e-12
C18_126 V18 V126 -2.0203256205740847e-21

R18_127 V18 V127 -5419.80064073227
L18_127 V18 V127 8.348176134485146e-12
C18_127 V18 V127 -3.2484600372799803e-22

R18_128 V18 V128 -58114.5850038893
L18_128 V18 V128 7.163484182397213e-10
C18_128 V18 V128 -1.0703883170886265e-21

R18_129 V18 V129 -14840.191640714176
L18_129 V18 V129 2.1026353757329742e-11
C18_129 V18 V129 -1.073451446368638e-21

R18_130 V18 V130 20089.89671718057
L18_130 V18 V130 -1.0491493289391796e-11
C18_130 V18 V130 7.382837818862695e-21

R18_131 V18 V131 16820.210254592446
L18_131 V18 V131 -4.828690596777809e-11
C18_131 V18 V131 -6.6738082649295044e-21

R18_132 V18 V132 21149.81392993419
L18_132 V18 V132 -4.056495128208435e-11
C18_132 V18 V132 -1.356155062091762e-21

R18_133 V18 V133 126457.14062785114
L18_133 V18 V133 -4.477062771487743e-10
C18_133 V18 V133 -1.0349502071889396e-20

R18_134 V18 V134 27760.88880281193
L18_134 V18 V134 -4.2343824651316104e-11
C18_134 V18 V134 -6.607553564898747e-23

R18_135 V18 V135 -8007.626969033082
L18_135 V18 V135 1.2646272346740357e-11
C18_135 V18 V135 4.259534115503364e-21

R18_136 V18 V136 -241862.84665998194
L18_136 V18 V136 2.2315236988201327e-10
C18_136 V18 V136 3.31449868694521e-21

R18_137 V18 V137 -180583.21180335002
L18_137 V18 V137 -4.793675487318482e-11
C18_137 V18 V137 6.139264141160506e-21

R18_138 V18 V138 4797.877650188076
L18_138 V18 V138 -6.567566426341995e-12
C18_138 V18 V138 8.218628135991729e-22

R18_139 V18 V139 -4128.43504845679
L18_139 V18 V139 6.156077065429159e-12
C18_139 V18 V139 -3.818395980642625e-21

R18_140 V18 V140 17112.11261705591
L18_140 V18 V140 -1.5593504854276466e-11
C18_140 V18 V140 4.0989934591985944e-21

R18_141 V18 V141 21320.49429320659
L18_141 V18 V141 -3.448521614452223e-11
C18_141 V18 V141 2.3078849767736723e-21

R18_142 V18 V142 16698.7008528272
L18_142 V18 V142 -1.2490217184249345e-11
C18_142 V18 V142 3.0874756171883356e-21

R18_143 V18 V143 13003.808419603898
L18_143 V18 V143 -2.1726058140249036e-11
C18_143 V18 V143 1.090119928794307e-21

R18_144 V18 V144 -34693.72966795582
L18_144 V18 V144 5.326821404697745e-11
C18_144 V18 V144 -4.9796806168598756e-21

R19_19 V19 0 480.68078035716917
L19_19 V19 0 -9.459080825921432e-13
C19_19 V19 0 -1.3264605127744094e-20

R19_20 V19 V20 707085.0123567327
L19_20 V19 V20 3.067855146029274e-10
C19_20 V19 V20 -9.877913380950378e-22

R19_21 V19 V21 45987.45971181707
L19_21 V19 V21 -1.207153722032175e-11
C19_21 V19 V21 -1.0657219282982817e-20

R19_22 V19 V22 -364478.5666078551
L19_22 V19 V22 2.2043174675745455e-11
C19_22 V19 V22 -4.040014482218333e-22

R19_23 V19 V23 70732.6714229624
L19_23 V19 V23 1.7231600367026417e-11
C19_23 V19 V23 -4.9339182288698586e-21

R19_24 V19 V24 -1168595.6146742427
L19_24 V19 V24 -5.923092090206711e-11
C19_24 V19 V24 3.089077446828709e-22

R19_25 V19 V25 53931.64247655753
L19_25 V19 V25 -2.1845862622931334e-11
C19_25 V19 V25 1.6776618377945094e-20

R19_26 V19 V26 140619.97079079985
L19_26 V19 V26 2.684176957047933e-11
C19_26 V19 V26 -1.4060563208705852e-21

R19_27 V19 V27 -226728.70410170325
L19_27 V19 V27 -1.409501585231167e-10
C19_27 V19 V27 2.21657092852583e-20

R19_28 V19 V28 109190.77180102663
L19_28 V19 V28 -1.0129899072286666e-10
C19_28 V19 V28 2.300498269850256e-21

R19_29 V19 V29 -21951.546803587116
L19_29 V19 V29 -1.513845087854564e-11
C19_29 V19 V29 -6.534921922729673e-21

R19_30 V19 V30 -81077.48140029675
L19_30 V19 V30 7.619145831582163e-11
C19_30 V19 V30 -7.195620583775543e-21

R19_31 V19 V31 -50259.18539084217
L19_31 V19 V31 9.849138345538644e-12
C19_31 V19 V31 -2.7438078108231223e-21

R19_32 V19 V32 -253070.54908892087
L19_32 V19 V32 -1.0630406374420832e-10
C19_32 V19 V32 -6.304089141780557e-21

R19_33 V19 V33 -10087.441287592745
L19_33 V19 V33 1.3729736002655896e-11
C19_33 V19 V33 -1.2416991036839096e-20

R19_34 V19 V34 15576.720553662302
L19_34 V19 V34 -1.7125092009309286e-10
C19_34 V19 V34 1.0833973956846998e-20

R19_35 V19 V35 -6798.98156582134
L19_35 V19 V35 -1.3942057924680494e-11
C19_35 V19 V35 1.1874612702651318e-21

R19_36 V19 V36 30483.663451766974
L19_36 V19 V36 -4.19193709011606e-10
C19_36 V19 V36 4.0039421263799054e-21

R19_37 V19 V37 9157.881029741939
L19_37 V19 V37 -1.0853938046820045e-11
C19_37 V19 V37 -9.55029185106766e-21

R19_38 V19 V38 -24544.648304332502
L19_38 V19 V38 -5.3902915207189517e-11
C19_38 V19 V38 1.1166983712892513e-20

R19_39 V19 V39 -203112.75396719787
L19_39 V19 V39 -6.132596160191906e-11
C19_39 V19 V39 -3.0960969712973007e-20

R19_40 V19 V40 -23294.910821749978
L19_40 V19 V40 -5.917137256142422e-11
C19_40 V19 V40 -8.689890918642912e-22

R19_41 V19 V41 -6365.14221052981
L19_41 V19 V41 2.4847394605971347e-12
C19_41 V19 V41 1.963445739660076e-20

R19_42 V19 V42 -73565.34628701863
L19_42 V19 V42 4.1748921173972515e-12
C19_42 V19 V42 1.1480307689917496e-20

R19_43 V19 V43 -24928.593643162534
L19_43 V19 V43 1.0456629747103558e-11
C19_43 V19 V43 3.9966307457826585e-20

R19_44 V19 V44 15278.151164132581
L19_44 V19 V44 1.174753411529128e-11
C19_44 V19 V44 -3.958199187433334e-20

R19_45 V19 V45 -407829.6448372287
L19_45 V19 V45 1.1600049821217811e-10
C19_45 V19 V45 -1.0386231980012538e-19

R19_46 V19 V46 -6235.612710130886
L19_46 V19 V46 -8.197756302012702e-12
C19_46 V19 V46 7.176075588488947e-20

R19_47 V19 V47 -3487.363337173427
L19_47 V19 V47 -1.9161356422323468e-11
C19_47 V19 V47 2.6655962813982135e-20

R19_48 V19 V48 8012.6539344853845
L19_48 V19 V48 9.948084125327139e-10
C19_48 V19 V48 1.072139804297398e-20

R19_49 V19 V49 3184.6853974753635
L19_49 V19 V49 2.676881182985063e-11
C19_49 V19 V49 3.0263347325709614e-20

R19_50 V19 V50 -3126.563952752812
L19_50 V19 V50 -8.379608355679448e-11
C19_50 V19 V50 -2.0228187875093722e-20

R19_51 V19 V51 16089.961143231549
L19_51 V19 V51 -8.635069175289303e-11
C19_51 V19 V51 -9.798334431063831e-21

R19_52 V19 V52 280874.82902270433
L19_52 V19 V52 1.94051233618785e-11
C19_52 V19 V52 1.6378946307242195e-20

R19_53 V19 V53 -18177.1589685564
L19_53 V19 V53 4.2942135974687434e-11
C19_53 V19 V53 1.0708440186080516e-20

R19_54 V19 V54 -10096.071910300789
L19_54 V19 V54 2.410482974161714e-11
C19_54 V19 V54 1.3987322939208012e-20

R19_55 V19 V55 23852.639007398073
L19_55 V19 V55 9.768344431531543e-12
C19_55 V19 V55 5.838747752542147e-20

R19_56 V19 V56 -14641.339867209115
L19_56 V19 V56 1.2962167366042193e-11
C19_56 V19 V56 2.254402827629119e-20

R19_57 V19 V57 -1284.4018897352541
L19_57 V19 V57 3.132464370852979e-12
C19_57 V19 V57 -8.777482928313509e-22

R19_58 V19 V58 -18963.631409972615
L19_58 V19 V58 1.7273923664926604e-11
C19_58 V19 V58 2.3452576287090125e-21

R19_59 V19 V59 -2084.319641414529
L19_59 V19 V59 -7.485553747614335e-12
C19_59 V19 V59 -1.7584964431077498e-20

R19_60 V19 V60 -7158.351819486716
L19_60 V19 V60 1.547452879730939e-11
C19_60 V19 V60 4.265927101020031e-21

R19_61 V19 V61 3591.352825487666
L19_61 V19 V61 -5.01551494997559e-11
C19_61 V19 V61 4.912777091506595e-22

R19_62 V19 V62 11175.739812476817
L19_62 V19 V62 -1.2225838202042258e-11
C19_62 V19 V62 -5.101840511965932e-21

R19_63 V19 V63 23979.925343707164
L19_63 V19 V63 1.7302008172369108e-11
C19_63 V19 V63 9.823146079341376e-21

R19_64 V19 V64 -16571.971045614624
L19_64 V19 V64 -8.076912906111465e-11
C19_64 V19 V64 -6.997433150505558e-21

R19_65 V19 V65 -3093.196825288313
L19_65 V19 V65 1.6885492936860065e-11
C19_65 V19 V65 -3.057627826400181e-20

R19_66 V19 V66 -5837.362426811419
L19_66 V19 V66 -2.4281340375017424e-11
C19_66 V19 V66 3.099648761747282e-20

R19_67 V19 V67 -10264.363987906556
L19_67 V19 V67 3.501559389209615e-11
C19_67 V19 V67 2.1438459972198278e-20

R19_68 V19 V68 26363.35809913364
L19_68 V19 V68 2.1658689562799952e-11
C19_68 V19 V68 -8.067652946362947e-21

R19_69 V19 V69 5262.446936447761
L19_69 V19 V69 6.307432982816126e-10
C19_69 V19 V69 -2.664145872893678e-20

R19_70 V19 V70 -38315.88141228427
L19_70 V19 V70 2.208366150655385e-11
C19_70 V19 V70 3.233837715660416e-20

R19_71 V19 V71 -240341.7372342151
L19_71 V19 V71 3.016081484310223e-10
C19_71 V19 V71 -1.0979041723063097e-21

R19_72 V19 V72 39801.50730732177
L19_72 V19 V72 1.2557791883495541e-11
C19_72 V19 V72 2.6249710451144973e-20

R19_73 V19 V73 36892.79990546939
L19_73 V19 V73 2.135343391317917e-11
C19_73 V19 V73 2.406146657614154e-21

R19_74 V19 V74 9759.320045279354
L19_74 V19 V74 7.679153415156311e-10
C19_74 V19 V74 -6.622395480839486e-21

R19_75 V19 V75 -91302.04977170868
L19_75 V19 V75 -2.4853377009015388e-11
C19_75 V19 V75 -8.651141797189116e-21

R19_76 V19 V76 -49756.351476050746
L19_76 V19 V76 -6.718244383584523e-11
C19_76 V19 V76 1.977849809191819e-22

R19_77 V19 V77 -365961.6363641308
L19_77 V19 V77 7.535466981851373e-11
C19_77 V19 V77 4.801921565966112e-23

R19_78 V19 V78 75952.3244582155
L19_78 V19 V78 -3.816797841735796e-11
C19_78 V19 V78 2.1529122874416717e-20

R19_79 V19 V79 41826.54152365506
L19_79 V19 V79 3.348371340316758e-11
C19_79 V19 V79 -1.9040901901198947e-21

R19_80 V19 V80 78664.62111308529
L19_80 V19 V80 2.052991963178426e-11
C19_80 V19 V80 -2.5807834055397382e-21

R19_81 V19 V81 -340332.4425904207
L19_81 V19 V81 -1.406431867762012e-11
C19_81 V19 V81 -6.92807103841628e-21

R19_82 V19 V82 -92932.0019182982
L19_82 V19 V82 -1.992313948775052e-11
C19_82 V19 V82 -8.660619428526454e-20

R19_83 V19 V83 -38818.58307873034
L19_83 V19 V83 -2.3603243020496992e-11
C19_83 V19 V83 -5.3169734531261996e-20

R19_84 V19 V84 -71278.88876463094
L19_84 V19 V84 -8.624741651087822e-11
C19_84 V19 V84 -3.753893357872631e-22

R19_85 V19 V85 100385.63206716118
L19_85 V19 V85 -1.9269324616892895e-10
C19_85 V19 V85 1.486579634792932e-20

R19_86 V19 V86 30495.04187538426
L19_86 V19 V86 3.854456763613146e-11
C19_86 V19 V86 4.1294596129559224e-20

R19_87 V19 V87 36508.08622590207
L19_87 V19 V87 -3.1309193946740985e-10
C19_87 V19 V87 4.485133040738911e-20

R19_88 V19 V88 69420.92723754478
L19_88 V19 V88 -2.8166525531721345e-11
C19_88 V19 V88 9.317244094459337e-21

R19_89 V19 V89 -82151.38190392373
L19_89 V19 V89 1.436196861697414e-11
C19_89 V19 V89 -3.1205091869100885e-20

R19_90 V19 V90 453411.1477167767
L19_90 V19 V90 3.410034003949623e-10
C19_90 V19 V90 1.0155420303926399e-20

R19_91 V19 V91 -28714.784228760796
L19_91 V19 V91 -1.0810411671796598e-11
C19_91 V19 V91 -1.0173847477597966e-19

R19_92 V19 V92 792639.8953401931
L19_92 V19 V92 2.914932925620017e-11
C19_92 V19 V92 -2.767401895200193e-20

R19_93 V19 V93 15058.799063959012
L19_93 V19 V93 -1.532965867656647e-10
C19_93 V19 V93 3.1496791704661158e-21

R19_94 V19 V94 26544.22481921096
L19_94 V19 V94 -2.1561182556563627e-11
C19_94 V19 V94 2.68286239264451e-20

R19_95 V19 V95 -117451.47922554644
L19_95 V19 V95 -2.478510494479471e-11
C19_95 V19 V95 -4.556814623442261e-20

R19_96 V19 V96 -53580.806875797505
L19_96 V19 V96 2.2622746295435272e-11
C19_96 V19 V96 3.1755206642730094e-21

R19_97 V19 V97 153235.5033094626
L19_97 V19 V97 2.7030346579441003e-11
C19_97 V19 V97 2.3164877294977005e-20

R19_98 V19 V98 -52481.389097658415
L19_98 V19 V98 1.1887953653424203e-11
C19_98 V19 V98 -2.8358547865952165e-20

R19_99 V19 V99 50439.8258484559
L19_99 V19 V99 4.376313896808637e-10
C19_99 V19 V99 9.093336309794097e-22

R19_100 V19 V100 -408037.4666453675
L19_100 V19 V100 -5.116087420692729e-11
C19_100 V19 V100 6.208335561508952e-21

R19_101 V19 V101 -1191520.9868630222
L19_101 V19 V101 1.0890717638227547e-11
C19_101 V19 V101 -3.56206691119458e-20

R19_102 V19 V102 34091.60893116936
L19_102 V19 V102 5.560776322114022e-11
C19_102 V19 V102 -7.728536894052783e-21

R19_103 V19 V103 160679.66997480328
L19_103 V19 V103 4.790633899846396e-11
C19_103 V19 V103 -2.2521527927734224e-20

R19_104 V19 V104 46555.175487788314
L19_104 V19 V104 1.731179409699574e-11
C19_104 V19 V104 2.4872475650511236e-20

R19_105 V19 V105 -171698.92800347504
L19_105 V19 V105 4.0848659308486293e-10
C19_105 V19 V105 3.6043710898719565e-20

R19_106 V19 V106 -47429.760614039864
L19_106 V19 V106 -1.0842841676100693e-11
C19_106 V19 V106 -7.941181925583711e-20

R19_107 V19 V107 -109580.1428709532
L19_107 V19 V107 -4.516728298099775e-11
C19_107 V19 V107 -3.0087696692727834e-21

R19_108 V19 V108 -38370.00224754991
L19_108 V19 V108 -2.3481971625994096e-11
C19_108 V19 V108 1.0736222472843823e-20

R19_109 V19 V109 -366706.6405355315
L19_109 V19 V109 1.743149060636144e-11
C19_109 V19 V109 1.0670245291255852e-20

R19_110 V19 V110 28627.248302416057
L19_110 V19 V110 5.055900698444273e-11
C19_110 V19 V110 6.60619763546219e-20

R19_111 V19 V111 -50082.91230470095
L19_111 V19 V111 1.6511643067793453e-11
C19_111 V19 V111 9.719586563051986e-21

R19_112 V19 V112 -28881.39419839287
L19_112 V19 V112 1.043654224727046e-11
C19_112 V19 V112 -2.531698818876152e-20

R19_113 V19 V113 -18706.436694115993
L19_113 V19 V113 1.1009524870742577e-10
C19_113 V19 V113 -1.665570786151751e-20

R19_114 V19 V114 241510.75810716907
L19_114 V19 V114 -2.1987519978935537e-10
C19_114 V19 V114 -4.04324559903539e-20

R19_115 V19 V115 40742.45253505308
L19_115 V19 V115 -3.839334860748281e-11
C19_115 V19 V115 -2.9262963411764917e-21

R19_116 V19 V116 -177143.26054314553
L19_116 V19 V116 -1.9646874852815295e-11
C19_116 V19 V116 3.650893575457912e-21

R19_117 V19 V117 47452.554907366895
L19_117 V19 V117 -4.0703027577576266e-11
C19_117 V19 V117 1.2454427279986679e-20

R19_118 V19 V118 56323.09090613917
L19_118 V19 V118 3.518905089745106e-11
C19_118 V19 V118 4.490335723762697e-20

R19_119 V19 V119 -28964.44520570414
L19_119 V19 V119 1.923230461116283e-11
C19_119 V19 V119 4.981869725696464e-20

R19_120 V19 V120 23215.980022841668
L19_120 V19 V120 -1.13732146687768e-11
C19_120 V19 V120 5.572079998611214e-21

R19_121 V19 V121 -14254.237019275422
L19_121 V19 V121 1.251188822427907e-11
C19_121 V19 V121 -7.966059805106005e-21

R19_122 V19 V122 -12701.168832595273
L19_122 V19 V122 1.193560287167759e-11
C19_122 V19 V122 -1.2767346514209432e-21

R19_123 V19 V123 51143.42587054007
L19_123 V19 V123 1.6425951859287994e-11
C19_123 V19 V123 1.0429317056520173e-20

R19_124 V19 V124 23485.767726962404
L19_124 V19 V124 3.230841902277816e-11
C19_124 V19 V124 7.262551911207558e-21

R19_125 V19 V125 10278.469222797901
L19_125 V19 V125 -7.073398679102734e-12
C19_125 V19 V125 6.38493140035843e-21

R19_126 V19 V126 22998.92278380902
L19_126 V19 V126 -1.1043502910982154e-10
C19_126 V19 V126 -2.450603514898766e-21

R19_127 V19 V127 1720167.6250565958
L19_127 V19 V127 -2.7685506014451835e-11
C19_127 V19 V127 -8.808305483118648e-22

R19_128 V19 V128 -40674.593219638846
L19_128 V19 V128 9.507603098603877e-11
C19_128 V19 V128 2.8512092662346843e-22

R19_129 V19 V129 19569.805390260586
L19_129 V19 V129 7.012262861967983e-11
C19_129 V19 V129 -5.338932010674096e-22

R19_130 V19 V130 -38516.73921015262
L19_130 V19 V130 -4.17884620954357e-11
C19_130 V19 V130 6.918369257906657e-21

R19_131 V19 V131 -72278.80821681049
L19_131 V19 V131 -2.7130937799023555e-11
C19_131 V19 V131 4.587975826826443e-21

R19_132 V19 V132 469960.5111770031
L19_132 V19 V132 -3.4449297122892914e-11
C19_132 V19 V132 -1.2970933196319258e-20

R19_133 V19 V133 -264285.33705158526
L19_133 V19 V133 -1.0140192445676793e-11
C19_133 V19 V133 -4.0257061938695013e-20

R19_134 V19 V134 102505.96938466515
L19_134 V19 V134 -2.7134914332852177e-11
C19_134 V19 V134 6.729796152587734e-21

R19_135 V19 V135 -55098.85302087587
L19_135 V19 V135 -6.474882128119279e-11
C19_135 V19 V135 -9.95396565576736e-22

R19_136 V19 V136 -85084.30748096287
L19_136 V19 V136 -2.9579238634933945e-10
C19_136 V19 V136 8.447803757223648e-21

R19_137 V19 V137 12206.599408150301
L19_137 V19 V137 -2.7989515785673584e-11
C19_137 V19 V137 2.0451433096870453e-20

R19_138 V19 V138 53283.4163642438
L19_138 V19 V138 -2.3169468376804023e-11
C19_138 V19 V138 -4.972163544420009e-21

R19_139 V19 V139 -391987.2894583922
L19_139 V19 V139 -2.4886697088090622e-11
C19_139 V19 V139 -4.800256990161306e-21

R19_140 V19 V140 -89907.97989531016
L19_140 V19 V140 -5.443400218154025e-11
C19_140 V19 V140 9.04313109941849e-21

R19_141 V19 V141 16115.566980630134
L19_141 V19 V141 -1.973601489596738e-10
C19_141 V19 V141 1.3082909786418335e-21

R19_142 V19 V142 -16891.967122060407
L19_142 V19 V142 -4.011629251695981e-11
C19_142 V19 V142 4.125246143029683e-22

R19_143 V19 V143 -48041.70771524032
L19_143 V19 V143 1.1525220611175897e-10
C19_143 V19 V143 -4.874076075558719e-21

R19_144 V19 V144 -29422.573510359816
L19_144 V19 V144 1.1460515107435593e-10
C19_144 V19 V144 -8.290882771974408e-21

R20_20 V20 0 4000.580903746037
L20_20 V20 0 -3.6143690464386485e-12
C20_20 V20 0 -1.31017667713119e-19

R20_21 V20 V21 -171249.7216070332
L20_21 V20 V21 5.312119539803912e-11
C20_21 V20 V21 2.224457530288229e-21

R20_22 V20 V22 -543674.8466499144
L20_22 V20 V22 6.984491070832958e-11
C20_22 V20 V22 -1.2968397312893259e-21

R20_23 V20 V23 -176934.58607461923
L20_23 V20 V23 6.539764849580767e-11
C20_23 V20 V23 -8.734383426182691e-22

R20_24 V20 V24 -2006252.6359208885
L20_24 V20 V24 1.3875237878863654e-11
C20_24 V20 V24 -2.2073242258364557e-21

R20_25 V20 V25 127077.77777433918
L20_25 V20 V25 -2.447919357548469e-10
C20_25 V20 V25 -4.804835206545243e-21

R20_26 V20 V26 325127.1896360949
L20_26 V20 V26 6.020471075707044e-10
C20_26 V20 V26 -3.2924072865417496e-21

R20_27 V20 V27 84034.96190773908
L20_27 V20 V27 -3.3168867720526756e-10
C20_27 V20 V27 -3.988954353229423e-21

R20_28 V20 V28 89360.46893466571
L20_28 V20 V28 4.5344886555527525e-11
C20_28 V20 V28 7.095022912514335e-21

R20_29 V20 V29 1015400.892876543
L20_29 V20 V29 7.010061570118363e-10
C20_29 V20 V29 9.365541620360802e-22

R20_30 V20 V30 -75785.62256716909
L20_30 V20 V30 1.4968694857327134e-10
C20_30 V20 V30 1.9905455101227222e-21

R20_31 V20 V31 -685470.0505244134
L20_31 V20 V31 -1.131522199852383e-10
C20_31 V20 V31 8.452934131882922e-22

R20_32 V20 V32 -1060674.8257749116
L20_32 V20 V32 1.1808120368580822e-11
C20_32 V20 V32 -9.682680358957968e-21

R20_33 V20 V33 36036.01455874599
L20_33 V20 V33 -9.973020410892675e-11
C20_33 V20 V33 2.5174912888496887e-21

R20_34 V20 V34 -193896.923908783
L20_34 V20 V34 -6.958717654101023e-10
C20_34 V20 V34 1.0144029321723532e-21

R20_35 V20 V35 26903.056678609635
L20_35 V20 V35 -2.74606830404498e-10
C20_35 V20 V35 2.71963039976389e-21

R20_36 V20 V36 -12401.753098322612
L20_36 V20 V36 -3.03317949814235e-11
C20_36 V20 V36 1.1100009396312023e-20

R20_37 V20 V37 -85976.4600913732
L20_37 V20 V37 6.571404476110194e-11
C20_37 V20 V37 6.6377216641082126e-21

R20_38 V20 V38 68076.32554430855
L20_38 V20 V38 -8.938389015878535e-11
C20_38 V20 V38 9.625069113798485e-21

R20_39 V20 V39 -107106.11090199386
L20_39 V20 V39 7.955159512071197e-11
C20_39 V20 V39 1.0172462795421567e-20

R20_40 V20 V40 -43382.85155220245
L20_40 V20 V40 1.0541813557109356e-11
C20_40 V20 V40 -6.734558165946851e-20

R20_41 V20 V41 24612.55604854765
L20_41 V20 V41 -1.9344388739762073e-11
C20_41 V20 V41 -4.808314463349642e-21

R20_42 V20 V42 25487.76319503409
L20_42 V20 V42 -1.9425985998702038e-11
C20_42 V20 V42 -2.8191110248894544e-20

R20_43 V20 V43 100138.94187819569
L20_43 V20 V43 -5.650244219827019e-11
C20_43 V20 V43 -3.3130218603639314e-21

R20_44 V20 V44 -13791.854020792585
L20_44 V20 V44 -8.98018582074175e-12
C20_44 V20 V44 1.1369464970226274e-19

R20_45 V20 V45 21827.69751130608
L20_45 V20 V45 1.457298579558856e-11
C20_45 V20 V45 -1.40313329992645e-20

R20_46 V20 V46 12448.410518356915
L20_46 V20 V46 -2.254593351128029e-11
C20_46 V20 V46 2.8596331878058284e-20

R20_47 V20 V47 -38106.99212272289
L20_47 V20 V47 -1.459947495409267e-09
C20_47 V20 V47 -6.7737194426185066e-21

R20_48 V20 V48 -5551.124876502002
L20_48 V20 V48 -2.561696699207954e-11
C20_48 V20 V48 -1.923221475997178e-20

R20_49 V20 V49 -18827.38787873168
L20_49 V20 V49 6.398161534813689e-11
C20_49 V20 V49 -2.604060679575106e-21

R20_50 V20 V50 18816.19825691145
L20_50 V20 V50 -3.610572978404025e-11
C20_50 V20 V50 3.5229720696656e-21

R20_51 V20 V51 -28289.64568851058
L20_51 V20 V51 9.252632051439304e-11
C20_51 V20 V51 5.670909942883187e-21

R20_52 V20 V52 22415.196313613982
L20_52 V20 V52 -7.871833595988559e-11
C20_52 V20 V52 1.1786012140279191e-20

R20_53 V20 V53 -15355.434445702345
L20_53 V20 V53 -1.6497981369592592e-10
C20_53 V20 V53 -3.048888387183366e-20

R20_54 V20 V54 -208591.90916105133
L20_54 V20 V54 3.315428612169054e-10
C20_54 V20 V54 -1.2612338071253294e-20

R20_55 V20 V55 61514.15466376213
L20_55 V20 V55 -3.499308559493136e-11
C20_55 V20 V55 -5.147975897151137e-21

R20_56 V20 V56 7870.751750897328
L20_56 V20 V56 1.63835634066373e-11
C20_56 V20 V56 6.479784954173648e-20

R20_57 V20 V57 4579.219762118841
L20_57 V20 V57 -2.2127992690875316e-11
C20_57 V20 V57 2.205454449943891e-21

R20_58 V20 V58 7018.261993707576
L20_58 V20 V58 3.630546166618e-11
C20_58 V20 V58 -1.3557057774268934e-21

R20_59 V20 V59 17085.489340669916
L20_59 V20 V59 5.886219354242879e-11
C20_59 V20 V59 2.209475187229452e-21

R20_60 V20 V60 -2276.921631139592
L20_60 V20 V60 -1.3170383095639596e-11
C20_60 V20 V60 -6.039526306879811e-21

R20_61 V20 V61 -17747.004016054492
L20_61 V20 V61 2.8659728226772605e-11
C20_61 V20 V61 -1.3334042174141509e-21

R20_62 V20 V62 -7555.7347503379815
L20_62 V20 V62 -1.1677755305973582e-10
C20_62 V20 V62 -4.18569500785995e-21

R20_63 V20 V63 170672.44354319965
L20_63 V20 V63 -7.648668866418213e-11
C20_63 V20 V63 2.754531280147052e-21

R20_64 V20 V64 19178.757626382663
L20_64 V20 V64 1.8581272353451197e-10
C20_64 V20 V64 4.080202540169513e-20

R20_65 V20 V65 19389.405637560645
L20_65 V20 V65 -9.3595624646145e-11
C20_65 V20 V65 -3.186399960033549e-21

R20_66 V20 V66 13910.332443138219
L20_66 V20 V66 3.5930974989383e-11
C20_66 V20 V66 1.0079015343567868e-20

R20_67 V20 V67 226725.73225904067
L20_67 V20 V67 -1.5594594812354036e-10
C20_67 V20 V67 4.327578615582799e-21

R20_68 V20 V68 -6578.578437157611
L20_68 V20 V68 -2.6247449859019437e-10
C20_68 V20 V68 1.2375133621160959e-20

R20_69 V20 V69 19922.5217402556
L20_69 V20 V69 1.6865615476622e-10
C20_69 V20 V69 -1.871155637045028e-21

R20_70 V20 V70 -26323.644545263665
L20_70 V20 V70 1.8062451567342897e-11
C20_70 V20 V70 3.3619083657201828e-21

R20_71 V20 V71 -541127.3236561156
L20_71 V20 V71 -1.2798553682652528e-10
C20_71 V20 V71 -1.9683775884296976e-21

R20_72 V20 V72 84660.79914500291
L20_72 V20 V72 6.355027099908758e-11
C20_72 V20 V72 1.929803052029577e-21

R20_73 V20 V73 -24514.836885517492
L20_73 V20 V73 2.4503653419030713e-11
C20_73 V20 V73 1.5730271026188158e-21

R20_74 V20 V74 -252139.21187159416
L20_74 V20 V74 8.103912480202721e-11
C20_74 V20 V74 3.704821886391229e-21

R20_75 V20 V75 47256.863422166665
L20_75 V20 V75 -4.7755476115081126e-11
C20_75 V20 V75 4.2325558300740106e-21

R20_76 V20 V76 50370.8658113236
L20_76 V20 V76 2.6326425682120985e-11
C20_76 V20 V76 4.417386508946693e-21

R20_77 V20 V77 92947.74384977426
L20_77 V20 V77 -3.922641323517696e-11
C20_77 V20 V77 -7.246304684566541e-21

R20_78 V20 V78 907456.595729205
L20_78 V20 V78 4.340192448843851e-11
C20_78 V20 V78 -3.659604796407626e-21

R20_79 V20 V79 593867.6345462671
L20_79 V20 V79 3.3770449950974683e-11
C20_79 V20 V79 2.441541190916621e-21

R20_80 V20 V80 -165086.5224542966
L20_80 V20 V80 -1.0875054615728234e-11
C20_80 V20 V80 -1.4413164064145548e-20

R20_81 V20 V81 390976.14961900236
L20_81 V20 V81 6.707357061396914e-12
C20_81 V20 V81 3.205766054725524e-20

R20_82 V20 V82 -110031.50816807403
L20_82 V20 V82 -1.1010530551984453e-11
C20_82 V20 V82 -5.61974407453796e-22

R20_83 V20 V83 -365734.06911813054
L20_83 V20 V83 -8.254969993864803e-12
C20_83 V20 V83 -1.552067474529862e-20

R20_84 V20 V84 78127.93496779118
L20_84 V20 V84 1.347133670397936e-10
C20_84 V20 V84 -4.0107157474166044e-21

R20_85 V20 V85 -311885.97207517794
L20_85 V20 V85 1.6775310143371755e-11
C20_85 V20 V85 7.48850811677247e-22

R20_86 V20 V86 -72643.01893072782
L20_86 V20 V86 3.018947374103003e-11
C20_86 V20 V86 -3.305446877217183e-21

R20_87 V20 V87 159730.1871723591
L20_87 V20 V87 1.1876463614976678e-11
C20_87 V20 V87 5.54222211195987e-21

R20_88 V20 V88 1337146.0196650263
L20_88 V20 V88 2.1381729609981218e-11
C20_88 V20 V88 6.270991353994469e-21

R20_89 V20 V89 306441.57606864994
L20_89 V20 V89 -1.7824639781869845e-11
C20_89 V20 V89 -1.72721487636866e-21

R20_90 V20 V90 -238339681.7374681
L20_90 V20 V90 -8.36353433710072e-11
C20_90 V20 V90 2.1671125290965494e-21

R20_91 V20 V91 245767.75936813667
L20_91 V20 V91 -2.3680786042221176e-11
C20_91 V20 V91 9.555431202194653e-21

R20_92 V20 V92 -100026.35053939259
L20_92 V20 V92 -6.2000015067891466e-12
C20_92 V20 V92 -3.046113997283403e-20

R20_93 V20 V93 -50451.29246752129
L20_93 V20 V93 4.740817944960058e-11
C20_93 V20 V93 4.47749083376966e-21

R20_94 V20 V94 -89191.82500313519
L20_94 V20 V94 1.4025843582931174e-11
C20_94 V20 V94 9.216667474956032e-21

R20_95 V20 V95 11387356.462161208
L20_95 V20 V95 -2.4468542256716484e-11
C20_95 V20 V95 1.734569183064567e-21

R20_96 V20 V96 754876.7640801878
L20_96 V20 V96 -6.383609706740258e-12
C20_96 V20 V96 -3.132291917025566e-20

R20_97 V20 V97 169047.4487708619
L20_97 V20 V97 1.9232209944768495e-11
C20_97 V20 V97 8.980715272179336e-21

R20_98 V20 V98 185683.32361578444
L20_98 V20 V98 -1.0453019827844922e-11
C20_98 V20 V98 -1.0669323730270143e-20

R20_99 V20 V99 -129880.79876207793
L20_99 V20 V99 4.1640882434216e-11
C20_99 V20 V99 3.3233706739855743e-21

R20_100 V20 V100 102524.40117649772
L20_100 V20 V100 1.6342454396786523e-11
C20_100 V20 V100 6.496687781210496e-21

R20_101 V20 V101 -77021.34385406262
L20_101 V20 V101 -1.011392276088945e-11
C20_101 V20 V101 -3.050105682652122e-21

R20_102 V20 V102 193681.3624818064
L20_102 V20 V102 -1.4192504732557564e-11
C20_102 V20 V102 9.586024419337615e-22

R20_103 V20 V103 330694.2208756725
L20_103 V20 V103 3.7989021264556296e-11
C20_103 V20 V103 -1.94659871920846e-21

R20_104 V20 V104 -82342.91419079316
L20_104 V20 V104 -1.0922574117985631e-11
C20_104 V20 V104 -1.6829159314127835e-20

R20_105 V20 V105 83023.7493057412
L20_105 V20 V105 9.674353070098556e-12
C20_105 V20 V105 5.162904024559951e-21

R20_106 V20 V106 -1106950.9667088862
L20_106 V20 V106 -7.369247554663014e-12
C20_106 V20 V106 -2.2472482608308984e-21

R20_107 V20 V107 -1269949.8516602437
L20_107 V20 V107 -1.720980044301081e-11
C20_107 V20 V107 -1.754663759114359e-21

R20_108 V20 V108 37071.153198973014
L20_108 V20 V108 7.886397759625333e-12
C20_108 V20 V108 8.576020194143249e-21

R20_109 V20 V109 -97749.19536097109
L20_109 V20 V109 -1.2789260187227323e-11
C20_109 V20 V109 -1.5751099741906883e-20

R20_110 V20 V110 92415.32511516947
L20_110 V20 V110 7.7995167211544e-12
C20_110 V20 V110 2.8336370784641015e-21

R20_111 V20 V111 99403.70011991009
L20_111 V20 V111 1.3653022497746572e-11
C20_111 V20 V111 8.039391504346997e-21

R20_112 V20 V112 51909.016149023715
L20_112 V20 V112 -9.826942720027956e-12
C20_112 V20 V112 -6.353702627956604e-21

R20_113 V20 V113 47527.11785976186
L20_113 V20 V113 3.618179256137911e-10
C20_113 V20 V113 9.403539518824161e-21

R20_114 V20 V114 45618.470714198134
L20_114 V20 V114 -1.2555724302556166e-11
C20_114 V20 V114 -7.564763834741936e-21

R20_115 V20 V115 247966.56861298694
L20_115 V20 V115 -3.376799014845186e-11
C20_115 V20 V115 -1.690109250016743e-21

R20_116 V20 V116 312436.37467254204
L20_116 V20 V116 1.1029230289063124e-11
C20_116 V20 V116 1.0509507413701425e-20

R20_117 V20 V117 -210754.83457152708
L20_117 V20 V117 3.1025290880547957e-10
C20_117 V20 V117 -9.329938927768079e-21

R20_118 V20 V118 -180062.2558501276
L20_118 V20 V118 3.012606964236559e-11
C20_118 V20 V118 -6.659846817206558e-21

R20_119 V20 V119 219619.6435215876
L20_119 V20 V119 9.201986457305733e-12
C20_119 V20 V119 1.5402548183586485e-20

R20_120 V20 V120 -1100629.6662721164
L20_120 V20 V120 1.4623677322114567e-11
C20_120 V20 V120 1.1183869911932053e-20

R20_121 V20 V121 35014.329313632865
L20_121 V20 V121 -7.68245397661022e-11
C20_121 V20 V121 3.638940115256347e-21

R20_122 V20 V122 14377.06754316721
L20_122 V20 V122 -4.9814988003514307e-11
C20_122 V20 V122 1.1177265589209691e-21

R20_123 V20 V123 33652.75800623512
L20_123 V20 V123 7.501268527256003e-11
C20_123 V20 V123 1.770853586551624e-21

R20_124 V20 V124 48050.40860410082
L20_124 V20 V124 1.3139289103238407e-11
C20_124 V20 V124 1.0362303052813908e-20

R20_125 V20 V125 -37716.734041504475
L20_125 V20 V125 2.6935212496259685e-11
C20_125 V20 V125 1.6132448860955938e-21

R20_126 V20 V126 -19233.30241890654
L20_126 V20 V126 -1.3977273101693045e-09
C20_126 V20 V126 1.3382396091618009e-23

R20_127 V20 V127 43538.28606326186
L20_127 V20 V127 -2.723968146139539e-10
C20_127 V20 V127 7.232505350888199e-22

R20_128 V20 V128 -181137.61298741834
L20_128 V20 V128 -2.5428691430954508e-11
C20_128 V20 V128 -5.9927462349086165e-21

R20_129 V20 V129 28578.425648167264
L20_129 V20 V129 4.9864106534398925e-11
C20_129 V20 V129 -8.743293289520599e-22

R20_130 V20 V130 -23645.811175107116
L20_130 V20 V130 -6.638165332857471e-11
C20_130 V20 V130 -6.174066484499464e-21

R20_131 V20 V131 -22035.01211620079
L20_131 V20 V131 -2.9267851980904885e-11
C20_131 V20 V131 -2.5955125824259118e-21

R20_132 V20 V132 -79307.92722986217
L20_132 V20 V132 3.226499557699712e-11
C20_132 V20 V132 5.415576130558633e-21

R20_133 V20 V133 -100157.57282470564
L20_133 V20 V133 -2.256364355643852e-11
C20_133 V20 V133 1.504280287651346e-22

R20_134 V20 V134 -126934.50939860482
L20_134 V20 V134 1.4160106184323075e-10
C20_134 V20 V134 1.0071884521772283e-21

R20_135 V20 V135 46560.31054496346
L20_135 V20 V135 2.0306710435547804e-10
C20_135 V20 V135 -1.0316232838375387e-23

R20_136 V20 V136 -196157.26001302758
L20_136 V20 V136 6.138041911590815e-10
C20_136 V20 V136 5.671286046522125e-21

R20_137 V20 V137 -60444.66658888404
L20_137 V20 V137 2.8511567691471093e-11
C20_137 V20 V137 -1.3929752035552672e-21

R20_138 V20 V138 -14340.538535606478
L20_138 V20 V138 7.679907566860033e-11
C20_138 V20 V138 4.68240980604073e-21

R20_139 V20 V139 35082.40904019955
L20_139 V20 V139 -9.15166679710374e-11
C20_139 V20 V139 3.0404227389386062e-21

R20_140 V20 V140 -137293.35730436453
L20_140 V20 V140 1.1415701697543066e-10
C20_140 V20 V140 3.774761964288531e-21

R20_141 V20 V141 -218132.54407343853
L20_141 V20 V141 4.18621283415974e-11
C20_141 V20 V141 3.510051820993874e-21

R20_142 V20 V142 -42051.2944931342
L20_142 V20 V142 4.0048393237782247e-10
C20_142 V20 V142 2.381047147906892e-21

R20_143 V20 V143 -69089.46688415445
L20_143 V20 V143 -1.7003054571155418e-10
C20_143 V20 V143 -4.9626018534877495e-22

R20_144 V20 V144 69503.15338586505
L20_144 V20 V144 -4.898393155245603e-11
C20_144 V20 V144 -3.867482079555713e-21

R21_21 V21 0 -525.1938568020133
L21_21 V21 0 -7.773552232300757e-14
C21_21 V21 0 4.2060434394389155e-19

R21_22 V21 V22 528418.1336567977
L21_22 V21 V22 9.360717242335395e-12
C21_22 V21 V22 -3.622501567776438e-21

R21_23 V21 V23 167687.06573193675
L21_23 V21 V23 1.1456591728982672e-11
C21_23 V21 V23 -9.779824007162075e-22

R21_24 V21 V24 1308857.1901042655
L21_24 V21 V24 9.673111407821857e-12
C21_24 V21 V24 -1.291199054212055e-21

R21_25 V21 V25 -13155.21602339235
L21_25 V21 V25 -3.494727286191874e-12
C21_25 V21 V25 -5.754285894567268e-20

R21_26 V21 V26 -43558.23413883088
L21_26 V21 V26 8.644000947159234e-11
C21_26 V21 V26 -8.895819368150729e-21

R21_27 V21 V27 -42614.69408643973
L21_27 V21 V27 -2.6205199491025902e-11
C21_27 V21 V27 -8.278747910659954e-21

R21_28 V21 V28 -66874.4904925492
L21_28 V21 V28 -5.030525236838991e-11
C21_28 V21 V28 -4.427860886654958e-21

R21_29 V21 V29 8092.117747417247
L21_29 V21 V29 -1.3338739125251386e-12
C21_29 V21 V29 2.4540456357297517e-20

R21_30 V21 V30 32228.022602859102
L21_30 V21 V30 2.5714536291295e-10
C21_30 V21 V30 1.9482063174494626e-20

R21_31 V21 V31 48448.498520517314
L21_31 V21 V31 -1.1947394157322435e-10
C21_31 V21 V31 6.0137594589742565e-21

R21_32 V21 V32 51533.64938186854
L21_32 V21 V32 4.3229729867705083e-11
C21_32 V21 V32 1.1679394962367732e-20

R21_33 V21 V33 13440.821638494072
L21_33 V21 V33 1.4347890291767377e-12
C21_33 V21 V33 1.3446141469139407e-20

R21_34 V21 V34 -23451.56678520386
L21_34 V21 V34 -3.3612710922384937e-12
C21_34 V21 V34 -4.232651392585661e-21

R21_35 V21 V35 24883.971879685112
L21_35 V21 V35 2.4192376613337238e-12
C21_35 V21 V35 1.1127955823429598e-21

R21_36 V21 V36 -34171.926689713684
L21_36 V21 V36 -6.981901568055105e-12
C21_36 V21 V36 -5.3236518608032974e-21

R21_37 V21 V37 -59503.18934406599
L21_37 V21 V37 -1.0092970265696714e-12
C21_37 V21 V37 5.19155781671938e-20

R21_38 V21 V38 -152639.21038960924
L21_38 V21 V38 4.136487248819336e-11
C21_38 V21 V38 2.360914761017525e-21

R21_39 V21 V39 -23865.512950084787
L21_39 V21 V39 -1.1736872007699123e-12
C21_39 V21 V39 2.7893690383596093e-20

R21_40 V21 V40 -1596469.3363668316
L21_40 V21 V40 3.720165271374455e-11
C21_40 V21 V40 -1.6384063964450426e-21

R21_41 V21 V41 5550.201508772941
L21_41 V21 V41 2.840763696177723e-13
C21_41 V21 V41 -1.8581857491362912e-19

R21_42 V21 V42 13680.08611416498
L21_42 V21 V42 3.958844153032208e-13
C21_42 V21 V42 -1.3417246864189048e-19

R21_43 V21 V43 26903.02554070656
L21_43 V21 V43 7.805744351326969e-13
C21_43 V21 V43 -6.041826914788346e-20

R21_44 V21 V44 -171636.12916977084
L21_44 V21 V44 2.6080762818033274e-11
C21_44 V21 V44 2.9838758550161615e-21

R21_45 V21 V45 4726.729226652921
L21_45 V21 V45 -7.664435279423329e-13
C21_45 V21 V45 1.431298571817223e-19

R21_46 V21 V46 5141.823424783919
L21_46 V21 V46 -5.384039513833096e-12
C21_46 V21 V46 7.687359385479631e-20

R21_47 V21 V47 8176.092844816451
L21_47 V21 V47 1.626997454480065e-11
C21_47 V21 V47 2.2348851800152147e-20

R21_48 V21 V48 -38288.83199951152
L21_48 V21 V48 -4.3306164774486775e-12
C21_48 V21 V48 4.127288350972046e-21

R21_49 V21 V49 -9947.624352982486
L21_49 V21 V49 3.153162357742828e-12
C21_49 V21 V49 -3.046808132605926e-20

R21_50 V21 V50 25020.530193821432
L21_50 V21 V50 1.3686505398260807e-12
C21_50 V21 V50 -3.018704783032178e-20

R21_51 V21 V51 -19993.056661638097
L21_51 V21 V51 -1.6509333484951156e-12
C21_51 V21 V51 2.821666221849912e-20

R21_52 V21 V52 -10312.715298443238
L21_52 V21 V52 7.52643076500554e-13
C21_52 V21 V52 -8.52428062597232e-20

R21_53 V21 V53 -25457.821149429456
L21_53 V21 V53 1.061488886426731e-12
C21_53 V21 V53 -4.481432640885212e-20

R21_54 V21 V54 12778.48949905665
L21_54 V21 V54 2.4853848555393903e-12
C21_54 V21 V54 -1.004191892141525e-20

R21_55 V21 V55 11886.162641201734
L21_55 V21 V55 1.2526695037157537e-12
C21_55 V21 V55 -2.4894086534507534e-20

R21_56 V21 V56 21527.48706350681
L21_56 V21 V56 2.0445161997480917e-12
C21_56 V21 V56 -2.0903931191617493e-20

R21_57 V21 V57 1079.1697504964723
L21_57 V21 V57 3.2581133752468346e-13
C21_57 V21 V57 8.131743631415468e-21

R21_58 V21 V58 4798.486078829252
L21_58 V21 V58 1.629663945938622e-12
C21_58 V21 V58 8.897481858972151e-21

R21_59 V21 V59 17015.523107774297
L21_59 V21 V59 1.753223706738395e-10
C21_59 V21 V59 1.1340989924797004e-20

R21_60 V21 V60 7783.888572727881
L21_60 V21 V60 2.3139749105499032e-12
C21_60 V21 V60 3.1966324199049453e-21

R21_61 V21 V61 -3292.450285975497
L21_61 V21 V61 -1.241203411873803e-11
C21_61 V21 V61 -4.366138981566815e-20

R21_62 V21 V62 -3482.822488230624
L21_62 V21 V62 -5.050155006131831e-12
C21_62 V21 V62 -4.033405390641694e-20

R21_63 V21 V63 -63359.672540333726
L21_63 V21 V63 2.8069929457147703e-11
C21_63 V21 V63 -7.55299082149922e-21

R21_64 V21 V64 208265.33927202242
L21_64 V21 V64 9.662213455675201e-12
C21_64 V21 V64 -3.0403146213783225e-21

R21_65 V21 V65 3389.410948052226
L21_65 V21 V65 5.701448572785899e-13
C21_65 V21 V65 -9.697267388785505e-21

R21_66 V21 V66 4219.649559685791
L21_66 V21 V66 6.668999347090055e-13
C21_66 V21 V66 -3.87111441933554e-21

R21_67 V21 V67 20090.59834835691
L21_67 V21 V67 3.292388787191402e-12
C21_67 V21 V67 -6.2341050514012805e-21

R21_68 V21 V68 50521.816758570545
L21_68 V21 V68 4.8595183404003385e-12
C21_68 V21 V68 -4.584064466341992e-21

R21_69 V21 V69 -38058.479735972054
L21_69 V21 V69 -2.6782743236613642e-12
C21_69 V21 V69 4.510180312659152e-21

R21_70 V21 V70 -24707.027165675205
L21_70 V21 V70 -3.4704231493891124e-12
C21_70 V21 V70 -1.5119557493676663e-20

R21_71 V21 V71 60718.99526896353
L21_71 V21 V71 -1.044232341541987e-11
C21_71 V21 V71 -5.4029151559802306e-21

R21_72 V21 V72 -20437.4559759319
L21_72 V21 V72 -1.76295737627629e-12
C21_72 V21 V72 -1.1099716837040994e-20

R21_73 V21 V73 214136.39493310542
L21_73 V21 V73 -1.2603468665322208e-11
C21_73 V21 V73 -1.1401898816732322e-20

R21_74 V21 V74 -29495.991985705656
L21_74 V21 V74 -2.5275118230115986e-12
C21_74 V21 V74 5.7408691768695104e-21

R21_75 V21 V75 27621.629303699705
L21_75 V21 V75 3.038331699270692e-12
C21_75 V21 V75 -1.3318831265104511e-21

R21_76 V21 V76 40058.829791767945
L21_76 V21 V76 2.9304857880545975e-12
C21_76 V21 V76 -4.891979324993527e-21

R21_77 V21 V77 172979.9035923949
L21_77 V21 V77 4.781178836980659e-12
C21_77 V21 V77 -1.1991630598924924e-22

R21_78 V21 V78 -62585.716860935434
L21_78 V21 V78 2.900880682420526e-11
C21_78 V21 V78 -7.451937019986444e-21

R21_79 V21 V79 -212461.62066143408
L21_79 V21 V79 -2.9792667578004444e-11
C21_79 V21 V79 6.062680175216473e-21

R21_80 V21 V80 -87109.93426386669
L21_80 V21 V80 1.2140793297863357e-11
C21_80 V21 V80 -9.665262195394765e-22

R21_81 V21 V81 204924.349550523
L21_81 V21 V81 -6.318931784215526e-12
C21_81 V21 V81 2.1183157961714005e-21

R21_82 V21 V82 -84766.16190119596
L21_82 V21 V82 2.3860145968572897e-12
C21_82 V21 V82 2.125024149434053e-20

R21_83 V21 V83 79046.0233106186
L21_83 V21 V83 -4.302067109156558e-11
C21_83 V21 V83 -2.756854197489367e-21

R21_84 V21 V84 70991.03159399159
L21_84 V21 V84 -2.5600860985857595e-12
C21_84 V21 V84 -9.250250308792601e-21

R21_85 V21 V85 -194192.07933395082
L21_85 V21 V85 -2.71538940787453e-12
C21_85 V21 V85 -1.0325586635835417e-20

R21_86 V21 V86 -109769.04961741144
L21_86 V21 V86 -4.46465568515492e-12
C21_86 V21 V86 -9.94335149183123e-21

R21_87 V21 V87 -703567.5736574243
L21_87 V21 V87 -3.459091025424998e-12
C21_87 V21 V87 -9.387224988500022e-21

R21_88 V21 V88 -84286.70327597702
L21_88 V21 V88 -3.9382923288793346e-11
C21_88 V21 V88 -2.3717126020778927e-22

R21_89 V21 V89 86540.99394528121
L21_89 V21 V89 1.5649026309648434e-12
C21_89 V21 V89 2.219669460101049e-20

R21_90 V21 V90 -728264.3375412798
L21_90 V21 V90 9.46405195924809e-12
C21_90 V21 V90 -4.708031109927584e-21

R21_91 V21 V91 292559.33598901593
L21_91 V21 V91 4.189754588680135e-12
C21_91 V21 V91 1.5095253270076937e-20

R21_92 V21 V92 658483.1958808803
L21_92 V21 V92 7.79443456148614e-12
C21_92 V21 V92 -1.4421134566010756e-21

R21_93 V21 V93 -18392.703759072534
L21_93 V21 V93 -1.54447366588146e-11
C21_93 V21 V93 7.122776846596457e-21

R21_94 V21 V94 -33750.494086292594
L21_94 V21 V94 -3.965374106105509e-12
C21_94 V21 V94 -8.126667984116842e-21

R21_95 V21 V95 430419.4922119996
L21_95 V21 V95 1.385895512362471e-11
C21_95 V21 V95 9.87714925414296e-21

R21_96 V21 V96 99428.19623719332
L21_96 V21 V96 -3.07541591948865e-11
C21_96 V21 V96 -3.962324191843623e-21

R21_97 V21 V97 -79775.83543162329
L21_97 V21 V97 4.828067217597173e-12
C21_97 V21 V97 -2.6808404416561245e-21

R21_98 V21 V98 -133848.04355865062
L21_98 V21 V98 1.84708636574034e-12
C21_98 V21 V98 4.962844862436186e-21

R21_99 V21 V99 -57592.2021925199
L21_99 V21 V99 1.0789379461220757e-10
C21_99 V21 V99 -9.664368604720173e-23

R21_100 V21 V100 162504.33749993026
L21_100 V21 V100 -2.11916119562745e-11
C21_100 V21 V100 2.1293426459369806e-23

R21_101 V21 V101 -78267.65566642319
L21_101 V21 V101 1.527279639910326e-12
C21_101 V21 V101 1.8799894408288908e-20

R21_102 V21 V102 -63473.52490785559
L21_102 V21 V102 2.247369338911465e-12
C21_102 V21 V102 -2.593639319146487e-21

R21_103 V21 V103 -233670.578156974
L21_103 V21 V103 1.0682752316096445e-11
C21_103 V21 V103 8.385996222757961e-21

R21_104 V21 V104 -560903.5555653331
L21_104 V21 V104 -1.236615120739995e-11
C21_104 V21 V104 -4.472173339828656e-21

R21_105 V21 V105 62924.9165687287
L21_105 V21 V105 -4.555861222552417e-12
C21_105 V21 V105 -1.2965453282926546e-21

R21_106 V21 V106 74485.5584239963
L21_106 V21 V106 8.127130620392157e-12
C21_106 V21 V106 1.1633066920205006e-20

R21_107 V21 V107 -156420.93459515693
L21_107 V21 V107 1.0438509929180382e-11
C21_107 V21 V107 -1.0780546059021979e-20

R21_108 V21 V108 70751.75524901101
L21_108 V21 V108 -2.5302679327962527e-12
C21_108 V21 V108 -2.769474757255835e-21

R21_109 V21 V109 237059.5663619034
L21_109 V21 V109 -1.51607181976339e-11
C21_109 V21 V109 -4.712060864635374e-21

R21_110 V21 V110 1190098.4563272577
L21_110 V21 V110 -2.31495616726601e-12
C21_110 V21 V110 -1.4491805623327173e-20

R21_111 V21 V111 58867.64712713703
L21_111 V21 V111 8.145068093081255e-12
C21_111 V21 V111 3.1988681719268267e-21

R21_112 V21 V112 33754.96509236359
L21_112 V21 V112 1.3523293094755233e-12
C21_112 V21 V112 7.203312445762569e-21

R21_113 V21 V113 41404.424460773276
L21_113 V21 V113 3.106519603779586e-12
C21_113 V21 V113 7.045694074394613e-21

R21_114 V21 V114 1143418.4639894562
L21_114 V21 V114 5.1257074881637245e-12
C21_114 V21 V114 9.075425227123393e-21

R21_115 V21 V115 -86809.4723971271
L21_115 V21 V115 -1.7648946262283098e-11
C21_115 V21 V115 -5.543684585989589e-21

R21_116 V21 V116 -264132.96316817234
L21_116 V21 V116 -2.7179306560006177e-12
C21_116 V21 V116 8.409709992363513e-22

R21_117 V21 V117 -50580.253270646295
L21_117 V21 V117 -3.0339956766234758e-12
C21_117 V21 V117 -7.034278844975703e-21

R21_118 V21 V118 108541.20684652108
L21_118 V21 V118 -3.3066704256763804e-12
C21_118 V21 V118 -5.913267692537409e-21

R21_119 V21 V119 44167.17535269184
L21_119 V21 V119 -1.534473577119852e-11
C21_119 V21 V119 -5.785496332841262e-21

R21_120 V21 V120 -48186.007591621405
L21_120 V21 V120 -2.8848026836706363e-12
C21_120 V21 V120 1.913935556714287e-21

R21_121 V21 V121 21056.182357360278
L21_121 V21 V121 1.8828555228938513e-12
C21_121 V21 V121 2.0179338335074539e-22

R21_122 V21 V122 16349.275520656907
L21_122 V21 V122 1.9038433737377588e-12
C21_122 V21 V122 1.9868607784522816e-21

R21_123 V21 V123 201657.27964653962
L21_123 V21 V123 1.3360866479681637e-11
C21_123 V21 V123 1.000690907969791e-21

R21_124 V21 V124 -267682.6388312736
L21_124 V21 V124 1.5842478448784288e-11
C21_124 V21 V124 -7.174457578710306e-23

R21_125 V21 V125 -15773.26545786812
L21_125 V21 V125 -1.2760266844785092e-12
C21_125 V21 V125 -1.8138876442612404e-21

R21_126 V21 V126 -19184.98913450457
L21_126 V21 V126 -4.955444595549404e-12
C21_126 V21 V126 -1.9636864034769933e-21

R21_127 V21 V127 1573557.3708742994
L21_127 V21 V127 2.58094148445566e-10
C21_127 V21 V127 -3.057831087630996e-21

R21_128 V21 V128 -121908.95050953579
L21_128 V21 V128 3.574739583534471e-11
C21_128 V21 V128 -2.757373619059594e-21

R21_129 V21 V129 -82111.66394110324
L21_129 V21 V129 -8.975284064534934e-11
C21_129 V21 V129 -4.586975945633914e-21

R21_130 V21 V130 -82343.90839863269
L21_130 V21 V130 -9.485507263191665e-12
C21_130 V21 V130 -4.479156419829615e-21

R21_131 V21 V131 -56155.653528416144
L21_131 V21 V131 -1.0675089675112478e-11
C21_131 V21 V131 -3.3988176165912855e-21

R21_132 V21 V132 -412463.12608434696
L21_132 V21 V132 -2.4445399336141912e-11
C21_132 V21 V132 2.3676645609819755e-21

R21_133 V21 V133 -155691.4940353394
L21_133 V21 V133 -7.307333741049593e-12
C21_133 V21 V133 3.2427172525139814e-21

R21_134 V21 V134 134231.08552162698
L21_134 V21 V134 -5.020473426037691e-12
C21_134 V21 V134 -1.4185261381993954e-21

R21_135 V21 V135 46750.978728912996
L21_135 V21 V135 7.255926315529955e-11
C21_135 V21 V135 2.4516619284976707e-21

R21_136 V21 V136 -183602.29735452798
L21_136 V21 V136 -2.12258304490779e-11
C21_136 V21 V136 3.877981205147319e-22

R21_137 V21 V137 -22447.050916841377
L21_137 V21 V137 -2.739957195684663e-12
C21_137 V21 V137 -5.4657052292107414e-21

R21_138 V21 V138 -32083.826660396116
L21_138 V21 V138 -3.916655791158371e-12
C21_138 V21 V138 9.672873677738087e-22

R21_139 V21 V139 -402175.30446149525
L21_139 V21 V139 5.419444795155457e-11
C21_139 V21 V139 -2.64087584311265e-22

R21_140 V21 V140 -83213.17144465644
L21_140 V21 V140 -5.403412222689818e-12
C21_140 V21 V140 -4.319411270136445e-21

R21_141 V21 V141 -24259.46171102982
L21_141 V21 V141 -1.1820832805318885e-11
C21_141 V21 V141 -5.8515347180963334e-21

R21_142 V21 V142 70600.06036857444
L21_142 V21 V142 -1.079213493442703e-11
C21_142 V21 V142 1.7645331735287225e-21

R21_143 V21 V143 104424.64617432059
L21_143 V21 V143 2.5355162263778927e-11
C21_143 V21 V143 3.457586910379582e-21

R21_144 V21 V144 27648.520550446032
L21_144 V21 V144 1.573990242355445e-11
C21_144 V21 V144 1.4041457947948393e-21

R22_22 V22 0 7568.775676874245
L22_22 V22 0 1.9612004880578952e-13
C22_22 V22 0 -2.3427063592631236e-19

R22_23 V22 V23 -1706838.8139168527
L22_23 V22 V23 7.20445832051486e-12
C22_23 V22 V23 1.2544585154633644e-21

R22_24 V22 V24 1244396.1768021185
L22_24 V22 V24 7.32147605213455e-12
C22_24 V22 V24 4.1559515169764773e-22

R22_25 V22 V25 102180.32042719802
L22_25 V22 V25 1.1400582728137903e-11
C22_25 V22 V25 8.113098619002669e-21

R22_26 V22 V26 -1485914.4189394077
L22_26 V22 V26 -2.048788281010356e-12
C22_26 V22 V26 5.589886148318522e-22

R22_27 V22 V27 254622.57276913934
L22_27 V22 V27 -8.771289950984123e-12
C22_27 V22 V27 2.4506731993625204e-21

R22_28 V22 V28 865776.1957972856
L22_28 V22 V28 -1.5374602150088922e-11
C22_28 V22 V28 1.513820775615921e-21

R22_29 V22 V29 -58707.27933481238
L22_29 V22 V29 5.661480294836498e-12
C22_29 V22 V29 -6.672783479111068e-21

R22_30 V22 V30 -554975.4000844863
L22_30 V22 V30 -2.1457792051716355e-12
C22_30 V22 V30 3.1041716365038696e-21

R22_31 V22 V31 -207368.6170537459
L22_31 V22 V31 6.92523829882123e-12
C22_31 V22 V31 -5.586396116162948e-21

R22_32 V22 V32 -283383.4470351544
L22_32 V22 V32 9.292328888875385e-12
C22_32 V22 V32 -3.6131740832798464e-21

R22_33 V22 V33 -182446.6469578729
L22_33 V22 V33 -5.134356879253977e-12
C22_33 V22 V33 -5.63064360413445e-22

R22_34 V22 V34 -268153755.77702048
L22_34 V22 V34 1.2793862456973639e-11
C22_34 V22 V34 -1.939444883414187e-21

R22_35 V22 V35 62842076.37331157
L22_35 V22 V35 -1.1773273167317764e-11
C22_35 V22 V35 4.332563434027104e-21

R22_36 V22 V36 426479.3782537713
L22_36 V22 V36 -4.630369436422102e-11
C22_36 V22 V36 1.725770908404971e-21

R22_37 V22 V37 -216897.87189673085
L22_37 V22 V37 4.450306697224491e-12
C22_37 V22 V37 -1.5846140938123928e-20

R22_38 V22 V38 69756.45074835733
L22_38 V22 V38 -3.716542309746792e-12
C22_38 V22 V38 1.6775777875741494e-20

R22_39 V22 V39 -534129.8292130302
L22_39 V22 V39 6.6483604564927406e-12
C22_39 V22 V39 -1.4564126282919566e-20

R22_40 V22 V40 -212064.3282925421
L22_40 V22 V40 1.0949638991748743e-11
C22_40 V22 V40 -8.408865435967412e-21

R22_41 V22 V41 106570.58849313331
L22_41 V22 V41 -1.112518349498815e-12
C22_41 V22 V41 7.175361362944563e-20

R22_42 V22 V42 -30150.92389533191
L22_42 V22 V42 3.4765700986217928e-12
C22_42 V22 V42 -2.4083197103709725e-20

R22_43 V22 V43 56397.4039999346
L22_43 V22 V43 -3.4234253831988945e-12
C22_43 V22 V43 2.5493234512411996e-20

R22_44 V22 V44 223040.21407445817
L22_44 V22 V44 -1.807745055865603e-11
C22_44 V22 V44 4.356675319002288e-21

R22_45 V22 V45 -32388.23529668886
L22_45 V22 V45 4.826383741859924e-12
C22_45 V22 V45 -4.0833284885578043e-20

R22_46 V22 V46 -170377.94753258643
L22_46 V22 V46 -9.367466342931695e-12
C22_46 V22 V46 1.7896373444877195e-20

R22_47 V22 V47 -69895.95426621521
L22_47 V22 V47 -5.029238376500181e-12
C22_47 V22 V47 -6.912925535146219e-21

R22_48 V22 V48 1169121.6701013255
L22_48 V22 V48 -9.64411325112415e-12
C22_48 V22 V48 2.2033375106137525e-21

R22_49 V22 V49 88016.02002284415
L22_49 V22 V49 -3.1320539023555495e-11
C22_49 V22 V49 1.4438359969373593e-20

R22_50 V22 V50 33529222.232322544
L22_50 V22 V50 2.2237757191347335e-11
C22_50 V22 V50 -1.6930227032710634e-21

R22_51 V22 V51 -699076.2974127338
L22_51 V22 V51 -4.178733148083019e-12
C22_51 V22 V51 1.8442937513468234e-20

R22_52 V22 V52 91794.4965684311
L22_52 V22 V52 -1.13776463712529e-11
C22_52 V22 V52 1.9156541297897213e-20

R22_53 V22 V53 69348.55107070436
L22_53 V22 V53 -2.238018440561341e-12
C22_53 V22 V53 2.6568969547781827e-20

R22_54 V22 V54 -97558.71021514352
L22_54 V22 V54 -1.5475091077306424e-11
C22_54 V22 V54 -6.924603206977535e-21

R22_55 V22 V55 -708349.39453365
L22_55 V22 V55 -2.0034549364684364e-11
C22_55 V22 V55 1.4380128688728673e-20

R22_56 V22 V56 175036.18722920422
L22_56 V22 V56 -2.7669338214944518e-12
C22_56 V22 V56 3.1922092636589884e-20

R22_57 V22 V57 -11446.027049888586
L22_57 V22 V57 -1.9483219296973675e-12
C22_57 V22 V57 -9.203715123647985e-21

R22_58 V22 V58 -26571.316384645736
L22_58 V22 V58 3.0452283904979572e-12
C22_58 V22 V58 7.071132098603945e-21

R22_59 V22 V59 -248349.7605426739
L22_59 V22 V59 -9.176806506223133e-12
C22_59 V22 V59 1.9550459453473912e-21

R22_60 V22 V60 -55443.68890991617
L22_60 V22 V60 -4.242036408667754e-12
C22_60 V22 V60 3.033969981368009e-21

R22_61 V22 V61 26430.970996830012
L22_61 V22 V61 -4.338283714978704e-12
C22_61 V22 V61 2.6135137611048106e-20

R22_62 V22 V62 39013.96477223447
L22_62 V22 V62 5.616796957087626e-12
C22_62 V22 V62 -3.695423093298602e-21

R22_63 V22 V63 5933599.892083116
L22_63 V22 V63 -2.0064274275326002e-11
C22_63 V22 V63 3.5995935130324675e-20

R22_64 V22 V64 92635.42220310152
L22_64 V22 V64 -3.260321196005404e-12
C22_64 V22 V64 2.476369794015318e-20

R22_65 V22 V65 -36621.07383957526
L22_65 V22 V65 -6.1963602900218716e-12
C22_65 V22 V65 1.5921616735793488e-21

R22_66 V22 V66 -369819.7166797545
L22_66 V22 V66 -2.4786995805125005e-12
C22_66 V22 V66 5.686258386872323e-21

R22_67 V22 V67 -39003.93135403811
L22_67 V22 V67 -3.887506394708945e-12
C22_67 V22 V67 1.1190324368552803e-20

R22_68 V22 V68 -89652.94540223319
L22_68 V22 V68 -2.7734175862757596e-11
C22_68 V22 V68 5.208427346513978e-21

R22_69 V22 V69 -152656.72944632306
L22_69 V22 V69 -1.2017906030628697e-11
C22_69 V22 V69 8.884276591903184e-22

R22_70 V22 V70 48608.890011672
L22_70 V22 V70 -3.7583436402581594e-12
C22_70 V22 V70 1.8346250382321646e-20

R22_71 V22 V71 21640.937393965247
L22_71 V22 V71 -9.413287877434273e-12
C22_71 V22 V71 7.072048264984755e-21

R22_72 V22 V72 -101713.39282768343
L22_72 V22 V72 -3.582112548886358e-11
C22_72 V22 V72 3.816402204501421e-21

R22_73 V22 V73 -52051.77040878926
L22_73 V22 V73 -7.182578379138336e-12
C22_73 V22 V73 2.1830001414045816e-21

R22_74 V22 V74 -154168.6218380479
L22_74 V22 V74 -4.034915523834507e-12
C22_74 V22 V74 3.153261514410688e-21

R22_75 V22 V75 -226983.69863233823
L22_75 V22 V75 4.21551264472922e-12
C22_75 V22 V75 -5.1450263578582786e-21

R22_76 V22 V76 183392.6750517324
L22_76 V22 V76 -1.6050301419761701e-12
C22_76 V22 V76 1.4940630411921956e-20

R22_77 V22 V77 -2737144.937541631
L22_77 V22 V77 -7.179885468788441e-12
C22_77 V22 V77 1.5620159930111943e-22

R22_78 V22 V78 1189762.5869739945
L22_78 V22 V78 -4.044664183038475e-12
C22_78 V22 V78 1.2674995946210196e-21

R22_79 V22 V79 97777.3224750824
L22_79 V22 V79 -1.383028892018685e-12
C22_79 V22 V79 3.5046226338973877e-20

R22_80 V22 V80 -105791.53066328306
L22_80 V22 V80 2.1535721376463998e-12
C22_80 V22 V80 -3.35860386571087e-20

R22_81 V22 V81 740454.1947174509
L22_81 V22 V81 8.47181642259057e-12
C22_81 V22 V81 -4.801003128033213e-22

R22_82 V22 V82 -145268.71193440116
L22_82 V22 V82 3.2464964392816355e-12
C22_82 V22 V82 -1.2161712338685383e-20

R22_83 V22 V83 315201.3690506223
L22_83 V22 V83 1.9949963869421566e-12
C22_83 V22 V83 -2.2049924073749497e-20

R22_84 V22 V84 -211412.47295459206
L22_84 V22 V84 -2.741556266499581e-12
C22_84 V22 V84 1.1951716614952263e-20

R22_85 V22 V85 210179.1201161937
L22_85 V22 V85 -1.841371643732437e-12
C22_85 V22 V85 2.016721205088258e-20

R22_86 V22 V86 -139918.01480759092
L22_86 V22 V86 -9.987645558136196e-12
C22_86 V22 V86 3.840751119953766e-21

R22_87 V22 V87 132178.3696954016
L22_87 V22 V87 -1.9711168553676602e-12
C22_87 V22 V87 1.7353655490607232e-20

R22_88 V22 V88 397101.7702264958
L22_88 V22 V88 5.582852580664996e-11
C22_88 V22 V88 -2.313575914484239e-21

R22_89 V22 V89 -321980.4217013249
L22_89 V22 V89 -5.076112008031516e-11
C22_89 V22 V89 -6.4321353919140146e-21

R22_90 V22 V90 -183824.70232265381
L22_90 V22 V90 1.2851041929816258e-12
C22_90 V22 V90 -3.3927453595031064e-20

R22_91 V22 V91 -1113681.5713806301
L22_91 V22 V91 3.2152093861661846e-12
C22_91 V22 V91 -7.453625943817982e-21

R22_92 V22 V92 -183977.59420460527
L22_92 V22 V92 6.582007748048602e-12
C22_92 V22 V92 -1.6307184396001666e-20

R22_93 V22 V93 140673.08278809136
L22_93 V22 V93 -4.980702241910664e-12
C22_93 V22 V93 5.840732308723504e-21

R22_94 V22 V94 -195147.27285102144
L22_94 V22 V94 1.205043493419386e-11
C22_94 V22 V94 -1.747311161629841e-21

R22_95 V22 V95 -10987102.444928588
L22_95 V22 V95 5.3596999074359904e-12
C22_95 V22 V95 -6.327958957313181e-21

R22_96 V22 V96 -199752.2573729881
L22_96 V22 V96 7.166896197786202e-12
C22_96 V22 V96 -1.2067812767379127e-20

R22_97 V22 V97 -516575.0004389916
L22_97 V22 V97 2.376457574584659e-12
C22_97 V22 V97 -1.4274673517024548e-20

R22_98 V22 V98 -8754673.392375048
L22_98 V22 V98 2.6567558859608618e-12
C22_98 V22 V98 -1.625405652963842e-20

R22_99 V22 V99 -487310.62072744634
L22_99 V22 V99 -2.6187472833688027e-12
C22_99 V22 V99 7.706210184825177e-21

R22_100 V22 V100 -813863.649407034
L22_100 V22 V100 3.163804034330265e-11
C22_100 V22 V100 -2.6508613843600125e-21

R22_101 V22 V101 -382164.72726257937
L22_101 V22 V101 8.15758556997253e-12
C22_101 V22 V101 -6.039597294748063e-21

R22_102 V22 V102 -47510.645400388275
L22_102 V22 V102 5.999470064727374e-13
C22_102 V22 V102 -6.53923762982259e-20

R22_103 V22 V103 58465.68074639382
L22_103 V22 V103 -1.0609002567374424e-12
C22_103 V22 V103 3.9841785707411465e-20

R22_104 V22 V104 -265808.066692713
L22_104 V22 V104 -9.156020994832161e-12
C22_104 V22 V104 -4.574513273164729e-21

R22_105 V22 V105 147353.4402531902
L22_105 V22 V105 -1.4751672885056563e-12
C22_105 V22 V105 1.783133296197174e-20

R22_106 V22 V106 -51795.808726373856
L22_106 V22 V106 9.561198330141073e-13
C22_106 V22 V106 -3.862153177620666e-20

R22_107 V22 V107 -41472.693026126784
L22_107 V22 V107 7.020661757484142e-13
C22_107 V22 V107 -6.263322380332862e-20

R22_108 V22 V108 46811.36440876266
L22_108 V22 V108 -9.25176352431719e-13
C22_108 V22 V108 4.924519846555895e-20

R22_109 V22 V109 120091.20319681456
L22_109 V22 V109 -1.5988351569055498e-12
C22_109 V22 V109 2.1235140356475445e-20

R22_110 V22 V110 57971.264352528015
L22_110 V22 V110 -2.7576128603898142e-12
C22_110 V22 V110 2.4455811035245873e-20

R22_111 V22 V111 258583.9974087685
L22_111 V22 V111 -1.095526505910489e-12
C22_111 V22 V111 2.7514660458925795e-20

R22_112 V22 V112 -111158.13897277178
L22_112 V22 V112 9.56860201187363e-13
C22_112 V22 V112 -3.663016770995751e-20

R22_113 V22 V113 -264910.08708469506
L22_113 V22 V113 1.9937766705084134e-12
C22_113 V22 V113 -1.4269192819888113e-20

R22_114 V22 V114 -491658.72662833467
L22_114 V22 V114 1.935908801949253e-12
C22_114 V22 V114 -1.2626003198253231e-20

R22_115 V22 V115 -120208.88610363573
L22_115 V22 V115 1.3654325717377562e-12
C22_115 V22 V115 -3.712930776253456e-20

R22_116 V22 V116 133696.6330150317
L22_116 V22 V116 -1.7406615673294686e-12
C22_116 V22 V116 3.02693146204732e-20

R22_117 V22 V117 68041.45964956877
L22_117 V22 V117 -2.9785870298917616e-12
C22_117 V22 V117 2.073967218023923e-20

R22_118 V22 V118 543353.902093454
L22_118 V22 V118 -2.221865454131493e-12
C22_118 V22 V118 1.558968860349459e-20

R22_119 V22 V119 2878525.8559171273
L22_119 V22 V119 -1.668188687886056e-12
C22_119 V22 V119 1.8807437331067536e-20

R22_120 V22 V120 40020.54701881984
L22_120 V22 V120 1.6235632209108456e-12
C22_120 V22 V120 1.1713246109098561e-20

R22_121 V22 V121 -569617.602760262
L22_121 V22 V121 6.9211706438135906e-12
C22_121 V22 V121 -1.7658808570565034e-21

R22_122 V22 V122 38012.343620080916
L22_122 V22 V122 1.1654357457942518e-12
C22_122 V22 V122 1.4189990977792932e-21

R22_123 V22 V123 135777.1241120729
L22_123 V22 V123 5.8110860788871275e-12
C22_123 V22 V123 3.362613486102903e-21

R22_124 V22 V124 407363.88914018736
L22_124 V22 V124 -7.511674815561808e-12
C22_124 V22 V124 7.510286542432616e-21

R22_125 V22 V125 94772.37110977725
L22_125 V22 V125 6.54706228482879e-12
C22_125 V22 V125 6.346639413945974e-21

R22_126 V22 V126 -27627.262424767432
L22_126 V22 V126 -8.980289124701667e-13
C22_126 V22 V126 -1.5412942798161046e-21

R22_127 V22 V127 36187.138681554265
L22_127 V22 V127 9.861383792115694e-13
C22_127 V22 V127 -2.4316385262078514e-21

R22_128 V22 V128 414979.2828448093
L22_128 V22 V128 1.351091791755359e-11
C22_128 V22 V128 -1.3462347508039396e-21

R22_129 V22 V129 75705.3623068358
L22_129 V22 V129 2.670387497089786e-12
C22_129 V22 V129 -2.755932344261247e-21

R22_130 V22 V130 -460910.7745663476
L22_130 V22 V130 -1.4358373405972447e-12
C22_130 V22 V130 1.1909651308304989e-20

R22_131 V22 V131 -65819.82596079768
L22_131 V22 V131 1.5881080755277225e-11
C22_131 V22 V131 -1.1515968249738884e-20

R22_132 V22 V132 -153196.41401848782
L22_132 V22 V132 -4.401699022240952e-12
C22_132 V22 V132 1.610438885251643e-21

R22_133 V22 V133 -203556.92253717297
L22_133 V22 V133 4.0202758833874825e-12
C22_133 V22 V133 -8.840285061996906e-21

R22_134 V22 V134 -140865.5820899949
L22_134 V22 V134 -1.037564574088069e-11
C22_134 V22 V134 -3.1738269133002716e-21

R22_135 V22 V135 49687.691235019076
L22_135 V22 V135 1.7001637571834219e-12
C22_135 V22 V135 1.0187064946698611e-20

R22_136 V22 V136 -7102679.568259255
L22_136 V22 V136 2.925855923929094e-11
C22_136 V22 V136 3.6019607441892486e-21

R22_137 V22 V137 163500.60376995103
L22_137 V22 V137 -1.4884624706392997e-11
C22_137 V22 V137 4.4672145506954376e-21

R22_138 V22 V138 -35164.7284661301
L22_138 V22 V138 -9.33569647426606e-13
C22_138 V22 V138 2.5026562733494658e-21

R22_139 V22 V139 30499.47755581889
L22_139 V22 V139 7.153938643342579e-13
C22_139 V22 V139 -6.967925454654727e-21

R22_140 V22 V140 -154198.99177686573
L22_140 V22 V140 -1.857590240623099e-12
C22_140 V22 V140 3.218817200023267e-21

R22_141 V22 V141 -607758.5131174237
L22_141 V22 V141 -3.476864089366681e-12
C22_141 V22 V141 1.866004014763748e-21

R22_142 V22 V142 -93388.87277065073
L22_142 V22 V142 -1.7201120082601747e-12
C22_142 V22 V142 3.63251210749056e-21

R22_143 V22 V143 -78451.24926558042
L22_143 V22 V143 -2.708795222054878e-12
C22_143 V22 V143 5.508339619209993e-21

R22_144 V22 V144 1347070.4582936985
L22_144 V22 V144 4.075185127303798e-12
C22_144 V22 V144 -7.43189604015602e-21

R23_23 V23 0 3351.40234835509
L23_23 V23 0 6.517648002087113e-13
C23_23 V23 0 -1.24358530856589e-19

R23_24 V23 V24 1045354.3565415987
L23_24 V23 V24 1.8707366158598693e-11
C23_24 V23 V24 -4.4310985582392586e-23

R23_25 V23 V25 168086.70046589238
L23_25 V23 V25 9.590657261892538e-12
C23_25 V23 V25 8.774541422448868e-21

R23_26 V23 V26 99309.60671680151
L23_26 V23 V26 6.155197673029354e-12
C23_26 V23 V26 3.496138718085289e-21

R23_27 V23 V27 -564060.9892953979
L23_27 V23 V27 -7.0826807530928504e-12
C23_27 V23 V27 -1.6490536179280085e-20

R23_28 V23 V28 -8781804.061342772
L23_28 V23 V28 -2.839185899961686e-11
C23_28 V23 V28 2.138867101532882e-22

R23_29 V23 V29 -56965.57471566583
L23_29 V23 V29 5.678842350563443e-12
C23_29 V23 V29 -7.892973894499709e-21

R23_30 V23 V30 -151847.4894089235
L23_30 V23 V30 6.822805706628553e-12
C23_30 V23 V30 -1.8263778694530648e-21

R23_31 V23 V31 62804.11931316199
L23_31 V23 V31 -1.9527254246727375e-12
C23_31 V23 V31 -1.1700730463468306e-20

R23_32 V23 V32 1937306.8880246284
L23_32 V23 V32 2.6291580010990543e-11
C23_32 V23 V32 -6.387743474632613e-22

R23_33 V23 V33 391326.6216751498
L23_33 V23 V33 -4.9356894632118225e-12
C23_33 V23 V33 -4.402434557109391e-21

R23_34 V23 V34 223675.69608215112
L23_34 V23 V34 -9.561371224212571e-11
C23_34 V23 V34 -2.5128539178139004e-21

R23_35 V23 V35 65790.23115911784
L23_35 V23 V35 2.3123502024042033e-12
C23_35 V23 V35 8.330303281821226e-21

R23_36 V23 V36 -100210.7668012653
L23_36 V23 V36 -2.0369660882455022e-11
C23_36 V23 V36 1.2620483392578165e-21

R23_37 V23 V37 -32881.27906480879
L23_37 V23 V37 -1.0459362622474244e-11
C23_37 V23 V37 -1.8103225709240392e-20

R23_38 V23 V38 150728.19269375192
L23_38 V23 V38 5.1653130864440475e-12
C23_38 V23 V38 -7.58284907375668e-21

R23_39 V23 V39 203552.1720419422
L23_39 V23 V39 -3.4391507291213668e-12
C23_39 V23 V39 -3.603850972769919e-21

R23_40 V23 V40 991812.2200695493
L23_40 V23 V40 8.459638068678262e-12
C23_40 V23 V40 -1.3999712457694224e-20

R23_41 V23 V41 -45226.91547338891
L23_41 V23 V41 -1.3702774208710028e-12
C23_41 V23 V41 6.953604557391374e-20

R23_42 V23 V42 -491487.49423166807
L23_42 V23 V42 -1.6779746115230833e-12
C23_42 V23 V42 6.883847507714696e-20

R23_43 V23 V43 -474804.26496420597
L23_43 V23 V43 1.648812764238415e-11
C23_43 V23 V43 7.10115116200626e-21

R23_44 V23 V44 -61627.538468647035
L23_44 V23 V44 -2.0686319734712238e-12
C23_44 V23 V44 3.574725651990109e-20

R23_45 V23 V45 -12173.908394505394
L23_45 V23 V45 -1.5013124769802716e-12
C23_45 V23 V45 -3.295009504588676e-20

R23_46 V23 V46 -37857.18987089205
L23_46 V23 V46 1.352023793139735e-12
C23_46 V23 V46 -5.652363996865461e-20

R23_47 V23 V47 40756.33399858576
L23_47 V23 V47 2.2917976803433814e-12
C23_47 V23 V47 -1.2640727502698664e-20

R23_48 V23 V48 -23242.99809147883
L23_48 V23 V48 -2.5059296904508367e-11
C23_48 V23 V48 -1.054212826986141e-20

R23_49 V23 V49 -20743.56348203067
L23_49 V23 V49 -7.952128232869354e-12
C23_49 V23 V49 1.6254361445522936e-21

R23_50 V23 V50 15147.440570288243
L23_50 V23 V50 1.2231837858434794e-11
C23_50 V23 V50 2.4737591930202968e-20

R23_51 V23 V51 -3400692.408074646
L23_51 V23 V51 7.284447124948678e-12
C23_51 V23 V51 -1.760966433059308e-20

R23_52 V23 V52 27509.242932086978
L23_52 V23 V52 -5.9477498223259475e-12
C23_52 V23 V52 3.536843743042055e-20

R23_53 V23 V53 151293.08025952426
L23_53 V23 V53 -6.17095327646306e-12
C23_53 V23 V53 8.838082870003371e-21

R23_54 V23 V54 -86770.66877444889
L23_54 V23 V54 -6.8972746799319865e-12
C23_54 V23 V54 9.63419980468418e-22

R23_55 V23 V55 -18827.686308541033
L23_55 V23 V55 4.3013644504944235e-11
C23_55 V23 V55 -9.042829970885837e-21

R23_56 V23 V56 111729.03236794277
L23_56 V23 V56 -5.3567943259901186e-11
C23_56 V23 V56 1.3230975378835581e-20

R23_57 V23 V57 -6448.800102720748
L23_57 V23 V57 -2.2992636179158052e-12
C23_57 V23 V57 -3.959667025873151e-21

R23_58 V23 V58 -17186.489705003707
L23_58 V23 V58 -2.4686007162723647e-12
C23_58 V23 V58 -7.836304849479089e-21

R23_59 V23 V59 8943.10904591307
L23_59 V23 V59 1.6826605639065961e-12
C23_59 V23 V59 -3.409743398685415e-21

R23_60 V23 V60 -13864.062789861187
L23_60 V23 V60 -1.3505926892256155e-11
C23_60 V23 V60 -4.467122298390922e-21

R23_61 V23 V61 21971.662868882315
L23_61 V23 V61 -1.4898021909235052e-11
C23_61 V23 V61 1.7047463963595295e-20

R23_62 V23 V62 11105.241229150306
L23_62 V23 V62 6.470511890143721e-12
C23_62 V23 V62 2.0873588879135848e-20

R23_63 V23 V63 -290732.4339461386
L23_63 V23 V63 5.2819697942520846e-11
C23_63 V23 V63 -1.5074986265456062e-21

R23_64 V23 V64 56025.850150037004
L23_64 V23 V64 7.093527297944149e-11
C23_64 V23 V64 7.354216198578184e-21

R23_65 V23 V65 -21012.54209487264
L23_65 V23 V65 -6.148867459257986e-12
C23_65 V23 V65 1.5864454288485155e-20

R23_66 V23 V66 -12181.861691064903
L23_66 V23 V66 -1.925932098518673e-12
C23_66 V23 V66 -8.634594893850581e-21

R23_67 V23 V67 130768.17665775846
L23_67 V23 V67 2.1252055806117187e-11
C23_67 V23 V67 -8.434627098541959e-21

R23_68 V23 V68 -30792.83324137185
L23_68 V23 V68 -3.7444069491160485e-11
C23_68 V23 V68 6.291655036428858e-21

R23_69 V23 V69 -50964.335129496
L23_69 V23 V69 2.8631405584115156e-11
C23_69 V23 V69 -7.659048999885822e-22

R23_70 V23 V70 41704.45859924731
L23_70 V23 V70 -5.938452422902299e-12
C23_70 V23 V70 -7.427196011280944e-21

R23_71 V23 V71 -76992.17889954374
L23_71 V23 V71 1.2400047258730313e-11
C23_71 V23 V71 -2.278469580594375e-21

R23_72 V23 V72 28841.44835215748
L23_72 V23 V72 -4.930239863064193e-12
C23_72 V23 V72 -4.0592366132500736e-21

R23_73 V23 V73 1214808.647095365
L23_73 V23 V73 2.3688039532410585e-11
C23_73 V23 V73 3.125448922615048e-21

R23_74 V23 V74 1269947.8618386409
L23_74 V23 V74 3.1775127667568825e-12
C23_74 V23 V74 6.210685703549825e-21

R23_75 V23 V75 -64025.53727033063
L23_75 V23 V75 1.634020419260423e-11
C23_75 V23 V75 1.134354369311718e-20

R23_76 V23 V76 -119855.18534140932
L23_76 V23 V76 -1.8130331887849202e-11
C23_76 V23 V76 2.6473045926177315e-21

R23_77 V23 V77 -283992.9142708712
L23_77 V23 V77 -1.9075960258273673e-10
C23_77 V23 V77 1.139784828422637e-21

R23_78 V23 V78 -692094.1086690107
L23_78 V23 V78 -2.9893208987729448e-12
C23_78 V23 V78 -1.9279235600764702e-20

R23_79 V23 V79 269227.84037645516
L23_79 V23 V79 4.701853768289837e-12
C23_79 V23 V79 5.645520712119158e-22

R23_80 V23 V80 269884.38487425697
L23_80 V23 V80 -4.011011954552225e-12
C23_80 V23 V80 -1.6353698662780472e-21

R23_81 V23 V81 333884.3566434437
L23_81 V23 V81 4.669671543504025e-12
C23_81 V23 V81 4.501942947874124e-21

R23_82 V23 V82 102683.61277676842
L23_82 V23 V82 8.060687761706131e-13
C23_82 V23 V82 3.22765966254964e-20

R23_83 V23 V83 294310.3639196891
L23_83 V23 V83 1.3420305301250255e-12
C23_83 V23 V83 2.1145037324927265e-20

R23_84 V23 V84 219884.41373563925
L23_84 V23 V84 5.466716102967932e-12
C23_84 V23 V84 -7.190577038326643e-22

R23_85 V23 V85 309545.1821144675
L23_85 V23 V85 -1.066590757491742e-11
C23_85 V23 V85 -9.364183386532871e-21

R23_86 V23 V86 -304709.34089049726
L23_86 V23 V86 -1.7675529951368788e-12
C23_86 V23 V86 -1.1824837598233057e-20

R23_87 V23 V87 -106360.47041633495
L23_87 V23 V87 -2.1896584626041077e-12
C23_87 V23 V87 -1.1934244475565432e-20

R23_88 V23 V88 -7183977.3985816585
L23_88 V23 V88 -5.061946146108188e-12
C23_88 V23 V88 -3.018014766580851e-21

R23_89 V23 V89 716874.4165036874
L23_89 V23 V89 8.404330615352264e-12
C23_89 V23 V89 8.262007538906671e-21

R23_90 V23 V90 -757038.5184942844
L23_90 V23 V90 -3.219680513321674e-12
C23_90 V23 V90 4.330625812688127e-21

R23_91 V23 V91 75870.22694213143
L23_91 V23 V91 7.473495163917702e-13
C23_91 V23 V91 2.980681274499887e-20

R23_92 V23 V92 771348.7862950801
L23_92 V23 V92 4.6914241341028676e-12
C23_92 V23 V92 6.331992617260831e-21

R23_93 V23 V93 89451.02628256209
L23_93 V23 V93 -1.431602817955311e-11
C23_93 V23 V93 -2.9627926826225165e-21

R23_94 V23 V94 836967.2098045953
L23_94 V23 V94 -3.2326530113424816e-12
C23_94 V23 V94 -1.0045720313819213e-20

R23_95 V23 V95 178216.95632997708
L23_95 V23 V95 1.529415084721166e-12
C23_95 V23 V95 1.6134211943612043e-20

R23_96 V23 V96 -2770733.980865808
L23_96 V23 V96 -3.7926135705082295e-12
C23_96 V23 V96 -4.125090378282261e-21

R23_97 V23 V97 245336.29963951907
L23_97 V23 V97 -1.7327226260781793e-12
C23_97 V23 V97 -6.75643004959836e-21

R23_98 V23 V98 153866.5608688212
L23_98 V23 V98 4.544094877310698e-12
C23_98 V23 V98 9.906039498856661e-21

R23_99 V23 V99 1177216.2088556876
L23_99 V23 V99 1.0908270950478474e-11
C23_99 V23 V99 -5.732549584245852e-22

R23_100 V23 V100 1920407.2645667994
L23_100 V23 V100 -1.2625165642740736e-11
C23_100 V23 V100 -1.4401451568836452e-21

R23_101 V23 V101 114326.60959827038
L23_101 V23 V101 3.0468889368573933e-12
C23_101 V23 V101 1.2889403829980152e-20

R23_102 V23 V102 213148.6813404256
L23_102 V23 V102 -4.609011815908349e-12
C23_102 V23 V102 1.6395659578935247e-20

R23_103 V23 V103 266126.88127162243
L23_103 V23 V103 3.2006471436670205e-12
C23_103 V23 V103 -7.100134301093077e-22

R23_104 V23 V104 -335574.0632082344
L23_104 V23 V104 -2.108548668810302e-12
C23_104 V23 V104 -5.767692525719982e-21

R23_105 V23 V105 -100355.97738892368
L23_105 V23 V105 -2.2839544677778662e-12
C23_105 V23 V105 -1.919069394590127e-20

R23_106 V23 V106 112313.40893309872
L23_106 V23 V106 9.366704261214076e-13
C23_106 V23 V106 3.0441445664034756e-20

R23_107 V23 V107 209463.12126073788
L23_107 V23 V107 -6.523910451454769e-12
C23_107 V23 V107 9.734847231436488e-21

R23_108 V23 V108 -206423.61558845287
L23_108 V23 V108 5.436034463832841e-12
C23_108 V23 V108 -8.472045414011857e-21

R23_109 V23 V109 -213737.2857747208
L23_109 V23 V109 -6.488794821258331e-12
C23_109 V23 V109 -7.650739433974754e-21

R23_110 V23 V110 -78617.67142421968
L23_110 V23 V110 -1.0440551846046014e-12
C23_110 V23 V110 -3.119364620325664e-20

R23_111 V23 V111 -217173.57831182567
L23_111 V23 V111 -9.734985287328888e-12
C23_111 V23 V111 -8.01722711946106e-21

R23_112 V23 V112 -403223.49220227473
L23_112 V23 V112 -2.7946619287373635e-11
C23_112 V23 V112 8.884958867457441e-21

R23_113 V23 V113 -890822.4042796826
L23_113 V23 V113 6.8818135842133976e-12
C23_113 V23 V113 8.342906758660634e-21

R23_114 V23 V114 90588.02662776141
L23_114 V23 V114 2.3729060981485214e-12
C23_114 V23 V114 1.4117534141947698e-20

R23_115 V23 V115 495306.0690087795
L23_115 V23 V115 -2.1178741879685387e-11
C23_115 V23 V115 4.3010619224901175e-21

R23_116 V23 V116 1152602.2756411142
L23_116 V23 V116 1.8165730366321772e-11
C23_116 V23 V116 -8.211942381506992e-21

R23_117 V23 V117 543687.7600359787
L23_117 V23 V117 -8.66686431718197e-12
C23_117 V23 V117 -1.0998859383376217e-20

R23_118 V23 V118 -106281.55186474427
L23_118 V23 V118 -1.932480862458353e-12
C23_118 V23 V118 -1.540232838752031e-20

R23_119 V23 V119 -75545.89453536716
L23_119 V23 V119 -2.1754986868740596e-12
C23_119 V23 V119 -1.4579170406310025e-20

R23_120 V23 V120 135615.79398044012
L23_120 V23 V120 -1.1620456236929334e-11
C23_120 V23 V120 1.1077754766533631e-21

R23_121 V23 V121 -131615.20035748303
L23_121 V23 V121 3.833321876075447e-11
C23_121 V23 V121 7.070135782882761e-21

R23_122 V23 V122 -101636.99774908127
L23_122 V23 V122 -2.8848257509919433e-12
C23_122 V23 V122 -1.4074084283741357e-21

R23_123 V23 V123 256632.29620599424
L23_123 V23 V123 -4.752449637029998e-12
C23_123 V23 V123 -4.028091003131042e-21

R23_124 V23 V124 2197523.173752139
L23_124 V23 V124 -1.9243567197283972e-11
C23_124 V23 V124 -5.240826075957796e-22

R23_125 V23 V125 90518.04442568697
L23_125 V23 V125 7.111925714034216e-11
C23_125 V23 V125 -3.651058598453357e-21

R23_126 V23 V126 145992.47614972384
L23_126 V23 V126 2.5707887636187116e-12
C23_126 V23 V126 8.663617196947862e-22

R23_127 V23 V127 -2365560.7575792763
L23_127 V23 V127 -6.9322252182220206e-12
C23_127 V23 V127 4.764688170749971e-22

R23_128 V23 V128 1504951.567742802
L23_128 V23 V128 4.0861042771543484e-11
C23_128 V23 V128 -4.0592417836167585e-21

R23_129 V23 V129 199219.74832283647
L23_129 V23 V129 -9.390178945169547e-12
C23_129 V23 V129 -3.0418453298713825e-21

R23_130 V23 V130 -135827.57419067482
L23_130 V23 V130 3.8501788618277794e-12
C23_130 V23 V130 -2.964112318546961e-21

R23_131 V23 V131 -781926.6822583809
L23_131 V23 V131 7.912792800652805e-12
C23_131 V23 V131 3.922401653856338e-21

R23_132 V23 V132 1259697.4434270284
L23_132 V23 V132 4.486001732708295e-12
C23_132 V23 V132 -5.440520734678208e-22

R23_133 V23 V133 289418.2798078943
L23_133 V23 V133 2.1520429705797915e-12
C23_133 V23 V133 5.3061837200469376e-21

R23_134 V23 V134 -169965.73137433792
L23_134 V23 V134 1.1080733173263909e-11
C23_134 V23 V134 1.233445807316123e-21

R23_135 V23 V135 -1360139.4309773576
L23_135 V23 V135 -6.355139379168019e-12
C23_135 V23 V135 -5.0845704819446305e-22

R23_136 V23 V136 2892570.4156034575
L23_136 V23 V136 -2.1943345574177298e-11
C23_136 V23 V136 2.997559091366626e-21

R23_137 V23 V137 152439.63234747454
L23_137 V23 V137 -1.5040473005591853e-11
C23_137 V23 V137 -1.5049387585958793e-22

R23_138 V23 V138 599628.9432155536
L23_138 V23 V138 1.99703261312263e-12
C23_138 V23 V138 -4.371602178120049e-22

R23_139 V23 V139 232619.45603224507
L23_139 V23 V139 -4.150303486128436e-12
C23_139 V23 V139 6.582501094032725e-22

R23_140 V23 V140 -339328.27850091795
L23_140 V23 V140 7.913138588839783e-12
C23_140 V23 V140 1.7504746443835383e-21

R23_141 V23 V141 217329.02426347768
L23_141 V23 V141 1.645798336364953e-11
C23_141 V23 V141 9.495460916579352e-22

R23_142 V23 V142 -115276.71263054843
L23_142 V23 V142 6.386873380427422e-12
C23_142 V23 V142 -6.988826974712063e-21

R23_143 V23 V143 -381790.54919983994
L23_143 V23 V143 7.373951422873328e-12
C23_143 V23 V143 -3.027578052965858e-21

R23_144 V23 V144 -484871.78866520646
L23_144 V23 V144 -1.245780074783596e-11
C23_144 V23 V144 -3.808346593385866e-22

R24_24 V24 0 -82077.1080317995
L24_24 V24 0 9.664401567418853e-13
C24_24 V24 0 -8.381728125724595e-20

R24_25 V24 V25 233906.72526785295
L24_25 V24 V25 3.0314640732911594e-11
C24_25 V24 V25 2.7246499711259738e-21

R24_26 V24 V26 311301.3641051659
L24_26 V24 V26 8.015460219411155e-12
C24_26 V24 V26 8.083458648732317e-22

R24_27 V24 V27 496336.2053439099
L24_27 V24 V27 1.5224851131058954e-11
C24_27 V24 V27 1.1727697423064325e-21

R24_28 V24 V28 -54278.14780208325
L24_28 V24 V28 -3.2727677805573167e-12
C24_28 V24 V28 -5.379462158448864e-21

R24_29 V24 V29 -237764.98278398404
L24_29 V24 V29 9.460774334312426e-12
C24_29 V24 V29 -1.2272096290310615e-21

R24_30 V24 V30 -492676.1416734716
L24_30 V24 V30 8.66797113279946e-12
C24_30 V24 V30 -8.426543329204946e-22

R24_31 V24 V31 24496212.660995513
L24_31 V24 V31 2.2135695011076e-11
C24_31 V24 V31 7.451596665099327e-22

R24_32 V24 V32 74291.21253362056
L24_32 V24 V32 -3.4249999088579007e-12
C24_32 V24 V32 4.983753153941554e-21

R24_33 V24 V33 2546626.696791408
L24_33 V24 V33 -1.5955549875023888e-11
C24_33 V24 V33 7.960279541997537e-22

R24_34 V24 V34 742422.6139771778
L24_34 V24 V34 4.5735385383570804e-11
C24_34 V24 V34 -3.262221336361905e-23

R24_35 V24 V35 235927.2187046816
L24_35 V24 V35 -7.086349481995106e-12
C24_35 V24 V35 2.0170863419586283e-21

R24_36 V24 V36 -375296.39623036864
L24_36 V24 V36 7.269148010366094e-12
C24_36 V24 V36 2.259971693651423e-21

R24_37 V24 V37 -302950.5709544089
L24_37 V24 V37 8.985403092856273e-12
C24_37 V24 V37 -6.378546172954407e-21

R24_38 V24 V38 -1471801.3279733986
L24_38 V24 V38 1.5009478238822734e-11
C24_38 V24 V38 -3.252929944788351e-21

R24_39 V24 V39 -240428.7119294559
L24_39 V24 V39 8.393611664246375e-12
C24_39 V24 V39 -6.542554603369454e-21

R24_40 V24 V40 -75655.07479457239
L24_40 V24 V40 -2.3663525860217856e-12
C24_40 V24 V40 9.467467727350559e-21

R24_41 V24 V41 111864.29935024198
L24_41 V24 V41 -5.356468192734708e-12
C24_41 V24 V41 1.2734441813907624e-20

R24_42 V24 V42 58291.194775509895
L24_42 V24 V42 -2.7412986454836682e-12
C24_42 V24 V42 2.008621201275746e-20

R24_43 V24 V43 3505607.835928999
L24_43 V24 V43 -9.259435464342078e-12
C24_43 V24 V43 6.344355852053417e-21

R24_44 V24 V44 -139311.1172846114
L24_44 V24 V44 1.378960858900782e-12
C24_44 V24 V44 -3.2848479952285966e-20

R24_45 V24 V45 -106104.48463369584
L24_45 V24 V45 -2.0658822089782686e-11
C24_45 V24 V45 -4.505553179444055e-21

R24_46 V24 V46 289318.52900107054
L24_46 V24 V46 4.331198834387242e-12
C24_46 V24 V46 -1.0180931506978394e-20

R24_47 V24 V47 -421652.66149094753
L24_47 V24 V47 3.691301755722586e-11
C24_47 V24 V47 -1.1824611461754424e-21

R24_48 V24 V48 77407.5582294472
L24_48 V24 V48 5.4890020468404836e-12
C24_48 V24 V48 1.7842526913478235e-20

R24_49 V24 V49 -141910.99282841376
L24_49 V24 V49 -1.6045851687747085e-11
C24_49 V24 V49 -1.0187423706398122e-21

R24_50 V24 V50 104375.14696984997
L24_50 V24 V50 -3.8486104416041366e-11
C24_50 V24 V50 5.7970494591353275e-21

R24_51 V24 V51 -346666.3390327277
L24_51 V24 V51 7.816225443934503e-12
C24_51 V24 V51 -7.641400358719285e-21

R24_52 V24 V52 -85071075.5021207
L24_52 V24 V52 -2.018264605228595e-11
C24_52 V24 V52 9.726556773662278e-21

R24_53 V24 V53 101864.11264181195
L24_53 V24 V53 -1.4589967234866783e-11
C24_53 V24 V53 9.227333645747318e-21

R24_54 V24 V54 363152.02553727356
L24_54 V24 V54 -1.4156283322547888e-11
C24_54 V24 V54 6.155654745143654e-21

R24_55 V24 V55 621179.8656627882
L24_55 V24 V55 -6.369664331157268e-11
C24_55 V24 V55 3.746073892273583e-21

R24_56 V24 V56 -27828.434492264285
L24_56 V24 V56 1.462942429485129e-11
C24_56 V24 V56 -3.583909362671213e-21

R24_57 V24 V57 96392.86459811305
L24_57 V24 V57 -3.2930078712027235e-12
C24_57 V24 V57 -4.125303635337079e-21

R24_58 V24 V58 95252.54066655107
L24_58 V24 V58 -2.923258230853315e-12
C24_58 V24 V58 6.839166735566248e-22

R24_59 V24 V59 1004301.4865502607
L24_59 V24 V59 -1.4641354503602343e-11
C24_59 V24 V59 -2.4738498112961415e-22

R24_60 V24 V60 -65826.21715346834
L24_60 V24 V60 1.8215893828542735e-12
C24_60 V24 V60 -3.671860551190213e-21

R24_61 V24 V61 -257948.26897523346
L24_61 V24 V61 -2.41476571676351e-11
C24_61 V24 V61 1.0833284393342828e-20

R24_62 V24 V62 -176486.61200869153
L24_62 V24 V62 1.457004629850375e-11
C24_62 V24 V62 2.0553980874699306e-21

R24_63 V24 V63 398446.30360501586
L24_63 V24 V63 1.110412027638037e-11
C24_63 V24 V63 -7.624934116971932e-21

R24_64 V24 V64 56688.22466624142
L24_64 V24 V64 -1.864967004883008e-11
C24_64 V24 V64 -3.964666461262333e-21

R24_65 V24 V65 -13079480.454957522
L24_65 V24 V65 -6.409701032318738e-12
C24_65 V24 V65 1.188201482693383e-21

R24_66 V24 V66 87809.33827869991
L24_66 V24 V66 -3.7308516296550996e-12
C24_66 V24 V66 6.48702805658251e-21

R24_67 V24 V67 430051.2994902617
L24_67 V24 V67 1.9220279364965746e-11
C24_67 V24 V67 -3.99400619962398e-21

R24_68 V24 V68 -53846.98814731855
L24_68 V24 V68 4.670843750794154e-12
C24_68 V24 V68 9.845796999709442e-21

R24_69 V24 V69 104012.91461637281
L24_69 V24 V69 -1.179746191168347e-11
C24_69 V24 V69 -1.2346643913181819e-21

R24_70 V24 V70 -210041.43622039072
L24_70 V24 V70 -8.501340592227788e-12
C24_70 V24 V70 1.393544068600246e-20

R24_71 V24 V71 -1008921.0063115981
L24_71 V24 V71 4.627018096623635e-11
C24_71 V24 V71 -2.661082203891299e-21

R24_72 V24 V72 262262.43520542793
L24_72 V24 V72 5.374214163953022e-11
C24_72 V24 V72 4.723585805307244e-21

R24_73 V24 V73 -125931.71259486835
L24_73 V24 V73 -6.60755024895895e-12
C24_73 V24 V73 7.951504598279781e-21

R24_74 V24 V74 -3171025.1513910135
L24_74 V24 V74 3.093689286528103e-11
C24_74 V24 V74 7.498366788822266e-21

R24_75 V24 V75 290576.5054238721
L24_75 V24 V75 9.41794347473354e-11
C24_75 V24 V75 7.22647388815279e-22

R24_76 V24 V76 105884.81328332833
L24_76 V24 V76 -9.5642973105972e-12
C24_76 V24 V76 9.695464185644896e-21

R24_77 V24 V77 -95352.87993515763
L24_77 V24 V77 4.748868634808058e-12
C24_77 V24 V77 -8.290944217857934e-21

R24_78 V24 V78 203374.73793767852
L24_78 V24 V78 -2.3889553948004983e-11
C24_78 V24 V78 1.438359122642978e-22

R24_79 V24 V79 572223.1612954834
L24_79 V24 V79 -1.411267620170764e-10
C24_79 V24 V79 6.522286762922903e-21

R24_80 V24 V80 -83101.09133847417
L24_80 V24 V80 2.993347891642766e-12
C24_80 V24 V80 -3.8277315604068943e-20

R24_81 V24 V81 36278.80939408339
L24_81 V24 V81 -1.1650191821567492e-12
C24_81 V24 V81 7.141970640690774e-20

R24_82 V24 V82 -286365.3652510456
L24_82 V24 V82 8.567633367003702e-12
C24_82 V24 V82 -1.888107847665768e-20

R24_83 V24 V83 -71025.83956201034
L24_83 V24 V83 2.6156753962216847e-12
C24_83 V24 V83 -4.4119287938766146e-20

R24_84 V24 V84 -676100.7943902733
L24_84 V24 V84 7.175135409758028e-12
C24_84 V24 V84 -5.619103156131712e-21

R24_85 V24 V85 1335070.5406954593
L24_85 V24 V85 -8.941234839352663e-12
C24_85 V24 V85 7.212299175302727e-21

R24_86 V24 V86 -188496.68214458696
L24_86 V24 V86 -1.8898215088167302e-11
C24_86 V24 V86 -6.680535076487965e-21

R24_87 V24 V87 108698.4142140542
L24_87 V24 V87 -6.9681068023596366e-12
C24_87 V24 V87 2.327626416379158e-20

R24_88 V24 V88 112339.32195225307
L24_88 V24 V88 -4.957928944495868e-12
C24_88 V24 V88 2.0097137945883893e-20

R24_89 V24 V89 -343995.1906492538
L24_89 V24 V89 1.218339641162789e-11
C24_89 V24 V89 -1.3792992903734626e-20

R24_90 V24 V90 2040141.2722467608
L24_90 V24 V90 -7.753719381023479e-12
C24_90 V24 V90 2.760700930728941e-21

R24_91 V24 V91 1833027.103112567
L24_91 V24 V91 -8.912675185446241e-12
C24_91 V24 V91 4.995706590784301e-21

R24_92 V24 V92 -41853.307856904685
L24_92 V24 V92 1.4604477379181321e-12
C24_92 V24 V92 -7.939009668970362e-20

R24_93 V24 V93 671453.0571397784
L24_93 V24 V93 -1.655737022985086e-11
C24_93 V24 V93 7.656911530937254e-21

R24_94 V24 V94 109135.0469257851
L24_94 V24 V94 -3.354454866521137e-12
C24_94 V24 V94 3.0963665948813285e-20

R24_95 V24 V95 -8438342.01487133
L24_95 V24 V95 2.122250660612307e-11
C24_95 V24 V95 -6.690182137098196e-21

R24_96 V24 V96 -34921.637420965526
L24_96 V24 V96 1.154611709313567e-12
C24_96 V24 V96 -7.815682972995385e-20

R24_97 V24 V97 112213.98746140888
L24_97 V24 V97 -2.7172599996165397e-12
C24_97 V24 V97 2.4699731455205477e-20

R24_98 V24 V98 -154732.30040515197
L24_98 V24 V98 5.206187039916679e-12
C24_98 V24 V98 -2.852120936131419e-20

R24_99 V24 V99 520231.01449337567
L24_99 V24 V99 -2.7170859802863005e-11
C24_99 V24 V99 1.0013616543260989e-20

R24_100 V24 V100 87454.45002263799
L24_100 V24 V100 -2.925304172872901e-12
C24_100 V24 V100 2.949407783573738e-20

R24_101 V24 V101 -138500.93848254113
L24_101 V24 V101 3.95021915517988e-12
C24_101 V24 V101 -2.1210702396258748e-20

R24_102 V24 V102 2388902.416575104
L24_102 V24 V102 -6.2368453741984044e-12
C24_102 V24 V102 2.247290601682931e-21

R24_103 V24 V103 -644250.3720128324
L24_103 V24 V103 4.367325453691371e-10
C24_103 V24 V103 -2.2350714148453546e-21

R24_104 V24 V104 -56254.468308048316
L24_104 V24 V104 1.741071350983571e-12
C24_104 V24 V104 -4.7991422646228123e-20

R24_105 V24 V105 83803.31379968849
L24_105 V24 V105 -3.9317353011684e-12
C24_105 V24 V105 2.9540966381902785e-20

R24_106 V24 V106 -88636.62450509232
L24_106 V24 V106 3.9167947552662315e-12
C24_106 V24 V106 -2.828693403646469e-20

R24_107 V24 V107 1093231.980955807
L24_107 V24 V107 -1.5118857163065343e-11
C24_107 V24 V107 -5.05888088859071e-21

R24_108 V24 V108 146558.5458813278
L24_108 V24 V108 -4.099503166489982e-12
C24_108 V24 V108 3.3144821099775245e-20

R24_109 V24 V109 -73911.03629811149
L24_109 V24 V109 1.9975686738484773e-12
C24_109 V24 V109 -5.116790093933871e-20

R24_110 V24 V110 149417.98257736352
L24_110 V24 V110 -3.2941445541106003e-12
C24_110 V24 V110 2.5279115544133857e-20

R24_111 V24 V111 765037.3352155694
L24_111 V24 V111 -7.946033580636515e-12
C24_111 V24 V111 2.130617035614745e-20

R24_112 V24 V112 -482593.35855377634
L24_112 V24 V112 2.13415511959243e-11
C24_112 V24 V112 -2.3657689056503512e-20

R24_113 V24 V113 179625.32465382747
L24_113 V24 V113 -4.797967242804481e-12
C24_113 V24 V113 2.4794558206202672e-20

R24_114 V24 V114 -98938.4322410497
L24_114 V24 V114 7.312293150944142e-12
C24_114 V24 V114 -2.722902411895218e-20

R24_115 V24 V115 -491515.6537318115
L24_115 V24 V115 -1.5910843121542496e-10
C24_115 V24 V115 -7.912437556715373e-21

R24_116 V24 V116 147512.5891059537
L24_116 V24 V116 -5.9549676159713465e-12
C24_116 V24 V116 2.5432497473030526e-20

R24_117 V24 V117 -157699.59052686414
L24_117 V24 V117 8.86368047423231e-12
C24_117 V24 V117 -2.0111954067572367e-20

R24_118 V24 V118 -321525.8466651256
L24_118 V24 V118 1.1277565998550926e-11
C24_118 V24 V118 -9.692205097823765e-21

R24_119 V24 V119 63858.85016967183
L24_119 V24 V119 -3.780757455265666e-12
C24_119 V24 V119 4.7695010477881526e-20

R24_120 V24 V120 127413.7841958899
L24_120 V24 V120 -3.939268195006186e-12
C24_120 V24 V120 2.9498940637822746e-20

R24_121 V24 V121 491169.43147490703
L24_121 V24 V121 -1.1521709266619532e-11
C24_121 V24 V121 3.0714479976705898e-21

R24_122 V24 V122 954326.5379076169
L24_122 V24 V122 -3.923005666079068e-12
C24_122 V24 V122 1.0575146196379053e-21

R24_123 V24 V123 -132827.46090941402
L24_123 V24 V123 -1.1731313992922055e-11
C24_123 V24 V123 3.038957937079876e-21

R24_124 V24 V124 -625756.0292892327
L24_124 V24 V124 -5.958902663154106e-12
C24_124 V24 V124 3.208031610057931e-20

R24_125 V24 V125 -319984.24852255336
L24_125 V24 V125 5.939988672984398e-11
C24_125 V24 V125 1.0368264978689686e-21

R24_126 V24 V126 -341373.29499433155
L24_126 V24 V126 3.3778473062877062e-12
C24_126 V24 V126 4.945497726893298e-22

R24_127 V24 V127 250460.38222604612
L24_127 V24 V127 -5.065478850949595e-12
C24_127 V24 V127 9.153341276412353e-21

R24_128 V24 V128 122996.53231730833
L24_128 V24 V128 1.5401907669514322e-11
C24_128 V24 V128 -9.520954283150627e-21

R24_129 V24 V129 -96889.5947338059
L24_129 V24 V129 -6.521818407044789e-12
C24_129 V24 V129 4.861676694009184e-21

R24_130 V24 V130 79801.42318894196
L24_130 V24 V130 5.29472561158804e-12
C24_130 V24 V130 -8.762177894765319e-21

R24_131 V24 V131 97697.49417420819
L24_131 V24 V131 6.7005116906978005e-12
C24_131 V24 V131 -7.40899852060429e-21

R24_132 V24 V132 124009.40340308336
L24_132 V24 V132 -1.0523274159366115e-11
C24_132 V24 V132 1.0100543736227271e-20

R24_133 V24 V133 -376357.4985791952
L24_133 V24 V133 8.870125576663093e-12
C24_133 V24 V133 -5.91345186220957e-21

R24_134 V24 V134 1505737.7346187027
L24_134 V24 V134 1.5382900434007822e-11
C24_134 V24 V134 2.5978728512601297e-21

R24_135 V24 V135 426821.29820236727
L24_135 V24 V135 -7.477701989903523e-12
C24_135 V24 V135 1.7441445218060565e-21

R24_136 V24 V136 -450193.002858054
L24_136 V24 V136 3.575310842031187e-11
C24_136 V24 V136 1.2235009882971714e-20

R24_137 V24 V137 9503800.423573809
L24_137 V24 V137 -1.7336031489384723e-10
C24_137 V24 V137 1.14665793044903e-20

R24_138 V24 V138 200405.911856482
L24_138 V24 V138 3.5740098333101823e-12
C24_138 V24 V138 1.7279123269507803e-20

R24_139 V24 V139 428277.1883551035
L24_139 V24 V139 -4.065252133806084e-12
C24_139 V24 V139 2.784780817434411e-21

R24_140 V24 V140 204084.63375370592
L24_140 V24 V140 1.2063573582120066e-11
C24_140 V24 V140 6.2172946056015716e-21

R24_141 V24 V141 -71003.6728371452
L24_141 V24 V141 7.633297758820222e-11
C24_141 V24 V141 8.410768043590923e-21

R24_142 V24 V142 69258.16450439648
L24_142 V24 V142 6.278917784165947e-12
C24_142 V24 V142 8.08866308992153e-21

R24_143 V24 V143 228326.51413972725
L24_143 V24 V143 1.0525745376151869e-11
C24_143 V24 V143 7.8176158144707705e-22

R24_144 V24 V144 751103.1755145285
L24_144 V24 V144 1.2150162156458597e-11
C24_144 V24 V144 -5.330865180602668e-21

R25_25 V25 0 693.9714618490914
L25_25 V25 0 -6.968170041079715e-13
C25_25 V25 0 8.69964729382038e-19

R25_26 V25 V26 70341.56638051482
L25_26 V25 V26 2.1147085274462356e-11
C25_26 V25 V26 -3.1429243060217433e-21

R25_27 V25 V27 72403.83160978109
L25_27 V25 V27 2.316568447536647e-11
C25_27 V25 V27 4.008105433888347e-22

R25_28 V25 V28 178484.64821658732
L25_28 V25 V28 2.2577964177263486e-11
C25_28 V25 V28 2.9108045746058764e-22

R25_29 V25 V29 -117181.1470394602
L25_29 V25 V29 -2.586952550441897e-12
C25_29 V25 V29 6.391283787705923e-20

R25_30 V25 V30 -46772.39635748962
L25_30 V25 V30 -5.364351474480467e-11
C25_30 V25 V30 -2.152611483474041e-21

R25_31 V25 V31 89735.97427058152
L25_31 V25 V31 2.077013429077073e-09
C25_31 V25 V31 4.526714703806555e-21

R25_32 V25 V32 -77228.97487599433
L25_32 V25 V32 -3.7606191159876776e-11
C25_32 V25 V32 -2.2165036923430634e-21

R25_33 V25 V33 -8569.756839106425
L25_33 V25 V33 5.693819208245239e-12
C25_33 V25 V33 -3.0261990217495246e-20

R25_34 V25 V34 22739.270752365963
L25_34 V25 V34 -1.7610289949695974e-11
C25_34 V25 V34 4.602672972730801e-21

R25_35 V25 V35 -23687.980879222978
L25_35 V25 V35 1.2714953752783497e-11
C25_35 V25 V35 3.257549990940308e-21

R25_36 V25 V36 34303.4463046225
L25_36 V25 V36 -1.1457626474842773e-10
C25_36 V25 V36 -2.0514051697819056e-22

R25_37 V25 V37 14929.055926788687
L25_37 V25 V37 -1.5816392056892553e-11
C25_37 V25 V37 1.3351905808098616e-19

R25_38 V25 V38 133088.70726174777
L25_38 V25 V38 2.2710960830411422e-11
C25_38 V25 V38 9.603616160812854e-21

R25_39 V25 V39 12530.280911862192
L25_39 V25 V39 -1.518594827120718e-11
C25_39 V25 V39 7.781218568727807e-20

R25_40 V25 V40 165863.58294371158
L25_40 V25 V40 4.34772239232048e-11
C25_40 V25 V40 6.774471884906909e-21

R25_41 V25 V41 -3103.6359608698376
L25_41 V25 V41 2.2684624458762e-12
C25_41 V25 V41 -4.0857817029150847e-19

R25_42 V25 V42 -4955.177673781552
L25_42 V25 V42 3.4395039697768527e-12
C25_42 V25 V42 -2.8376559465745705e-19

R25_43 V25 V43 -9539.23768209142
L25_43 V25 V43 5.784273224010596e-12
C25_43 V25 V43 -1.247445084716319e-19

R25_44 V25 V44 -119669.02024476646
L25_44 V25 V44 9.111536085538239e-11
C25_44 V25 V44 -6.6362426598076215e-21

R25_45 V25 V45 188394.9604124238
L25_45 V25 V45 -1.354547183898553e-11
C25_45 V25 V45 2.8905973230998344e-19

R25_46 V25 V46 -51244.49985059829
L25_46 V25 V46 -1.414707983958181e-11
C25_46 V25 V46 1.5520123266615426e-19

R25_47 V25 V47 -25817.641691566085
L25_47 V25 V47 -3.093969401963609e-11
C25_47 V25 V47 4.066257355061725e-20

R25_48 V25 V48 42398.37046889063
L25_48 V25 V48 -4.133904433967371e-11
C25_48 V25 V48 8.35379602892225e-21

R25_49 V25 V49 -52955.33847846544
L25_49 V25 V49 1.1845101585548993e-11
C25_49 V25 V49 -6.79394336242923e-20

R25_50 V25 V50 -17349.573355685076
L25_50 V25 V50 9.641740956800173e-12
C25_50 V25 V50 -6.524364596504535e-20

R25_51 V25 V51 17390.816244314145
L25_51 V25 V51 -1.2300277388811036e-11
C25_51 V25 V51 5.512920776715295e-20

R25_52 V25 V52 -10480.21423638014
L25_52 V25 V52 4.2158011928296016e-12
C25_52 V25 V52 -1.8560390263172108e-19

R25_53 V25 V53 -12618.970335778302
L25_53 V25 V53 3.979381629623927e-12
C25_53 V25 V53 -9.994015972945462e-20

R25_54 V25 V54 -16446.000533134087
L25_54 V25 V54 1.5429108243816918e-11
C25_54 V25 V54 -2.1085973856796352e-20

R25_55 V25 V55 -11628.471126618379
L25_55 V25 V55 1.0450897031973934e-11
C25_55 V25 V55 -5.414896859744795e-20

R25_56 V25 V56 -17688.231379853692
L25_56 V25 V56 1.5403130064772152e-11
C25_56 V25 V56 -5.626467584858002e-20

R25_57 V25 V57 -2043.4245759869825
L25_57 V25 V57 3.0991631244763144e-12
C25_57 V25 V57 2.9021342856454605e-20

R25_58 V25 V58 -15416.738934517538
L25_58 V25 V58 2.0284399304989776e-11
C25_58 V25 V58 1.6125966650305237e-20

R25_59 V25 V59 63679.52164619651
L25_59 V25 V59 -2.730723566347626e-11
C25_59 V25 V59 2.2381495704617398e-20

R25_60 V25 V60 -37286.333126092955
L25_60 V25 V60 3.3869051599496625e-11
C25_60 V25 V60 7.421686671484097e-21

R25_61 V25 V61 16664.319097333148
L25_61 V25 V61 1.6892116463340912e-11
C25_61 V25 V61 -1.1805100470500173e-19

R25_62 V25 V62 10677.050803981592
L25_62 V25 V62 -5.0628891761284985e-11
C25_62 V25 V62 -9.407494502751392e-20

R25_63 V25 V63 19858.199657547884
L25_63 V25 V63 -3.1119160022787764e-11
C25_63 V25 V63 -2.51176110616755e-20

R25_64 V25 V64 -54490.345100735925
L25_64 V25 V64 2.1474155750454233e-11
C25_64 V25 V64 -2.0718300632075042e-20

R25_65 V25 V65 -3710.7486044769153
L25_65 V25 V65 3.281568819285143e-12
C25_65 V25 V65 -3.237098914253013e-20

R25_66 V25 V66 -3873.5259643461095
L25_66 V25 V66 2.6083543182034664e-12
C25_66 V25 V66 -2.8396432825101206e-20

R25_67 V25 V67 -11320.202498765193
L25_67 V25 V67 5.827678157764318e-11
C25_67 V25 V67 -2.113255807344695e-20

R25_68 V25 V68 -125996.8391102212
L25_68 V25 V68 -3.7269878391333136e-10
C25_68 V25 V68 -1.3533576126685643e-20

R25_69 V25 V69 267703.67311904475
L25_69 V25 V69 -9.113642640231318e-12
C25_69 V25 V69 7.44905152566905e-21

R25_70 V25 V70 11230.849920066094
L25_70 V25 V70 -2.2771076920311427e-11
C25_70 V25 V70 -3.0007713649582234e-20

R25_71 V25 V71 15853.24109268416
L25_71 V25 V71 -8.561925568343089e-11
C25_71 V25 V71 -9.35344872672754e-21

R25_72 V25 V72 11781.554970034615
L25_72 V25 V72 -6.151443474160073e-12
C25_72 V25 V72 -1.3884503511289797e-20

R25_73 V25 V73 184295.091145965
L25_73 V25 V73 -1.1487477506866294e-11
C25_73 V25 V73 -2.4764614763446414e-20

R25_74 V25 V74 24196.413150931097
L25_74 V25 V74 -1.0372103282793641e-11
C25_74 V25 V74 1.5775974647830636e-20

R25_75 V25 V75 -14257.809652311753
L25_75 V25 V75 4.0531660941583326e-11
C25_75 V25 V75 -4.749860275062913e-21

R25_76 V25 V76 -13506.775872312734
L25_76 V25 V76 7.933756519861756e-12
C25_76 V25 V76 -2.4753775092145273e-20

R25_77 V25 V77 -41287.88558883284
L25_77 V25 V77 1.6442010778590302e-11
C25_77 V25 V77 2.367012405113191e-21

R25_78 V25 V78 -53681.05701400941
L25_78 V25 V78 1.6159438643974835e-11
C25_78 V25 V78 -2.0428631146362375e-20

R25_79 V25 V79 57230.189641640354
L25_79 V25 V79 1.868068961302237e-11
C25_79 V25 V79 -5.069767936495985e-21

R25_80 V25 V80 32729.786104207287
L25_80 V25 V80 4.8883706011761995e-11
C25_80 V25 V80 1.9375504944332132e-20

R25_81 V25 V81 84796.99188655018
L25_81 V25 V81 -1.8626764862534087e-11
C25_81 V25 V81 -1.75667459346331e-20

R25_82 V25 V82 525305.1898753139
L25_82 V25 V82 7.296008000747663e-11
C25_82 V25 V82 4.647116948599379e-20

R25_83 V25 V83 35367.8943935231
L25_83 V25 V83 -5.500207757168381e-12
C25_83 V25 V83 2.3011389313239244e-20

R25_84 V25 V84 241246.8982434121
L25_84 V25 V84 -5.3842946086052965e-12
C25_84 V25 V84 -1.1911029943616026e-20

R25_85 V25 V85 48615.312638874406
L25_85 V25 V85 -1.036671600896051e-11
C25_85 V25 V85 -2.4633864127444816e-20

R25_86 V25 V86 -312523.30125166697
L25_86 V25 V86 -3.3371888447491646e-11
C25_86 V25 V86 -1.4911310009485128e-20

R25_87 V25 V87 -55028.61159520394
L25_87 V25 V87 -1.0922564295074963e-10
C25_87 V25 V87 -2.819086406070282e-20

R25_88 V25 V88 -97342.40766038487
L25_88 V25 V88 3.9430365491534143e-11
C25_88 V25 V88 -9.204682580138883e-21

R25_89 V25 V89 -167640.1670259223
L25_89 V25 V89 3.531515777890666e-12
C25_89 V25 V89 3.014797572986978e-20

R25_90 V25 V90 87068.1658701582
L25_90 V25 V90 1.5476545671403778e-10
C25_90 V25 V90 4.64029440471523e-21

R25_91 V25 V91 51650.611984461895
L25_91 V25 V91 -1.1964470166391831e-11
C25_91 V25 V91 3.068750222987771e-20

R25_92 V25 V92 101312.29123728398
L25_92 V25 V92 -3.4291339842701044e-11
C25_92 V25 V92 2.6732793279623845e-20

R25_93 V25 V93 26031.51899123096
L25_93 V25 V93 2.920900578337252e-11
C25_93 V25 V93 4.661876680253972e-21

R25_94 V25 V94 -170663.1324170923
L25_94 V25 V94 -1.502767549225312e-11
C25_94 V25 V94 -2.037405242538008e-20

R25_95 V25 V95 89593.17704067177
L25_95 V25 V95 -1.4065348283597817e-11
C25_95 V25 V95 2.1495203214489537e-20

R25_96 V25 V96 1368878.682913289
L25_96 V25 V96 -1.8064847257414193e-11
C25_96 V25 V96 2.262031262513962e-20

R25_97 V25 V97 47484.53893596054
L25_97 V25 V97 7.0762437576319136e-12
C25_97 V25 V97 -7.265270578986602e-21

R25_98 V25 V98 23892.779910250116
L25_98 V25 V98 5.854267510460873e-12
C25_98 V25 V98 2.3523383333813404e-20

R25_99 V25 V99 -172902.28103882313
L25_99 V25 V99 2.1323497548685573e-11
C25_99 V25 V99 -3.703624416164727e-21

R25_100 V25 V100 -95137.11501301886
L25_100 V25 V100 2.4428135210293147e-10
C25_100 V25 V100 -9.385870264627789e-21

R25_101 V25 V101 44132.6498728003
L25_101 V25 V101 4.3154712285402925e-12
C25_101 V25 V101 3.139653012188466e-20

R25_102 V25 V102 44493.04109575174
L25_102 V25 V102 2.118837073859051e-11
C25_102 V25 V102 1.8543567965187374e-20

R25_103 V25 V103 182199.32315415452
L25_103 V25 V103 8.271909277297614e-12
C25_103 V25 V103 -6.6784644986936325e-21

R25_104 V25 V104 -502902.7427921176
L25_104 V25 V104 3.270286886032748e-10
C25_104 V25 V104 1.039404931923973e-20

R25_105 V25 V105 -41311.45099040617
L25_105 V25 V105 2.0806435265736374e-11
C25_105 V25 V105 -2.222915741256384e-20

R25_106 V25 V106 -201579.79895203846
L25_106 V25 V106 -4.6799336641412115e-12
C25_106 V25 V106 4.680216538237431e-20

R25_107 V25 V107 139937.77201749486
L25_107 V25 V107 -9.652686676217096e-12
C25_107 V25 V107 1.0778507719180584e-20

R25_108 V25 V108 1108327.1613781673
L25_108 V25 V108 -1.8905628579409057e-11
C25_108 V25 V108 -2.6065377743855318e-20

R25_109 V25 V109 140643.85893635202
L25_109 V25 V109 2.6822830502761668e-11
C25_109 V25 V109 3.42073792805423e-21

R25_110 V25 V110 932912.2332469322
L25_110 V25 V110 -3.62171808565008e-11
C25_110 V25 V110 -4.499594454800222e-20

R25_111 V25 V111 -37602.27490843365
L25_111 V25 V111 5.601335461973543e-12
C25_111 V25 V111 -1.535182062035712e-20

R25_112 V25 V112 43089.44820817142
L25_112 V25 V112 4.92181103254216e-12
C25_112 V25 V112 2.5865020243387028e-20

R25_113 V25 V113 131273.64785172074
L25_113 V25 V113 1.2849695821980934e-11
C25_113 V25 V113 9.145630741174443e-21

R25_114 V25 V114 59846.949306875256
L25_114 V25 V114 -3.13614878926617e-11
C25_114 V25 V114 2.764782031452772e-20

R25_115 V25 V115 52306.93599544312
L25_115 V25 V115 -9.975281389504395e-12
C25_115 V25 V115 8.496092747939116e-21

R25_116 V25 V116 -128495.31427222001
L25_116 V25 V116 -1.1427824474642858e-11
C25_116 V25 V116 -1.6492113233616403e-20

R25_117 V25 V117 42237.810164400944
L25_117 V25 V117 -1.0716689005016168e-11
C25_117 V25 V117 -9.536062559207806e-21

R25_118 V25 V118 -34387.16646018343
L25_118 V25 V118 -2.963026997084941e-11
C25_118 V25 V118 -1.9177906892201626e-20

R25_119 V25 V119 -33932.16065552629
L25_119 V25 V119 8.813594559160727e-12
C25_119 V25 V119 -3.000211045938597e-20

R25_120 V25 V120 18284.663107744676
L25_120 V25 V120 -4.639902636333305e-12
C25_120 V25 V120 -1.3213532369082134e-20

R25_121 V25 V121 -209914.43002447413
L25_121 V25 V121 4.6772934387454486e-12
C25_121 V25 V121 -3.4031715059494415e-22

R25_122 V25 V122 13618.127494769884
L25_122 V25 V122 4.981625318831431e-12
C25_122 V25 V122 6.772973774486718e-21

R25_123 V25 V123 101504.2187474795
L25_123 V25 V123 3.4758202904864124e-11
C25_123 V25 V123 -5.163331515508264e-21

R25_124 V25 V124 -98808.30654776188
L25_124 V25 V124 1.6708313055438263e-11
C25_124 V25 V124 -1.0667632494124039e-20

R25_125 V25 V125 31393.75218410997
L25_125 V25 V125 -2.7582828016633054e-12
C25_125 V25 V125 -4.134443029716092e-21

R25_126 V25 V126 -12411.73205793612
L25_126 V25 V126 -1.6464748216526265e-10
C25_126 V25 V126 1.9726224319304924e-21

R25_127 V25 V127 12152.247280189222
L25_127 V25 V127 -1.3176640165567327e-11
C25_127 V25 V127 -1.5425552566499105e-21

R25_128 V25 V128 66549.66171657029
L25_128 V25 V128 -1.915179384164683e-10
C25_128 V25 V128 -3.2132129380557097e-21

R25_129 V25 V129 33153.17348681641
L25_129 V25 V129 -5.471228550447108e-11
C25_129 V25 V129 -3.792086097143324e-21

R25_130 V25 V130 -96980.71000795202
L25_130 V25 V130 7.086803599159191e-10
C25_130 V25 V130 -7.34104426676401e-21

R25_131 V25 V131 -86060.73077031634
L25_131 V25 V131 -1.5665066683542607e-11
C25_131 V25 V131 3.179739897733061e-21

R25_132 V25 V132 -48081.42059367125
L25_132 V25 V132 -5.887220936361432e-11
C25_132 V25 V132 -1.6145045927665001e-21

R25_133 V25 V133 -655698.3734680368
L25_133 V25 V133 -6.769199724166105e-12
C25_133 V25 V133 1.2061986956575021e-20

R25_134 V25 V134 -29463.432874862287
L25_134 V25 V134 -9.762495096363594e-12
C25_134 V25 V134 -4.876426319407489e-21

R25_135 V25 V135 24713.248354340252
L25_135 V25 V135 -1.967590815359292e-11
C25_135 V25 V135 -3.155063250210962e-21

R25_136 V25 V136 232978.64141742786
L25_136 V25 V136 -4.7643830176629825e-11
C25_136 V25 V136 -2.3390763452525474e-21

R25_137 V25 V137 102075.684067341
L25_137 V25 V137 -6.582589836880777e-12
C25_137 V25 V137 -1.461651590365114e-20

R25_138 V25 V138 -11345.287359528449
L25_138 V25 V138 -1.1433066442852e-11
C25_138 V25 V138 -1.4451919696033428e-20

R25_139 V25 V139 8340.436874609337
L25_139 V25 V139 -1.0096686148651724e-11
C25_139 V25 V139 7.738242710294774e-21

R25_140 V25 V140 -63452.22658131531
L25_140 V25 V140 1.1260286446042164e-10
C25_140 V25 V140 9.513746163749924e-21

R25_141 V25 V141 586018.0946496035
L25_141 V25 V141 4.1383052279617324e-11
C25_141 V25 V141 1.7361685739711153e-21

R25_142 V25 V142 -31920.633056605693
L25_142 V25 V142 1.6944170689107013e-10
C25_142 V25 V142 2.9213038575284417e-21

R25_143 V25 V143 -25648.586385255538
L25_143 V25 V143 5.5337306543475404e-11
C25_143 V25 V143 -7.321679212619021e-21

R25_144 V25 V144 -84329.78486342776
L25_144 V25 V144 -3.835690057375089e-11
C25_144 V25 V144 -6.893183718961952e-21

R26_26 V26 0 -1425.4935043629268
L26_26 V26 0 3.7015632448141355e-13
C26_26 V26 0 2.2469727589205623e-19

R26_27 V26 V27 -72414.13150365495
L26_27 V26 V27 -1.6257718882738278e-11
C26_27 V26 V27 5.566438578534653e-22

R26_28 V26 V28 -172319.051463464
L26_28 V26 V28 1.83522193830698e-10
C26_28 V26 V28 -1.4559930662131662e-22

R26_29 V26 V29 45825.04077089299
L26_29 V26 V29 3.8361787603786156e-11
C26_29 V26 V29 1.3106328883812495e-20

R26_30 V26 V30 -73907.34612041661
L26_30 V26 V30 -3.777223095902143e-12
C26_30 V26 V30 6.598563317694599e-21

R26_31 V26 V31 236244.78644845844
L26_31 V26 V31 6.983128749324472e-12
C26_31 V26 V31 -7.363400509193886e-21

R26_32 V26 V32 113782.03866887091
L26_32 V26 V32 1.198471416253698e-11
C26_32 V26 V32 -4.1552993918017816e-21

R26_33 V26 V33 325081.29707827896
L26_33 V26 V33 -1.6369618522427665e-11
C26_33 V26 V33 -6.611729899688395e-21

R26_34 V26 V34 376781.3168959425
L26_34 V26 V34 3.578230323357956e-11
C26_34 V26 V34 -1.4616950370853381e-21

R26_35 V26 V35 -83004.1460968339
L26_35 V26 V35 -1.5260570651338423e-11
C26_35 V26 V35 1.489931276670137e-20

R26_36 V26 V36 -131223.8984637559
L26_36 V26 V36 -5.003059422213886e-11
C26_36 V26 V36 2.7355188514716565e-22

R26_37 V26 V37 45863.5240747253
L26_37 V26 V37 6.98672777559122e-12
C26_37 V26 V37 2.460770887700276e-20

R26_38 V26 V38 81743.93302911503
L26_38 V26 V38 -8.740628682649655e-12
C26_38 V26 V38 3.506836610232829e-20

R26_39 V26 V39 -122121.21193317685
L26_39 V26 V39 9.758151092716618e-12
C26_39 V26 V39 -8.134544702292095e-21

R26_40 V26 V40 -161284.74399383666
L26_40 V26 V40 1.1590108984689094e-11
C26_40 V26 V40 -1.9069589661376878e-20

R26_41 V26 V41 19900.77085593887
L26_41 V26 V41 -2.178508521944955e-12
C26_41 V26 V41 -8.017810528515608e-20

R26_42 V26 V42 -50241.93414008257
L26_42 V26 V42 2.7570971143015515e-11
C26_42 V26 V42 -1.4485599768053808e-19

R26_43 V26 V43 67824.99698002478
L26_43 V26 V43 -1.6162554268543055e-11
C26_43 V26 V43 6.182452560941256e-20

R26_44 V26 V44 826052.4514843203
L26_44 V26 V44 -2.1303549444526267e-11
C26_44 V26 V44 2.8984020971563006e-20

R26_45 V26 V45 14809.770866483013
L26_45 V26 V45 5.2628847346167915e-12
C26_45 V26 V45 2.0109999301846346e-20

R26_46 V26 V46 10613.83088201793
L26_46 V26 V46 -9.488853790682641e-12
C26_46 V26 V46 1.2833643428930569e-19

R26_47 V26 V47 -48746.35247478487
L26_47 V26 V47 -7.080925505431903e-12
C26_47 V26 V47 -4.0139420432726215e-20

R26_48 V26 V48 -91151.73658969534
L26_48 V26 V48 -1.6249774103186882e-11
C26_48 V26 V48 -2.0202590364369193e-20

R26_49 V26 V49 95612.95160663304
L26_49 V26 V49 6.400977779190278e-11
C26_49 V26 V49 -6.60715025507494e-21

R26_50 V26 V50 -27948.72537354906
L26_50 V26 V50 5.7891215025915255e-11
C26_50 V26 V50 -2.994376826635405e-20

R26_51 V26 V51 48814.139607151934
L26_51 V26 V51 -7.444462093321405e-12
C26_51 V26 V51 4.604269664310851e-20

R26_52 V26 V52 -36592.48297883498
L26_52 V26 V52 -4.4340017441059645e-11
C26_52 V26 V52 -4.2438622245587564e-20

R26_53 V26 V53 -40521.966805888565
L26_53 V26 V53 -6.656389132593049e-12
C26_53 V26 V53 -3.5449700894762596e-20

R26_54 V26 V54 97510.30359330283
L26_54 V26 V54 -4.152507168919951e-11
C26_54 V26 V54 -3.214902831276011e-20

R26_55 V26 V55 19086.786376181302
L26_55 V26 V55 -3.485967824077301e-11
C26_55 V26 V55 2.0843289340385113e-21

R26_56 V26 V56 26686.616084170775
L26_56 V26 V56 -5.477703947776029e-12
C26_56 V26 V56 -5.2751056970401325e-21

R26_57 V26 V57 3649.9961070987706
L26_57 V26 V57 -3.2412946997428055e-12
C26_57 V26 V57 8.97619871608656e-21

R26_58 V26 V58 6230.056225229457
L26_58 V26 V58 1.724265458347673e-11
C26_58 V26 V58 -6.441981701605456e-21

R26_59 V26 V59 -37511.38668617264
L26_59 V26 V59 -1.0068330483360885e-11
C26_59 V26 V59 -7.274946401215472e-21

R26_60 V26 V60 41876.93319301652
L26_60 V26 V60 -5.844975042869707e-12
C26_60 V26 V60 1.5975963734643551e-21

R26_61 V26 V61 -10257.459970343085
L26_61 V26 V61 -1.4470592855308323e-11
C26_61 V26 V61 -3.9378178385404086e-20

R26_62 V26 V62 -7448.115523249756
L26_62 V26 V62 9.273161651153315e-12
C26_62 V26 V62 -1.5842582390910406e-20

R26_63 V26 V63 18673.703799079616
L26_63 V26 V63 -8.555775238919843e-12
C26_63 V26 V63 -1.9178026471426183e-20

R26_64 V26 V64 169029.99966611507
L26_64 V26 V64 -6.628897542802678e-12
C26_64 V26 V64 -1.4170080855089134e-20

R26_65 V26 V65 11194.884554802318
L26_65 V26 V65 -7.821604206463078e-11
C26_65 V26 V65 -8.447155123129275e-21

R26_66 V26 V66 13063.001857886997
L26_66 V26 V66 -1.8361007432770813e-11
C26_66 V26 V66 -2.137088755565738e-21

R26_67 V26 V67 224066.5994596876
L26_67 V26 V67 -6.023142975235867e-12
C26_67 V26 V67 1.063983503738355e-21

R26_68 V26 V68 70136.42576974553
L26_68 V26 V68 -1.60513043576318e-11
C26_68 V26 V68 -5.433935961371332e-21

R26_69 V26 V69 -249695.6190938341
L26_69 V26 V69 -8.457506725887022e-12
C26_69 V26 V69 -1.2255189676446686e-20

R26_70 V26 V70 -40709.32821178747
L26_70 V26 V70 -8.347924848290293e-12
C26_70 V26 V70 -1.94439061038608e-20

R26_71 V26 V71 -158647.2198208718
L26_71 V26 V71 -6.07179835897888e-11
C26_71 V26 V71 -5.682634905889796e-21

R26_72 V26 V72 -48598.95898890634
L26_72 V26 V72 -1.2331423848980425e-11
C26_72 V26 V72 -7.691710703122856e-21

R26_73 V26 V73 275350.09549049014
L26_73 V26 V73 -7.483746730836645e-12
C26_73 V26 V73 -1.2527478674021684e-20

R26_74 V26 V74 -86112.72469661341
L26_74 V26 V74 -4.5146437991102174e-12
C26_74 V26 V74 3.0427737532039243e-21

R26_75 V26 V75 56932.23332955954
L26_75 V26 V75 6.274713439348715e-12
C26_75 V26 V75 1.435738811913525e-20

R26_76 V26 V76 -179035.37077958032
L26_76 V26 V76 -3.3504482649358376e-12
C26_76 V26 V76 -1.504367748503423e-20

R26_77 V26 V77 1375328.9033484254
L26_77 V26 V77 -1.046041766948136e-11
C26_77 V26 V77 3.857585128397912e-21

R26_78 V26 V78 -76135.8406352631
L26_78 V26 V78 -1.0064072425902438e-11
C26_78 V26 V78 -1.4584474283109804e-20

R26_79 V26 V79 -66067.1464682203
L26_79 V26 V79 -2.1296753376035135e-12
C26_79 V26 V79 -2.2427760016650184e-20

R26_80 V26 V80 246438.00528092124
L26_80 V26 V80 3.941655117619601e-12
C26_80 V26 V80 2.570055556103534e-20

R26_81 V26 V81 -368184.9558668555
L26_81 V26 V81 6.329470051742189e-12
C26_81 V26 V81 -9.309052757143551e-21

R26_82 V26 V82 218733.27967679402
L26_82 V26 V82 2.945368509604755e-11
C26_82 V26 V82 2.4243519801797046e-20

R26_83 V26 V83 75202.6442912419
L26_83 V26 V83 6.014967201255399e-12
C26_83 V26 V83 2.923004568337426e-20

R26_84 V26 V84 1796675.368220225
L26_84 V26 V84 -3.3602737486665327e-12
C26_84 V26 V84 -1.6551334256009207e-20

R26_85 V26 V85 -122654.95512546918
L26_85 V26 V85 -3.117451229539628e-12
C26_85 V26 V85 -2.7746349610044295e-20

R26_86 V26 V86 -217476.6107968881
L26_86 V26 V86 -5.297572167831331e-11
C26_86 V26 V86 -8.01557279215224e-21

R26_87 V26 V87 -99018.05462267369
L26_87 V26 V87 -4.845551745828109e-12
C26_87 V26 V87 -2.140840619367085e-20

R26_88 V26 V88 -74725.42821807656
L26_88 V26 V88 1.2521493656341096e-11
C26_88 V26 V88 -3.603844273156595e-21

R26_89 V26 V89 195199.84740019747
L26_89 V26 V89 -5.3302519688379576e-11
C26_89 V26 V89 1.6769328526987534e-20

R26_90 V26 V90 61109.8559564974
L26_90 V26 V90 1.8777575904394785e-12
C26_90 V26 V90 2.946327736132583e-20

R26_91 V26 V91 109888.60241044656
L26_91 V26 V91 1.9412401674973138e-11
C26_91 V26 V91 1.9134670100296578e-20

R26_92 V26 V92 107858.58044185204
L26_92 V26 V92 -3.092579555890579e-11
C26_92 V26 V92 2.2307280883624228e-20

R26_93 V26 V93 -26702.943827907573
L26_93 V26 V93 -1.0435638438201597e-11
C26_93 V26 V93 -2.635594386946728e-21

R26_94 V26 V94 -36240.86912143541
L26_94 V26 V94 8.666841517992476e-12
C26_94 V26 V94 -8.977217610088767e-21

R26_95 V26 V95 410081.49233427166
L26_95 V26 V95 2.793926046282821e-11
C26_95 V26 V95 1.4514404436645978e-20

R26_96 V26 V96 120685.60295383658
L26_96 V26 V96 -6.476654587982621e-11
C26_96 V26 V96 2.0382146227458378e-20

R26_97 V26 V97 73167.3439843243
L26_97 V26 V97 2.8001146927114428e-12
C26_97 V26 V97 6.4686149910837165e-21

R26_98 V26 V98 30952.557243133695
L26_98 V26 V98 5.984097418576334e-12
C26_98 V26 V98 2.039160015924354e-20

R26_99 V26 V99 -46770.02413069406
L26_99 V26 V99 -4.5558210770550394e-12
C26_99 V26 V99 -7.461885086020241e-21

R26_100 V26 V100 -1132978.2005934643
L26_100 V26 V100 1.1860268750510093e-11
C26_100 V26 V100 -1.9614781723687663e-21

R26_101 V26 V101 -209797.5958285306
L26_101 V26 V101 1.8492896935123122e-08
C26_101 V26 V101 2.133738708317039e-20

R26_102 V26 V102 39525.878849280765
L26_102 V26 V102 9.86155596185971e-13
C26_102 V26 V102 5.832006618852606e-20

R26_103 V26 V103 -116976.9123293752
L26_103 V26 V103 -1.6985519511724819e-12
C26_103 V26 V103 -3.6001976746735736e-20

R26_104 V26 V104 -295483.7329846408
L26_104 V26 V104 -1.1960236101638721e-11
C26_104 V26 V104 1.3135273487233416e-20

R26_105 V26 V105 -104525.76865248439
L26_105 V26 V105 -3.3998722721798422e-12
C26_105 V26 V105 -2.8184082105454243e-20

R26_106 V26 V106 200411.30962233545
L26_106 V26 V106 2.296868132937703e-12
C26_106 V26 V106 5.126053771989225e-20

R26_107 V26 V107 55196.532766486394
L26_107 V26 V107 1.1855345703039685e-12
C26_107 V26 V107 4.83660791073232e-20

R26_108 V26 V108 90985.94941813553
L26_108 V26 V108 -1.664975169700143e-12
C26_108 V26 V108 -4.4044679647622047e-20

R26_109 V26 V109 120980.14287925976
L26_109 V26 V109 -2.4045376381191116e-12
C26_109 V26 V109 -1.1140216778148308e-20

R26_110 V26 V110 115805.29309016495
L26_110 V26 V110 -1.5664254876442056e-11
C26_110 V26 V110 -4.2008522266116e-20

R26_111 V26 V111 -252067.9125287248
L26_111 V26 V111 -2.0604718492085706e-12
C26_111 V26 V111 -2.5346364801402384e-20

R26_112 V26 V112 16192.372325471231
L26_112 V26 V112 1.7156718366515225e-12
C26_112 V26 V112 3.447822630516811e-20

R26_113 V26 V113 32374.588723800425
L26_113 V26 V113 3.2631396264867085e-12
C26_113 V26 V113 1.5191313828703682e-20

R26_114 V26 V114 68933.7526576806
L26_114 V26 V114 4.737350218442908e-12
C26_114 V26 V114 2.1242495585559234e-20

R26_115 V26 V115 70777.4546015861
L26_115 V26 V115 2.289806458725508e-12
C26_115 V26 V115 2.7433702773003847e-20

R26_116 V26 V116 -58016.84840286328
L26_116 V26 V116 -3.050853258031833e-12
C26_116 V26 V116 -2.790807767309363e-20

R26_117 V26 V117 -313173.78008562064
L26_117 V26 V117 -4.85587761665546e-12
C26_117 V26 V117 -2.1413635434896896e-20

R26_118 V26 V118 -72098.64889644651
L26_118 V26 V118 -4.683403180971883e-12
C26_118 V26 V118 -1.8173726913129513e-20

R26_119 V26 V119 1565765.4585004183
L26_119 V26 V119 -4.010353016944195e-12
C26_119 V26 V119 -2.3689454832804393e-20

R26_120 V26 V120 56674.65229950523
L26_120 V26 V120 2.4744895016232006e-12
C26_120 V26 V120 -1.277467660011264e-20

R26_121 V26 V121 16438.54924172283
L26_121 V26 V121 1.1597523032063436e-11
C26_121 V26 V121 4.089310882408204e-21

R26_122 V26 V122 7209.681255104227
L26_122 V26 V122 1.7793062786969394e-12
C26_122 V26 V122 2.368157284141401e-21

R26_123 V26 V123 44508.01178050884
L26_123 V26 V123 7.632566079186613e-12
C26_123 V26 V123 -4.361074320265356e-21

R26_124 V26 V124 470844.85507507244
L26_124 V26 V124 -2.0751674687291323e-11
C26_124 V26 V124 -9.500913559340635e-21

R26_125 V26 V125 -18845.087255038678
L26_125 V26 V125 1.1488351188241941e-11
C26_125 V26 V125 -3.944280397846982e-21

R26_126 V26 V126 -7934.800094113753
L26_126 V26 V126 -1.3786860394897319e-12
C26_126 V26 V126 7.730610739898928e-21

R26_127 V26 V127 13152.408484233723
L26_127 V26 V127 1.5955096699592168e-12
C26_127 V26 V127 -1.9866600007805365e-21

R26_128 V26 V128 -673205.1289283944
L26_128 V26 V128 3.449869909073565e-11
C26_128 V26 V128 -4.779611755518514e-21

R26_129 V26 V129 32474.136393018533
L26_129 V26 V129 4.1234519369777425e-12
C26_129 V26 V129 -7.352696569106572e-21

R26_130 V26 V130 -30090.768218967136
L26_130 V26 V130 -2.2475968157993945e-12
C26_130 V26 V130 -1.427521271223267e-20

R26_131 V26 V131 -26077.629077012563
L26_131 V26 V131 -1.4590484380385396e-10
C26_131 V26 V131 1.3389672495026533e-20

R26_132 V26 V132 -39507.020988793534
L26_132 V26 V132 -6.6272044011572725e-12
C26_132 V26 V132 -4.918785084255641e-21

R26_133 V26 V133 -70331.30089927798
L26_133 V26 V133 1.6003645030761303e-11
C26_133 V26 V133 1.0393091123330938e-20

R26_134 V26 V134 -48518.52003106018
L26_134 V26 V134 -1.4158281089234274e-11
C26_134 V26 V134 8.278384894380188e-22

R26_135 V26 V135 18127.565467447457
L26_135 V26 V135 2.6934190494818516e-12
C26_135 V26 V135 -5.1631033313384325e-21

R26_136 V26 V136 -154638.09548215743
L26_136 V26 V136 3.950638106767929e-11
C26_136 V26 V136 2.0507560388040673e-21

R26_137 V26 V137 -24515.72400271074
L26_137 V26 V137 -4.902147056065224e-11
C26_137 V26 V137 -6.569379359306489e-21

R26_138 V26 V138 -8207.075688469073
L26_138 V26 V138 -1.4016620799461762e-12
C26_138 V26 V138 -1.105091757935446e-20

R26_139 V26 V139 10044.763468355555
L26_139 V26 V139 1.1575358904017532e-12
C26_139 V26 V139 6.747441774687996e-21

R26_140 V26 V140 -33820.59212198687
L26_140 V26 V140 -3.21453402758568e-12
C26_140 V26 V140 2.9661601410089345e-21

R26_141 V26 V141 -36953.84969540879
L26_141 V26 V141 -6.119366380383264e-12
C26_141 V26 V141 -7.7748431491290465e-22

R26_142 V26 V142 -35709.02508427685
L26_142 V26 V142 -2.764418965691155e-12
C26_142 V26 V142 -5.9147819781651106e-21

R26_143 V26 V143 -33970.38960475039
L26_143 V26 V143 -3.820754916110532e-12
C26_143 V26 V143 -6.249521945728415e-21

R26_144 V26 V144 35292.38890334274
L26_144 V26 V144 7.266929732504207e-12
C26_144 V26 V144 2.2393009028478735e-21

R27_27 V27 0 -1272.1702462939081
L27_27 V27 0 1.055443470872547e-12
C27_27 V27 0 2.0247269834162492e-19

R27_28 V27 V28 -377588.261567909
L27_28 V27 V28 6.452154692412963e-11
C27_28 V27 V28 1.1866366287369193e-21

R27_29 V27 V29 55268.25788569403
L27_29 V27 V29 -5.2743646994931705e-11
C27_29 V27 V29 1.0055071129130782e-20

R27_30 V27 V30 -3557603.854764376
L27_30 V27 V30 -1.8733902016073567e-11
C27_30 V27 V30 -1.4568381487631178e-21

R27_31 V27 V31 -22287.57468627628
L27_31 V27 V31 -1.587708780175062e-11
C27_31 V27 V31 5.166959685020803e-20

R27_32 V27 V32 -841948.8184052631
L27_32 V27 V32 3.5578086694813046e-11
C27_32 V27 V32 -4.557263936170785e-21

R27_33 V27 V33 -265286.76125790307
L27_33 V27 V33 -2.862232122319951e-11
C27_33 V27 V33 1.808211312799062e-20

R27_34 V27 V34 -61447.39733426601
L27_34 V27 V34 -4.949803046832948e-10
C27_34 V27 V34 5.889897224710512e-21

R27_35 V27 V35 71707.69282954476
L27_35 V27 V35 4.100038734268165e-11
C27_35 V27 V35 -3.8616890793442807e-20

R27_36 V27 V36 114437.81482155262
L27_36 V27 V36 -1.6328538328805145e-10
C27_36 V27 V36 1.6991192966267335e-21

R27_37 V27 V37 69536.03619640965
L27_37 V27 V37 1.557844728306796e-11
C27_37 V27 V37 3.06931131984587e-20

R27_38 V27 V38 -304830.59092450247
L27_38 V27 V38 -3.201604682448863e-11
C27_38 V27 V38 -6.736024182013312e-21

R27_39 V27 V39 20486.799002395917
L27_39 V27 V39 2.396047335978379e-11
C27_39 V27 V39 7.584016298199939e-20

R27_40 V27 V40 -1894090.7551327788
L27_40 V27 V40 3.092997927214723e-11
C27_40 V27 V40 -1.108538973956587e-20

R27_41 V27 V41 18028.00624164879
L27_41 V27 V41 -6.893111135374837e-12
C27_41 V27 V41 -4.9890560875784127e-20

R27_42 V27 V42 44943.946755259945
L27_42 V27 V42 8.044111325511509e-11
C27_42 V27 V42 -5.913821356208233e-20

R27_43 V27 V43 -27994.75596835832
L27_43 V27 V43 -1.354472033839996e-11
C27_43 V27 V43 -6.192828872023416e-20

R27_44 V27 V44 19128.705329461558
L27_44 V27 V44 3.153627547519127e-11
C27_44 V27 V44 8.282582512335766e-20

R27_45 V27 V45 8647.221818426262
L27_45 V27 V45 6.4846377276005355e-12
C27_45 V27 V45 1.6981018912400392e-19

R27_46 V27 V46 -78594.75663209883
L27_46 V27 V46 -6.247463548942376e-12
C27_46 V27 V46 -9.237531986808386e-20

R27_47 V27 V47 -46115.05553741393
L27_47 V27 V47 -8.146666208102039e-12
C27_47 V27 V47 -4.7918052043512195e-20

R27_48 V27 V48 858733.3466477738
L27_48 V27 V48 -5.946902135310318e-11
C27_48 V27 V48 -2.9158800611677164e-20

R27_49 V27 V49 -55250.49973781931
L27_49 V27 V49 3.314003598004506e-11
C27_49 V27 V49 -6.560573244771038e-20

R27_50 V27 V50 62396.009083329795
L27_50 V27 V50 3.06831191017767e-11
C27_50 V27 V50 4.130789761674451e-20

R27_51 V27 V51 -136586.43399090288
L27_51 V27 V51 -2.988412045816719e-11
C27_51 V27 V51 2.2512482631363676e-20

R27_52 V27 V52 -45860.053672076014
L27_52 V27 V52 9.793110810741913e-11
C27_52 V27 V52 -3.688710283057103e-20

R27_53 V27 V53 -382552.61969181907
L27_53 V27 V53 -5.636486188568424e-11
C27_53 V27 V53 -2.1144310280928105e-20

R27_54 V27 V54 33913.6916055161
L27_54 V27 V54 -2.3604929457109697e-11
C27_54 V27 V54 -1.6395959480396643e-20

R27_55 V27 V55 24481.31748078138
L27_55 V27 V55 -3.646408656416518e-11
C27_55 V27 V55 -7.085384315607998e-20

R27_56 V27 V56 83953.82790004164
L27_56 V27 V56 -1.1213208630165967e-11
C27_56 V27 V56 -2.0865861494167798e-20

R27_57 V27 V57 3582.262687297055
L27_57 V27 V57 -7.848631240453278e-12
C27_57 V27 V57 6.679369392242549e-21

R27_58 V27 V58 7295.6313117153895
L27_58 V27 V58 -9.058737082175285e-11
C27_58 V27 V58 -4.479640863417494e-21

R27_59 V27 V59 -30494.067706764858
L27_59 V27 V59 -7.667205124849037e-12
C27_59 V27 V59 1.1524751493580416e-20

R27_60 V27 V60 9334.88293575325
L27_60 V27 V60 -1.4425979336688599e-11
C27_60 V27 V60 -2.561486115174908e-21

R27_61 V27 V61 -10561.50007136229
L27_61 V27 V61 6.159343097160162e-11
C27_61 V27 V61 -2.350878626435192e-20

R27_62 V27 V62 -8495.686390372266
L27_62 V27 V62 -2.2137810618895335e-10
C27_62 V27 V62 -1.2706821365191712e-20

R27_63 V27 V63 44051.3219088873
L27_63 V27 V63 -1.682796867997409e-11
C27_63 V27 V63 -2.1275520304337312e-20

R27_64 V27 V64 298557.3707895368
L27_64 V27 V64 -2.4447238185411473e-11
C27_64 V27 V64 5.44003629273294e-22

R27_65 V27 V65 8297.472096118303
L27_65 V27 V65 1.5595671928906288e-11
C27_65 V27 V65 7.321911398069493e-21

R27_66 V27 V66 8338.052250210434
L27_66 V27 V66 2.558995894731856e-11
C27_66 V27 V66 -2.6926302199850512e-20

R27_67 V27 V67 -46365.138466096934
L27_67 V27 V67 -9.216274353943245e-12
C27_67 V27 V67 -2.1187044093627665e-20

R27_68 V27 V68 35506.51105723352
L27_68 V27 V68 4.637178176050183e-11
C27_68 V27 V68 -6.649646443809293e-22

R27_69 V27 V69 -27945.319614813343
L27_69 V27 V69 1.2529168878120977e-11
C27_69 V27 V69 1.8288945693398487e-20

R27_70 V27 V70 -52051.323799708385
L27_70 V27 V70 -5.7981121340586934e-12
C27_70 V27 V70 -1.7048782765740428e-20

R27_71 V27 V71 38707.45280655805
L27_71 V27 V71 3.305004580894866e-11
C27_71 V27 V71 2.0942169638088016e-22

R27_72 V27 V72 -19428.903117311427
L27_72 V27 V72 -5.0093625813633884e-12
C27_72 V27 V72 -6.717747471074213e-21

R27_73 V27 V73 -76993.82651866734
L27_73 V27 V73 -1.6743384146165096e-11
C27_73 V27 V73 -6.961107107554212e-21

R27_74 V27 V74 -30236.747422726392
L27_74 V27 V74 6.889084685045944e-11
C27_74 V27 V74 3.0767345965800327e-21

R27_75 V27 V75 64775.31405428626
L27_75 V27 V75 9.303717390733294e-12
C27_75 V27 V75 -1.803185385965453e-21

R27_76 V27 V76 107835.60362684446
L27_76 V27 V76 -2.8654336024789076e-11
C27_76 V27 V76 -8.551436159591949e-21

R27_77 V27 V77 153789.54297648623
L27_77 V27 V77 -8.468236304429944e-11
C27_77 V27 V77 4.625843327011593e-21

R27_78 V27 V78 -102474.00300431513
L27_78 V27 V78 -1.0009834883660565e-11
C27_78 V27 V78 -5.6275080852486586e-21

R27_79 V27 V79 -60543.54737848026
L27_79 V27 V79 -1.2100800164371049e-11
C27_79 V27 V79 -1.0671109079510223e-20

R27_80 V27 V80 -668122.646753427
L27_80 V27 V80 -4.47123392687256e-11
C27_80 V27 V80 1.792278574255242e-20

R27_81 V27 V81 -146317.75963690726
L27_81 V27 V81 8.370258995854236e-12
C27_81 V27 V81 -1.5683754870169872e-20

R27_82 V27 V82 2621409.9962169137
L27_82 V27 V82 2.8823690102621846e-12
C27_82 V27 V82 1.9567638459661046e-21

R27_83 V27 V83 81908.03167125492
L27_83 V27 V83 4.954201963868058e-12
C27_83 V27 V83 5.9058618032350856e-21

R27_84 V27 V84 -137500.492782503
L27_84 V27 V84 -1.1410171324224155e-11
C27_84 V27 V84 -8.123234035538101e-21

R27_85 V27 V85 -87753.86123397516
L27_85 V27 V85 -7.10104465869953e-12
C27_85 V27 V85 -1.061911714242895e-20

R27_86 V27 V86 -86707.09430435541
L27_86 V27 V86 -5.859502895718566e-12
C27_86 V27 V86 -4.615913018268034e-21

R27_87 V27 V87 -269357.4759168906
L27_87 V27 V87 -5.686393636565939e-12
C27_87 V27 V87 -1.3053769300999133e-20

R27_88 V27 V88 -96564.85555118136
L27_88 V27 V88 -1.063424952265195e-10
C27_88 V27 V88 -4.8096887473564525e-21

R27_89 V27 V89 249401.67444170653
L27_89 V27 V89 1.9419753317370873e-11
C27_89 V27 V89 7.759546460467692e-21

R27_90 V27 V90 72817.41355178201
L27_90 V27 V90 1.46151428755357e-11
C27_90 V27 V90 9.467881679382577e-21

R27_91 V27 V91 1118256.5058203978
L27_91 V27 V91 2.6963148744426926e-12
C27_91 V27 V91 7.200934883589005e-22

R27_92 V27 V92 157875.38277292295
L27_92 V27 V92 6.81268849759793e-11
C27_92 V27 V92 1.8064821400219154e-20

R27_93 V27 V93 -26503.90183913454
L27_93 V27 V93 -2.6320958775281378e-11
C27_93 V27 V93 -9.451892692604762e-22

R27_94 V27 V94 -38097.29277719266
L27_94 V27 V94 -2.962152244613898e-11
C27_94 V27 V94 -2.345634994566819e-21

R27_95 V27 V95 -921020.9714495227
L27_95 V27 V95 5.723967498020256e-12
C27_95 V27 V95 4.1556749076633434e-22

R27_96 V27 V96 212444.13880375706
L27_96 V27 V96 -8.484316164972004e-12
C27_96 V27 V96 1.599311097118176e-20

R27_97 V27 V97 255825.93003885896
L27_97 V27 V97 -3.109282343633858e-11
C27_97 V27 V97 3.910287585170769e-22

R27_98 V27 V98 39306.766478485435
L27_98 V27 V98 9.764167693819698e-12
C27_98 V27 V98 8.00952544708398e-21

R27_99 V27 V99 -59582.36787057087
L27_99 V27 V99 -3.857723223581195e-11
C27_99 V27 V99 -1.5212730083145933e-21

R27_100 V27 V100 -151346.5687152697
L27_100 V27 V100 6.36272070931799e-11
C27_100 V27 V100 -7.090410530309571e-21

R27_101 V27 V101 -169480.39980397376
L27_101 V27 V101 1.0265463494741804e-11
C27_101 V27 V101 1.1684579901452373e-20

R27_102 V27 V102 89140.74769543484
L27_102 V27 V102 4.4202566705153245e-12
C27_102 V27 V102 1.678923238041613e-20

R27_103 V27 V103 -140650.7381553328
L27_103 V27 V103 -1.2460949425132906e-11
C27_103 V27 V103 -1.5073520838536427e-20

R27_104 V27 V104 -195703.34892977666
L27_104 V27 V104 -5.610306346816921e-12
C27_104 V27 V104 1.2820316673616938e-20

R27_105 V27 V105 1302793.002211741
L27_105 V27 V105 -5.6838635882828994e-12
C27_105 V27 V105 -9.604082759886083e-21

R27_106 V27 V106 -113108.66474600077
L27_106 V27 V106 2.560349298015102e-12
C27_106 V27 V106 1.820495145304433e-20

R27_107 V27 V107 175263.683251639
L27_107 V27 V107 5.409105113666843e-12
C27_107 V27 V107 1.2940291255359197e-20

R27_108 V27 V108 60273.699809452904
L27_108 V27 V108 -8.483765353203391e-12
C27_108 V27 V108 -2.2970703095652398e-20

R27_109 V27 V109 69954.4612195279
L27_109 V27 V109 -5.690234376084248e-12
C27_109 V27 V109 7.821864101719425e-21

R27_110 V27 V110 53068.83019368767
L27_110 V27 V110 -3.804559420770583e-12
C27_110 V27 V110 -5.877642100981143e-21

R27_111 V27 V111 2801853.1937301788
L27_111 V27 V111 -6.7445985417688494e-12
C27_111 V27 V111 -7.711883214788016e-21

R27_112 V27 V112 19288.34640596558
L27_112 V27 V112 6.1434380438511796e-12
C27_112 V27 V112 1.7060232777661678e-20

R27_113 V27 V113 31680.39100673045
L27_113 V27 V113 7.2394880681192766e-12
C27_113 V27 V113 -8.565259381236544e-23

R27_114 V27 V114 -109576.47673548866
L27_114 V27 V114 6.349467780625417e-12
C27_114 V27 V114 4.279392390876789e-21

R27_115 V27 V115 133747.2070876883
L27_115 V27 V115 1.0015017564078828e-11
C27_115 V27 V115 1.101722656961963e-20

R27_116 V27 V116 -67576.34265328385
L27_116 V27 V116 -1.2278301635987299e-11
C27_116 V27 V116 -1.4066868582799362e-20

R27_117 V27 V117 -331304.1182083477
L27_117 V27 V117 -1.0046027949351267e-11
C27_117 V27 V117 -4.556428280788997e-21

R27_118 V27 V118 -246002.10419695725
L27_118 V27 V118 -4.721452061621504e-12
C27_118 V27 V118 -3.144269985894938e-21

R27_119 V27 V119 55844.052824046346
L27_119 V27 V119 -5.685043219745974e-12
C27_119 V27 V119 -1.0668715412406956e-20

R27_120 V27 V120 96211.15910611514
L27_120 V27 V120 1.1874985513365832e-11
C27_120 V27 V120 -9.380255084430229e-21

R27_121 V27 V121 17484.291212507156
L27_121 V27 V121 2.4115147336489806e-11
C27_121 V27 V121 -1.635324163194489e-21

R27_122 V27 V122 7970.77172072519
L27_122 V27 V122 1.1905186614350531e-11
C27_122 V27 V122 4.561527883680906e-21

R27_123 V27 V123 219875.1126903715
L27_123 V27 V123 -4.632258001157402e-11
C27_123 V27 V123 2.5866093828046638e-21

R27_124 V27 V124 -78004.77014997594
L27_124 V27 V124 -5.1587111264416024e-11
C27_124 V27 V124 -4.232329005148981e-21

R27_125 V27 V125 -18388.917792501823
L27_125 V27 V125 2.084539431764738e-10
C27_125 V27 V125 -1.726697251252346e-21

R27_126 V27 V126 -8929.052638880132
L27_126 V27 V126 -9.532273721168553e-12
C27_126 V27 V126 1.7954415435634873e-21

R27_127 V27 V127 14414.432823463829
L27_127 V27 V127 6.959339959430422e-12
C27_127 V27 V127 3.891447010638302e-22

R27_128 V27 V128 75739.37761466004
L27_128 V27 V128 7.351307055876e-11
C27_128 V27 V128 1.2803107754044708e-21

R27_129 V27 V129 110417.54302386903
L27_129 V27 V129 2.519333444117626e-11
C27_129 V27 V129 1.5505529566960568e-21

R27_130 V27 V130 19816191.274454236
L27_130 V27 V130 -1.9769362494252252e-11
C27_130 V27 V130 -3.598606789912206e-21

R27_131 V27 V131 -63374.39715428639
L27_131 V27 V131 3.510156011586814e-11
C27_131 V27 V131 3.619850348265751e-21

R27_132 V27 V132 -45838.038922985696
L27_132 V27 V132 3.77300154688173e-11
C27_132 V27 V132 -1.0214658922527083e-21

R27_133 V27 V133 -81502.51682947422
L27_133 V27 V133 7.01184462203989e-12
C27_133 V27 V133 7.084904455272482e-21

R27_134 V27 V134 -73502.62820298255
L27_134 V27 V134 2.344502416409549e-09
C27_134 V27 V134 -2.3802628371823838e-22

R27_135 V27 V135 21628.347650314525
L27_135 V27 V135 1.6282958702333043e-11
C27_135 V27 V135 -2.1552319979884062e-21

R27_136 V27 V136 580881.5622186037
L27_136 V27 V136 -7.643146694850887e-11
C27_136 V27 V136 -2.8508000506181363e-21

R27_137 V27 V137 -23929.572055964316
L27_137 V27 V137 -2.6490819885554604e-11
C27_137 V27 V137 -4.678051837226331e-21

R27_138 V27 V138 -10666.948301292952
L27_138 V27 V138 -1.4900477947447684e-11
C27_138 V27 V138 -1.347069382408722e-21

R27_139 V27 V139 11686.573702865784
L27_139 V27 V139 5.446997475287682e-12
C27_139 V27 V139 4.390005597738569e-21

R27_140 V27 V140 -69817.3368415734
L27_140 V27 V140 -1.9135757464008394e-11
C27_140 V27 V140 -7.108288729984781e-22

R27_141 V27 V141 -28813.570978030642
L27_141 V27 V141 -4.506640612180179e-11
C27_141 V27 V141 1.8932933057380108e-21

R27_142 V27 V142 -317849.3390255908
L27_142 V27 V142 -2.4190480346098748e-11
C27_142 V27 V142 1.46031056457285e-21

R27_143 V27 V143 -53087.34289976756
L27_143 V27 V143 -2.5294908465996615e-11
C27_143 V27 V143 -2.30466353171721e-21

R27_144 V27 V144 50192.663112133436
L27_144 V27 V144 9.56572651080951e-10
C27_144 V27 V144 -1.1681657460244261e-21

R28_28 V28 0 -4045.077438334116
L28_28 V28 0 7.546622258353273e-13
C28_28 V28 0 2.012252410122981e-19

R28_29 V28 V29 77845.69974938044
L28_29 V28 V29 1.7307972646179373e-10
C28_29 V28 V29 4.127912601407705e-21

R28_30 V28 V30 548838.2276327942
L28_30 V28 V30 -4.0735486514849955e-11
C28_30 V28 V30 -1.9393005408330263e-21

R28_31 V28 V31 -7232724.870305528
L28_31 V28 V31 -1.0921676388094775e-10
C28_31 V28 V31 -1.3205228152326811e-21

R28_32 V28 V32 -68341.74359894783
L28_32 V28 V32 -3.984289150657556e-12
C28_32 V28 V32 7.181974201980697e-21

R28_33 V28 V33 -4031781.0974631603
L28_33 V28 V33 -5.945193424726025e-11
C28_33 V28 V33 2.3672252363264297e-21

R28_34 V28 V34 -205026.10501055603
L28_34 V28 V34 -7.737852005295971e-10
C28_34 V28 V34 -2.356078149071189e-21

R28_35 V28 V35 6270839.0592221515
L28_35 V28 V35 -4.287878664941501e-11
C28_35 V28 V35 2.7971303900948734e-21

R28_36 V28 V36 -216902.41110952714
L28_36 V28 V36 1.508384536613095e-11
C28_36 V28 V36 -9.869876873734457e-21

R28_37 V28 V37 -6187808.959174854
L28_37 V28 V37 2.5891327534467364e-11
C28_37 V28 V37 7.460966223054042e-21

R28_38 V28 V38 -256933.86628114828
L28_38 V28 V38 6.711596152104364e-11
C28_38 V28 V38 -3.7826563388916504e-21

R28_39 V28 V39 602092.7124433054
L28_39 V28 V39 7.860719200028611e-11
C28_39 V28 V39 -1.2781274391901631e-21

R28_40 V28 V40 20082.484924404584
L28_40 V28 V40 -9.03030723600119e-12
C28_40 V28 V40 4.7600199513547934e-20

R28_41 V28 V41 69413.33176735684
L28_41 V28 V41 -9.834965697948373e-12
C28_41 V28 V41 -3.7933597953544736e-20

R28_42 V28 V42 71221.87416078769
L28_42 V28 V42 -1.100233318690979e-10
C28_42 V28 V42 -9.089866472490752e-21

R28_43 V28 V43 -601546.7430225624
L28_43 V28 V43 -5.131164248267835e-10
C28_43 V28 V43 -1.27572439998644e-22

R28_44 V28 V44 -16528.95785480844
L28_44 V28 V44 4.354662785484143e-12
C28_44 V28 V44 -7.761920087685165e-20

R28_45 V28 V45 24162.482486211087
L28_45 V28 V45 -1.3832049926039159e-11
C28_45 V28 V45 5.060733415558876e-20

R28_46 V28 V46 108059.62948067041
L28_46 V28 V46 8.012466614083877e-12
C28_46 V28 V46 -7.324257330903611e-21

R28_47 V28 V47 593909.3713278398
L28_47 V28 V47 -7.304389638066341e-11
C28_47 V28 V47 -4.752226835477754e-21

R28_48 V28 V48 -51646.35535983448
L28_48 V28 V48 2.224921619203118e-11
C28_48 V28 V48 1.1371325685475511e-20

R28_49 V28 V49 -121017.15827490266
L28_49 V28 V49 -4.041596452700866e-11
C28_49 V28 V49 -1.0681433889451228e-20

R28_50 V28 V50 10096691.703695672
L28_50 V28 V50 1.4633247014828472e-11
C28_50 V28 V50 -3.749767954710387e-21

R28_51 V28 V51 -137049.89521352228
L28_51 V28 V51 -5.5058158115889824e-11
C28_51 V28 V51 4.046019301398118e-21

R28_52 V28 V52 -132123.45430528978
L28_52 V28 V52 1.7790452566825053e-11
C28_52 V28 V52 -2.86563635958684e-20

R28_53 V28 V53 -94546.38573074418
L28_53 V28 V53 -3.256901117652138e-11
C28_53 V28 V53 1.0138060721285921e-20

R28_54 V28 V54 75815.3791680981
L28_54 V28 V54 -2.8752944271988593e-11
C28_54 V28 V54 1.6892615134974206e-21

R28_55 V28 V55 57534.51789824211
L28_55 V28 V55 1.8042883915313692e-11
C28_55 V28 V55 -9.742652500596957e-21

R28_56 V28 V56 37030.99098242232
L28_56 V28 V56 -3.425408774962445e-11
C28_56 V28 V56 -6.552329665568523e-20

R28_57 V28 V57 8986.56866160902
L28_57 V28 V57 -9.372444853685251e-12
C28_57 V28 V57 1.6828763357217049e-22

R28_58 V28 V58 15222.998439266756
L28_58 V28 V58 -6.889310250510303e-12
C28_58 V28 V58 -2.6288407204364818e-21

R28_59 V28 V59 79969.06566972332
L28_59 V28 V59 -3.2902264911763125e-11
C28_59 V28 V59 -1.5498632522982438e-21

R28_60 V28 V60 2001985.3359034173
L28_60 V28 V60 6.140631518958803e-12
C28_60 V28 V60 3.6869666768565526e-21

R28_61 V28 V61 -25701.283820471846
L28_61 V28 V61 -1.508311661349515e-11
C28_61 V28 V61 -1.367300899734443e-20

R28_62 V28 V62 -21961.31448029487
L28_62 V28 V62 2.0291200999450003e-11
C28_62 V28 V62 -1.8056747026576154e-21

R28_63 V28 V63 71000.01922315742
L28_63 V28 V63 2.575894682586186e-11
C28_63 V28 V63 -9.342862693461366e-21

R28_64 V28 V64 -34163.081128598526
L28_64 V28 V64 -6.766178688235636e-12
C28_64 V28 V64 -5.071414104495163e-20

R28_65 V28 V65 23688.195243923295
L28_65 V28 V65 2.560021461291004e-11
C28_65 V28 V65 1.0221645733990293e-20

R28_66 V28 V66 67910.42863097784
L28_66 V28 V66 -6.322646484970151e-12
C28_66 V28 V66 -2.2883756980452718e-20

R28_67 V28 V67 -75124.97982467948
L28_67 V28 V67 -4.5920613257427104e-11
C28_67 V28 V67 -1.1693523822844134e-20

R28_68 V28 V68 117178.49818822491
L28_68 V28 V68 1.4333145462310442e-11
C28_68 V28 V68 -1.0845818935699548e-20

R28_69 V28 V69 -47106.98711893173
L28_69 V28 V69 -9.796929406512101e-12
C28_69 V28 V69 -1.7141338147762827e-21

R28_70 V28 V70 568978.7952926045
L28_70 V28 V70 -4.591194235607807e-12
C28_70 V28 V70 -2.210164579458155e-20

R28_71 V28 V71 97310.94911807701
L28_71 V28 V71 9.740869011728466e-11
C28_71 V28 V71 -4.093054452563922e-21

R28_72 V28 V72 -96510.45086582066
L28_72 V28 V72 -9.577061946134636e-12
C28_72 V28 V72 -7.006134607830025e-21

R28_73 V28 V73 190072.75440651964
L28_73 V28 V73 -5.0720557988809265e-12
C28_73 V28 V73 -1.792135293027311e-20

R28_74 V28 V74 -114295.51538176011
L28_74 V28 V74 -2.0928648049089312e-11
C28_74 V28 V74 4.376988321291001e-21

R28_75 V28 V75 -978468.7234369877
L28_75 V28 V75 8.577907100520976e-12
C28_75 V28 V75 1.3094512972315305e-20

R28_76 V28 V76 -86560.11202909854
L28_76 V28 V76 -6.0948205559372544e-12
C28_76 V28 V76 -1.4718826561855923e-20

R28_77 V28 V77 79695.53223022015
L28_77 V28 V77 5.6643206828887846e-12
C28_77 V28 V77 2.2115355325118598e-20

R28_78 V28 V78 -78071.99333414569
L28_78 V28 V78 -8.521511528252252e-12
C28_78 V28 V78 -1.7514434879741005e-20

R28_79 V28 V79 -161043.8816687389
L28_79 V28 V79 -6.7056861272216485e-12
C28_79 V28 V79 -9.994567681756376e-21

R28_80 V28 V80 89489.92531588247
L28_80 V28 V80 2.716656134159711e-12
C28_80 V28 V80 3.437676999296108e-20

R28_81 V28 V81 -45565.87737126386
L28_81 V28 V81 -1.4617208315803801e-12
C28_81 V28 V81 -6.011444329037758e-20

R28_82 V28 V82 133445.61601134305
L28_82 V28 V82 2.8573923447846936e-12
C28_82 V28 V82 3.631461322347684e-20

R28_83 V28 V83 45323.706903124825
L28_83 V28 V83 1.9679586790792784e-12
C28_83 V28 V83 4.63494457512394e-20

R28_84 V28 V84 343019.51688788057
L28_84 V28 V84 7.18912422232188e-10
C28_84 V28 V84 -1.3243996507224388e-21

R28_85 V28 V85 -225112.80915476382
L28_85 V28 V85 -3.792680971589689e-12
C28_85 V28 V85 -2.4675620359633652e-20

R28_86 V28 V86 -176778.76026491026
L28_86 V28 V86 -6.4630644880550696e-12
C28_86 V28 V86 -1.3365010897282178e-20

R28_87 V28 V87 -71089.91251525069
L28_87 V28 V87 -3.3546865207217566e-12
C28_87 V28 V87 -2.8347151264792396e-20

R28_88 V28 V88 -74927.37342813314
L28_88 V28 V88 -5.7280120354036876e-12
C28_88 V28 V88 -1.6046882420862876e-20

R28_89 V28 V89 153371.7765462616
L28_89 V28 V89 6.003984750534867e-12
C28_89 V28 V89 2.4125465753258965e-20

R28_90 V28 V90 175361.00235478318
L28_90 V28 V90 1.8778625107169704e-11
C28_90 V28 V90 7.939242977509078e-21

R28_91 V28 V91 107711.44247682882
L28_91 V28 V91 6.6298307980392006e-12
C28_91 V28 V91 2.2520994037460743e-20

R28_92 V28 V92 47084.022578462915
L28_92 V28 V92 1.5345666254757297e-12
C28_92 V28 V92 5.927812429271601e-20

R28_93 V28 V93 -56059.98781529781
L28_93 V28 V93 -9.299769986428205e-12
C28_93 V28 V93 -7.410492788957072e-21

R28_94 V28 V94 -46826.19455466439
L28_94 V28 V94 -3.358697929818669e-12
C28_94 V28 V94 -3.1391580988337064e-20

R28_95 V28 V95 273025.8417000497
L28_95 V28 V95 6.567722036934978e-12
C28_95 V28 V95 1.6981032111356263e-20

R28_96 V28 V96 42547.45646436876
L28_96 V28 V96 1.409800560938635e-12
C28_96 V28 V96 6.147597043089564e-20

R28_97 V28 V97 -467107.53547723393
L28_97 V28 V97 -4.06787986694595e-12
C28_97 V28 V97 -1.9047591152949994e-20

R28_98 V28 V98 42459.05388784128
L28_98 V28 V98 3.013349693442163e-12
C28_98 V28 V98 3.1135983454423865e-20

R28_99 V28 V99 -98637.70251670181
L28_99 V28 V99 -1.0040301439677883e-11
C28_99 V28 V99 -8.205576072130466e-21

R28_100 V28 V100 -142550.62303663653
L28_100 V28 V100 -3.70898066602725e-12
C28_100 V28 V100 -1.920738368952526e-20

R28_101 V28 V101 142593.1444024444
L28_101 V28 V101 2.9661282774506185e-12
C28_101 V28 V101 3.582159945071926e-20

R28_102 V28 V102 90713.57298371167
L28_102 V28 V102 3.947806943069473e-12
C28_102 V28 V102 2.6181414368302504e-20

R28_103 V28 V103 -687708.8004538156
L28_103 V28 V103 -6.924782710765828e-12
C28_103 V28 V103 -9.516357334342872e-21

R28_104 V28 V104 133525.17330860082
L28_104 V28 V104 2.5427027518033034e-12
C28_104 V28 V104 4.0230476300619555e-20

R28_105 V28 V105 -88017.16160191773
L28_105 V28 V105 -2.4181782724139074e-12
C28_105 V28 V105 -4.184073821220991e-20

R28_106 V28 V106 86537.37719015604
L28_106 V28 V106 1.7987940157217772e-12
C28_106 V28 V106 5.589240836500423e-20

R28_107 V28 V107 146093.15232158673
L28_107 V28 V107 4.103168034522606e-12
C28_107 V28 V107 1.9222663211588747e-20

R28_108 V28 V108 322622.35271573556
L28_108 V28 V108 -2.2478738516379695e-12
C28_108 V28 V108 -3.945967465177262e-20

R28_109 V28 V109 110307.3624158833
L28_109 V28 V109 3.947374354500213e-12
C28_109 V28 V109 2.6222684858620693e-20

R28_110 V28 V110 -207218.04038798824
L28_110 V28 V110 -2.1347409093545193e-12
C28_110 V28 V110 -4.924580070890167e-20

R28_111 V28 V111 -430352.7186265255
L28_111 V28 V111 -3.458628291269688e-12
C28_111 V28 V111 -2.2200430336841302e-20

R28_112 V28 V112 32341.48875574867
L28_112 V28 V112 2.9682092661363323e-12
C28_112 V28 V112 2.8853254228265157e-20

R28_113 V28 V113 59773.90654202465
L28_113 V28 V113 -1.0822441528019665e-10
C28_113 V28 V113 1.1947643851066556e-21

R28_114 V28 V114 90913.44891555993
L28_114 V28 V114 3.589134520441585e-12
C28_114 V28 V114 2.8030534681509825e-20

R28_115 V28 V115 171491.63634119404
L28_115 V28 V115 7.261363948209884e-12
C28_115 V28 V115 1.1846492223861986e-20

R28_116 V28 V116 -81211.99660028977
L28_116 V28 V116 -3.3070584906896337e-12
C28_116 V28 V116 -2.955015687232527e-20

R28_117 V28 V117 -1617998.8331099171
L28_117 V28 V117 -3.4918107110593654e-11
C28_117 V28 V117 -7.604896166851763e-21

R28_118 V28 V118 -124077.34730841214
L28_118 V28 V118 -8.883741868969293e-12
C28_118 V28 V118 -1.2163189468401516e-20

R28_119 V28 V119 -141295.19091786846
L28_119 V28 V119 -2.5080211169844323e-12
C28_119 V28 V119 -3.9650336187056943e-20

R28_120 V28 V120 559415.353153689
L28_120 V28 V120 -6.897198448598241e-12
C28_120 V28 V120 -1.658621757243299e-20

R28_121 V28 V121 37307.39943384819
L28_121 V28 V121 6.652087624280805e-11
C28_121 V28 V121 3.5622030111832766e-21

R28_122 V28 V122 15882.324832227565
L28_122 V28 V122 1.6838481966052692e-10
C28_122 V28 V122 2.609044828113e-21

R28_123 V28 V123 104437.59301000478
L28_123 V28 V123 -1.589200714315734e-11
C28_123 V28 V123 -1.820516145270634e-21

R28_124 V28 V124 2459846.7914722105
L28_124 V28 V124 -5.815208413916828e-12
C28_124 V28 V124 -1.6945128880194085e-20

R28_125 V28 V125 -38603.53227039437
L28_125 V28 V125 -2.2794037270526408e-11
C28_125 V28 V125 -6.29284323546293e-21

R28_126 V28 V126 -19144.64348592474
L28_126 V28 V126 3.713033911587314e-11
C28_126 V28 V126 3.209384700513369e-21

R28_127 V28 V127 29502.04125127803
L28_127 V28 V127 2.328514002706012e-11
C28_127 V28 V127 -1.7526523143679854e-21

R28_128 V28 V128 -361998.79801188793
L28_128 V28 V128 1.72806419833012e-11
C28_128 V28 V128 -1.7484530925464035e-21

R28_129 V28 V129 63004.7418534029
L28_129 V28 V129 -1.6601916331946947e-11
C28_129 V28 V129 -5.644559839773881e-21

R28_130 V28 V130 -60838.398982825776
L28_130 V28 V130 5.7446951280485136e-11
C28_130 V28 V130 -1.080748565283873e-20

R28_131 V28 V131 -52788.211839014024
L28_131 V28 V131 7.457565051410522e-12
C28_131 V28 V131 4.841525105919835e-21

R28_132 V28 V132 -59530.699309599666
L28_132 V28 V132 -9.699433541999981e-12
C28_132 V28 V132 -8.374948958774645e-21

R28_133 V28 V133 -462283.2923316358
L28_133 V28 V133 5.498450911460708e-12
C28_133 V28 V133 1.7826549845309268e-20

R28_134 V28 V134 -96660.64661869922
L28_134 V28 V134 6.126611507254507e-11
C28_134 V28 V134 -1.6103822684984705e-21

R28_135 V28 V135 44449.38872697468
L28_135 V28 V135 -1.4321419517299527e-10
C28_135 V28 V135 -1.7025817903253102e-21

R28_136 V28 V136 604460.9108473036
L28_136 V28 V136 1.2048901056610907e-10
C28_136 V28 V136 3.844513888520143e-21

R28_137 V28 V137 -53091.54700708936
L28_137 V28 V137 -1.4584303960757537e-11
C28_137 V28 V137 -8.434114991517111e-21

R28_138 V28 V138 -19376.059976396624
L28_138 V28 V138 9.720118753907703e-11
C28_138 V28 V138 -1.584238045727144e-21

R28_139 V28 V139 22992.843532107025
L28_139 V28 V139 1.3841841766850992e-11
C28_139 V28 V139 5.045443432848431e-21

R28_140 V28 V140 -74322.63888832428
L28_140 V28 V140 -2.3513233502136123e-11
C28_140 V28 V140 -3.430055633975587e-21

R28_141 V28 V141 -172480.13128702482
L28_141 V28 V141 -2.977771301971928e-11
C28_141 V28 V141 3.9526441737590494e-21

R28_142 V28 V142 -67897.46479060309
L28_142 V28 V142 1.302852188932014e-10
C28_142 V28 V142 -4.992100223422333e-21

R28_143 V28 V143 -77211.27199743185
L28_143 V28 V143 1.933516832601799e-10
C28_143 V28 V143 -2.459615797616282e-21

R28_144 V28 V144 80266.34835972796
L28_144 V28 V144 1.0912343810410121e-11
C28_144 V28 V144 2.2285502993815606e-21

R29_29 V29 0 -694.8550317121048
L29_29 V29 0 -6.62441509170209e-14
C29_29 V29 0 -2.2504887370028026e-18

R29_30 V29 V30 -39137.65125297286
L29_30 V29 V30 1.608629761415951e-11
C29_30 V29 V30 -2.96451455310506e-20

R29_31 V29 V31 -17760.072762886888
L29_31 V29 V31 3.283479030560862e-11
C29_31 V29 V31 -3.4923277021197735e-20

R29_32 V29 V32 -59471.72074501733
L29_32 V29 V32 1.8256359571070924e-11
C29_32 V29 V32 -2.092770984725479e-20

R29_33 V29 V33 6817.976490814675
L29_33 V29 V33 1.5114923714613278e-12
C29_33 V29 V33 5.3882864883192404e-20

R29_34 V29 V34 -24745.33843961355
L29_34 V29 V34 -3.5946150553955956e-12
C29_34 V29 V34 -1.598710953399166e-20

R29_35 V29 V35 13600.619614442683
L29_35 V29 V35 2.8887597277415166e-12
C29_35 V29 V35 3.2104853533584765e-20

R29_36 V29 V36 -237857.88408365299
L29_36 V29 V36 -7.06748566407004e-12
C29_36 V29 V36 5.5040273539875645e-21

R29_37 V29 V37 -7762.8899384738215
L29_37 V29 V37 -8.904918328253458e-13
C29_37 V29 V37 -3.0883646133640073e-19

R29_38 V29 V38 53380.39913732654
L29_38 V29 V38 -1.1857536378710005e-10
C29_38 V29 V38 -5.787363113710448e-21

R29_39 V29 V39 -9170.314113631259
L29_39 V29 V39 -1.1022286071862322e-12
C29_39 V29 V39 -2.2247516297201225e-19

R29_40 V29 V40 -974455.9984909779
L29_40 V29 V40 -7.830117945921109e-11
C29_40 V29 V40 -2.4703475288745722e-20

R29_41 V29 V41 2208.5326363997488
L29_41 V29 V41 2.5516328227999877e-13
C29_41 V29 V41 9.693698329006797e-19

R29_42 V29 V42 3051.1606459652317
L29_42 V29 V42 3.711616799433919e-13
C29_42 V29 V42 6.879198984274756e-19

R29_43 V29 V43 5932.511611315017
L29_43 V29 V43 7.454280035693042e-13
C29_43 V29 V43 3.498626082837557e-19

R29_44 V29 V44 60954.14229320281
L29_44 V29 V44 1.6959371711718133e-11
C29_44 V29 V44 2.6455466912091724e-20

R29_45 V29 V45 -3342.6651160371002
L29_45 V29 V45 -7.206434872441803e-13
C29_45 V29 V45 -7.408490511689539e-19

R29_46 V29 V46 -8937.863408223844
L29_46 V29 V46 -4.2718211001886954e-12
C29_46 V29 V46 -3.0788936016322957e-19

R29_47 V29 V47 -34516.487425671956
L29_47 V29 V47 9.842669484518197e-12
C29_47 V29 V47 -1.0407283746438696e-19

R29_48 V29 V48 -27596.07456703768
L29_48 V29 V48 -4.36298700737592e-12
C29_48 V29 V48 -2.976648052177036e-20

R29_49 V29 V49 14698.136198572436
L29_49 V29 V49 3.794245248813694e-12
C29_49 V29 V49 1.807245862491168e-19

R29_50 V29 V50 8522.088549929693
L29_50 V29 V50 1.449224705867389e-12
C29_50 V29 V50 1.4315463892601847e-19

R29_51 V29 V51 -15114.477223145808
L29_51 V29 V51 -1.593675192433685e-12
C29_51 V29 V51 -1.3272746621527594e-19

R29_52 V29 V52 4049.147740196243
L29_52 V29 V52 7.981486146389077e-13
C29_52 V29 V52 4.523781783873767e-19

R29_53 V29 V53 6790.23663425428
L29_53 V29 V53 1.1601162232589195e-12
C29_53 V29 V53 2.270639617285086e-19

R29_54 V29 V54 28173.150960822957
L29_54 V29 V54 2.2489979458612267e-12
C29_54 V29 V54 3.7250840699915286e-20

R29_55 V29 V55 14590.173766316717
L29_55 V29 V55 1.2630864766915472e-12
C29_55 V29 V55 1.3972148560076387e-19

R29_56 V29 V56 16765.56586010909
L29_56 V29 V56 1.7684095062843315e-12
C29_56 V29 V56 1.2756187616836333e-19

R29_57 V29 V57 20752.601036015734
L29_57 V29 V57 2.894741572043625e-13
C29_57 V29 V57 -7.334629357031442e-20

R29_58 V29 V58 128534.85721102751
L29_58 V29 V58 1.3571670204510839e-12
C29_58 V29 V58 -5.064226064270004e-20

R29_59 V29 V59 49977.500455359026
L29_59 V29 V59 1.2303181544161356e-10
C29_59 V29 V59 -6.369659330191139e-20

R29_60 V29 V60 256727.86617484843
L29_60 V29 V60 2.0179434039564955e-12
C29_60 V29 V60 -1.9636394596138862e-20

R29_61 V29 V61 7237.235385239784
L29_61 V29 V61 -7.701760028007558e-12
C29_61 V29 V61 2.8041958133824195e-19

R29_62 V29 V62 8398.714890649024
L29_62 V29 V62 -3.5557265289338277e-12
C29_62 V29 V62 2.446785261707648e-19

R29_63 V29 V63 95887.1752351108
L29_63 V29 V63 1.0834194195474085e-11
C29_63 V29 V63 5.96549893427964e-20

R29_64 V29 V64 28630.348329118468
L29_64 V29 V64 6.924608277890431e-12
C29_64 V29 V64 3.4180763933621744e-20

R29_65 V29 V65 6225.517053270489
L29_65 V29 V65 6.028380003747641e-13
C29_65 V29 V65 9.055190298097059e-20

R29_66 V29 V66 6573.849995350262
L29_66 V29 V66 6.873108884890102e-13
C29_66 V29 V66 5.024887755310875e-20

R29_67 V29 V67 19855.65684339591
L29_67 V29 V67 3.0171720102073822e-12
C29_67 V29 V67 4.5612676171422735e-20

R29_68 V29 V68 289162.3933281493
L29_68 V29 V68 4.538198381733247e-12
C29_68 V29 V68 3.4462850318454024e-20

R29_69 V29 V69 -20470.116824956338
L29_69 V29 V69 -3.5286815589359085e-12
C29_69 V29 V69 -2.3050897059797722e-20

R29_70 V29 V70 -28368.52860971177
L29_70 V29 V70 -1.6467097889644737e-11
C29_70 V29 V70 2.952215298681611e-20

R29_71 V29 V71 -36245.9238402502
L29_71 V29 V71 -1.3412511405749147e-10
C29_71 V29 V71 1.4635474727756633e-20

R29_72 V29 V72 -16646.835378983724
L29_72 V29 V72 -3.089599280457056e-12
C29_72 V29 V72 1.0391632151884005e-20

R29_73 V29 V73 -149694.17846341286
L29_73 V29 V73 1.0590776237565679e-11
C29_73 V29 V73 4.2391393922746553e-20

R29_74 V29 V74 -18591.69215484723
L29_74 V29 V74 -3.0483198464504266e-12
C29_74 V29 V74 -2.819974916026306e-20

R29_75 V29 V75 18806.22137805584
L29_75 V29 V75 3.911237066221465e-12
C29_75 V29 V75 3.731705582834961e-20

R29_76 V29 V76 16125.99655997881
L29_76 V29 V76 2.43110906744586e-12
C29_76 V29 V76 3.9112276163127294e-20

R29_77 V29 V77 43498.931392097744
L29_77 V29 V77 6.7051722085595966e-12
C29_77 V29 V77 1.0865880363746108e-20

R29_78 V29 V78 58910.48675320524
L29_78 V29 V78 9.673371455472218e-12
C29_78 V29 V78 4.924257229673894e-21

R29_79 V29 V79 -79915.10014456318
L29_79 V29 V79 3.094662237642378e-11
C29_79 V29 V79 9.022100643622276e-21

R29_80 V29 V80 -68064.25258877598
L29_80 V29 V80 -1.599945595863664e-11
C29_80 V29 V80 5.146238994498194e-22

R29_81 V29 V81 -58972.788538314555
L29_81 V29 V81 -4.7505993114000474e-11
C29_81 V29 V81 -4.601454901778834e-21

R29_82 V29 V82 50605.285983867674
L29_82 V29 V82 -7.250538659040964e-11
C29_82 V29 V82 1.5956014888089343e-20

R29_83 V29 V83 -158548.1092582452
L29_83 V29 V83 -7.870833104307613e-12
C29_83 V29 V83 2.6483254566889778e-20

R29_84 V29 V84 -55132.16998990827
L29_84 V29 V84 -8.76699203417124e-12
C29_84 V29 V84 4.940073890564462e-21

R29_85 V29 V85 -41473.66181921171
L29_85 V29 V85 -1.7519370299457576e-11
C29_85 V29 V85 -1.23190148810303e-21

R29_86 V29 V86 -75091.878951954
L29_86 V29 V86 -7.182168404685057e-11
C29_86 V29 V86 -1.2378594572112265e-20

R29_87 V29 V87 -1041140.0882414693
L29_87 V29 V87 -9.746976497220676e-11
C29_87 V29 V87 -7.202743299945732e-21

R29_88 V29 V88 171798.34267396593
L29_88 V29 V88 5.955202212447145e-11
C29_88 V29 V88 5.764132488467827e-22

R29_89 V29 V89 57086.283391018995
L29_89 V29 V89 4.547736519670123e-12
C29_89 V29 V89 6.306813399304576e-21

R29_90 V29 V90 272980.5349671764
L29_90 V29 V90 9.974304728216323e-11
C29_90 V29 V90 2.3479702445979712e-21

R29_91 V29 V91 162974.70076980974
L29_91 V29 V91 -3.1441422779071016e-11
C29_91 V29 V91 2.6442506438544007e-20

R29_92 V29 V92 271054.2332311011
L29_92 V29 V92 -2.8418776674708315e-11
C29_92 V29 V92 1.366729357375304e-20

R29_93 V29 V93 -96442.82503714165
L29_93 V29 V93 -3.8524176471251206e-11
C29_93 V29 V93 -6.4362850763929116e-21

R29_94 V29 V94 -78508.72814670469
L29_94 V29 V94 -1.4770570379312346e-11
C29_94 V29 V94 -8.417860395215392e-21

R29_95 V29 V95 304726.6217894722
L29_95 V29 V95 -2.2304373890949954e-11
C29_95 V29 V95 7.363617213911317e-21

R29_96 V29 V96 1951372.830638611
L29_96 V29 V96 -1.4411938827874109e-11
C29_96 V29 V96 -2.4950830202528e-21

R29_97 V29 V97 -190296.41129912098
L29_97 V29 V97 7.911057439361606e-12
C29_97 V29 V97 -6.751762424718959e-21

R29_98 V29 V98 746900.3234291644
L29_98 V29 V98 7.161150772789266e-12
C29_98 V29 V98 1.1947160603588609e-20

R29_99 V29 V99 -104394.42957571725
L29_99 V29 V99 3.2312345229546135e-11
C29_99 V29 V99 -9.96101485944448e-22

R29_100 V29 V100 -42622359.06864902
L29_100 V29 V100 7.432571655045561e-11
C29_100 V29 V100 -3.0184941814192256e-21

R29_101 V29 V101 153171.20729443515
L29_101 V29 V101 5.235552091832545e-12
C29_101 V29 V101 1.7237817906862865e-20

R29_102 V29 V102 102996.81856815857
L29_102 V29 V102 1.655840055111904e-11
C29_102 V29 V102 2.2737539269506198e-20

R29_103 V29 V103 275067.23250776326
L29_103 V29 V103 1.1744882200784458e-11
C29_103 V29 V103 9.797028484856494e-21

R29_104 V29 V104 -213681.4616891338
L29_104 V29 V104 -3.718727620869364e-11
C29_104 V29 V104 -7.710211280923707e-21

R29_105 V29 V105 -5617050.747678003
L29_105 V29 V105 4.2558245922380804e-11
C29_105 V29 V105 -2.519532301581979e-20

R29_106 V29 V106 94840.02213203312
L29_106 V29 V106 -6.620559827936925e-12
C29_106 V29 V106 2.4457227350491785e-20

R29_107 V29 V107 -648670.4046001319
L29_107 V29 V107 -1.5889820557060075e-11
C29_107 V29 V107 8.87243903677286e-21

R29_108 V29 V108 -124666.15011172679
L29_108 V29 V108 -1.6661894299212914e-11
C29_108 V29 V108 -2.505418702829376e-20

R29_109 V29 V109 -126183.99588273192
L29_109 V29 V109 8.542513401277872e-10
C29_109 V29 V109 -1.2235645615358986e-20

R29_110 V29 V110 6760691.364714162
L29_110 V29 V110 -2.4852501173106322e-11
C29_110 V29 V110 -2.7568435115025095e-20

R29_111 V29 V111 -254032.47492720227
L29_111 V29 V111 6.494208866804564e-12
C29_111 V29 V111 -3.7557339673200795e-21

R29_112 V29 V112 74554.70310956401
L29_112 V29 V112 4.805532905652063e-12
C29_112 V29 V112 1.095027895728544e-20

R29_113 V29 V113 82922.22825483137
L29_113 V29 V113 1.0309174975972986e-11
C29_113 V29 V113 5.263830483522292e-21

R29_114 V29 V114 843802.942282072
L29_114 V29 V114 -6.181457426287842e-11
C29_114 V29 V114 8.36500646646644e-21

R29_115 V29 V115 -760869.1306779403
L29_115 V29 V115 -1.1728214335621292e-11
C29_115 V29 V115 -3.392841331595837e-21

R29_116 V29 V116 -87907.96838236137
L29_116 V29 V116 -9.56942942344837e-12
C29_116 V29 V116 -1.9787317320047642e-20

R29_117 V29 V117 -113063.84910870627
L29_117 V29 V117 -8.383108364731732e-12
C29_117 V29 V117 -1.292455719836529e-20

R29_118 V29 V118 -1043900.2877333814
L29_118 V29 V118 -2.283849911280579e-11
C29_118 V29 V118 -1.6334862738988385e-20

R29_119 V29 V119 -469099.54866539664
L29_119 V29 V119 1.2834296513324999e-11
C29_119 V29 V119 -1.4117224091751193e-20

R29_120 V29 V120 58585.99653629734
L29_120 V29 V120 -6.916901194165034e-12
C29_120 V29 V120 3.925263913349637e-21

R29_121 V29 V121 155108.8514151246
L29_121 V29 V121 4.304374272626926e-12
C29_121 V29 V121 6.560478344921583e-21

R29_122 V29 V122 37197.13006852789
L29_122 V29 V122 5.76452995413114e-12
C29_122 V29 V122 -9.968453501276102e-21

R29_123 V29 V123 1522669.5961870288
L29_123 V29 V123 1.9545863660802137e-11
C29_123 V29 V123 -2.14765461339678e-21

R29_124 V29 V124 -324254.38701615937
L29_124 V29 V124 1.9894469320059195e-11
C29_124 V29 V124 6.325670816654157e-21

R29_125 V29 V125 -164961.66177958748
L29_125 V29 V125 -2.816237709108977e-12
C29_125 V29 V125 -1.0033300197787522e-20

R29_126 V29 V126 -28506.71851864123
L29_126 V29 V126 -1.5541846875362124e-11
C29_126 V29 V126 3.7369330067150925e-21

R29_127 V29 V127 32921.77053785623
L29_127 V29 V127 -1.2400105123412727e-11
C29_127 V29 V127 5.36329633063994e-21

R29_128 V29 V128 157865.58727617658
L29_128 V29 V128 -1.2061883707629468e-10
C29_128 V29 V128 3.2873620495093344e-21

R29_129 V29 V129 204333.30754195226
L29_129 V29 V129 -3.214161166640647e-11
C29_129 V29 V129 4.699857927092945e-21

R29_130 V29 V130 -321948.69165343477
L29_130 V29 V130 -3.0736875320446636e-11
C29_130 V29 V130 -6.522175033911997e-22

R29_131 V29 V131 -156617.5784288194
L29_131 V29 V131 -1.3930496468922488e-11
C29_131 V29 V131 2.555567762626849e-21

R29_132 V29 V132 -154040.8831438489
L29_132 V29 V132 -1.3984842535483407e-10
C29_132 V29 V132 -8.248198432299198e-22

R29_133 V29 V133 265799.4989603004
L29_133 V29 V133 -7.122669517434208e-12
C29_133 V29 V133 8.483832971411672e-21

R29_134 V29 V134 177209.98991111544
L29_134 V29 V134 -1.2389664698318441e-11
C29_134 V29 V134 5.586548087836971e-21

R29_135 V29 V135 53738.2082771515
L29_135 V29 V135 -1.5290563171639425e-10
C29_135 V29 V135 1.1283175710388914e-21

R29_136 V29 V136 716850.4783684717
L29_136 V29 V136 -1.0372941232179653e-10
C29_136 V29 V136 2.822326938208176e-21

R29_137 V29 V137 -171962.58938548208
L29_137 V29 V137 -7.915744416774369e-12
C29_137 V29 V137 8.530913507779522e-21

R29_138 V29 V138 -40407.46006169601
L29_138 V29 V138 -1.873984762424945e-11
C29_138 V29 V138 1.6748882524064688e-20

R29_139 V29 V139 39277.49186868403
L29_139 V29 V139 -1.1133249544008498e-11
C29_139 V29 V139 -8.820421497853466e-21

R29_140 V29 V140 -1138028.3475090142
L29_140 V29 V140 -9.825488282901178e-12
C29_140 V29 V140 -1.0625950451298004e-20

R29_141 V29 V141 -131374.08173308207
L29_141 V29 V141 -1.5838769557953667e-11
C29_141 V29 V141 5.730676321774288e-21

R29_142 V29 V142 -559279.6537338553
L29_142 V29 V142 -3.766746285901172e-11
C29_142 V29 V142 -1.3880681819523538e-20

R29_143 V29 V143 -88911.58994334718
L29_143 V29 V143 2.1978721225822307e-11
C29_143 V29 V143 -8.141003319216494e-22

R29_144 V29 V144 103075.41538357586
L29_144 V29 V144 3.2961525617835006e-11
C29_144 V29 V144 9.873999594273004e-21

R30_30 V30 0 -2239.4355677579515
L30_30 V30 0 2.7461592472480372e-12
C30_30 V30 0 -4.1626588490526315e-19

R30_31 V30 V31 234213.87015574198
L30_31 V30 V31 1.0974328790053119e-11
C30_31 V30 V31 -1.2691390532253241e-20

R30_32 V30 V32 -267666.99346514593
L30_32 V30 V32 1.0232981829777816e-11
C30_32 V30 V32 1.2604880393984427e-22

R30_33 V30 V33 38926.90041169201
L30_33 V30 V33 -5.389307236203341e-11
C30_33 V30 V33 1.915046598626771e-20

R30_34 V30 V34 -899795.8021795063
L30_34 V30 V34 3.640623242242818e-11
C30_34 V30 V34 -2.7343706027660508e-21

R30_35 V30 V35 153396.39099313034
L30_35 V30 V35 -9.068365601755097e-11
C30_35 V30 V35 1.2468540286050997e-20

R30_36 V30 V36 -74941.81433291746
L30_36 V30 V36 -2.2539160843847782e-11
C30_36 V30 V36 -2.691984870437019e-22

R30_37 V30 V37 -33764.40724703808
L30_37 V30 V37 -3.367320285362834e-11
C30_37 V30 V37 -6.763396738381252e-20

R30_38 V30 V38 -35928.44914636568
L30_38 V30 V38 -4.1173726128939675e-12
C30_38 V30 V38 -3.9159769062147334e-20

R30_39 V30 V39 -29438.440686721653
L30_39 V30 V39 -4.3672002295702776e-11
C30_39 V30 V39 -5.86559121137114e-20

R30_40 V30 V40 -2953334.525209466
L30_40 V30 V40 1.3586130962654014e-11
C30_40 V30 V40 -4.914081378664237e-21

R30_41 V30 V41 13281.727562560141
L30_41 V30 V41 -3.9037388377253386e-11
C30_41 V30 V41 1.6051324027992535e-19

R30_42 V30 V42 5030.1622284968025
L30_42 V30 V42 1.149154934995541e-12
C30_42 V30 V42 2.8774396171534793e-19

R30_43 V30 V43 -69979.74696674265
L30_43 V30 V43 -6.869400161532714e-12
C30_43 V30 V43 2.790212630944608e-20

R30_44 V30 V44 -51123.96526300838
L30_44 V30 V44 -1.1203238631935562e-11
C30_44 V30 V44 -8.839103339443825e-21

R30_45 V30 V45 -15444.927207280141
L30_45 V30 V45 -1.088427032749807e-11
C30_45 V30 V45 -1.9145241382900588e-19

R30_46 V30 V46 -170225.13841171277
L30_46 V30 V46 -5.997706521036961e-12
C30_46 V30 V46 -1.0354087214968728e-19

R30_47 V30 V47 -13526.739330416764
L30_47 V30 V47 -9.507137601436684e-12
C30_47 V30 V47 3.485981848457558e-20

R30_48 V30 V48 -20422.854382354926
L30_48 V30 V48 -8.10372523391406e-12
C30_48 V30 V48 5.229955845284342e-21

R30_49 V30 V49 45653.70555267325
L30_49 V30 V49 3.975721069095834e-11
C30_49 V30 V49 5.175329066920602e-20

R30_50 V30 V50 39653.22157519564
L30_50 V30 V50 7.603993559290392e-12
C30_50 V30 V50 3.157118394043973e-20

R30_51 V30 V51 -20193.03118687688
L30_51 V30 V51 -2.793012884506869e-12
C30_51 V30 V51 -9.213369890185121e-20

R30_52 V30 V52 15201.858934826361
L30_52 V30 V52 6.937267869075069e-12
C30_52 V30 V52 1.1251998566221422e-19

R30_53 V30 V53 -34993.728007577214
L30_53 V30 V53 -4.496335722023679e-12
C30_53 V30 V53 2.5872706513283664e-20

R30_54 V30 V54 103749.85715458743
L30_54 V30 V54 1.050056639941718e-11
C30_54 V30 V54 3.879052605569841e-20

R30_55 V30 V55 37346.33088304989
L30_55 V30 V55 1.171072083246495e-11
C30_55 V30 V55 3.8521990331298785e-20

R30_56 V30 V56 -104351.40510321918
L30_56 V30 V56 -5.998317421420035e-12
C30_56 V30 V56 1.4419676337739037e-20

R30_57 V30 V57 40357.61687740157
L30_57 V30 V57 4.098091474737367e-12
C30_57 V30 V57 -1.2362163546307306e-20

R30_58 V30 V58 4599.376234454985
L30_58 V30 V58 1.539490942475439e-12
C30_58 V30 V58 -1.7560044626368693e-20

R30_59 V30 V59 -89786.34118790735
L30_59 V30 V59 -1.9943871837792095e-11
C30_59 V30 V59 -1.901968138434187e-20

R30_60 V30 V60 -15534.240422612218
L30_60 V30 V60 -9.200408721852027e-12
C30_60 V30 V60 -1.0840727082405255e-20

R30_61 V30 V61 66145.64802290454
L30_61 V30 V61 -5.805926607263218e-12
C30_61 V30 V61 5.485072447400445e-20

R30_62 V30 V62 236859.28696440035
L30_62 V30 V62 1.9672236342492885e-11
C30_62 V30 V62 7.397671206702469e-20

R30_63 V30 V63 18065.110843523446
L30_63 V30 V63 3.688022467101884e-11
C30_63 V30 V63 -1.367982650589086e-20

R30_64 V30 V64 -298871.0559733308
L30_64 V30 V64 -6.3844297584071264e-12
C30_64 V30 V64 -1.1279648321472162e-20

R30_65 V30 V65 45905.48628968786
L30_65 V30 V65 8.42365808023087e-12
C30_65 V30 V65 2.2228954845420773e-20

R30_66 V30 V66 18813.97246968655
L30_66 V30 V66 1.2211787354783807e-11
C30_66 V30 V66 1.4660465569775485e-20

R30_67 V30 V67 -16221.566046785501
L30_67 V30 V67 -4.263161680388569e-12
C30_67 V30 V67 4.782843799005008e-21

R30_68 V30 V68 -53960.457564882614
L30_68 V30 V68 -4.566676390202886e-11
C30_68 V30 V68 7.894811265892838e-21

R30_69 V30 V69 -149604.2448081116
L30_69 V30 V69 -9.928557113322828e-12
C30_69 V30 V69 -1.1263372602269702e-20

R30_70 V30 V70 -99943.8002682812
L30_70 V30 V70 -1.2685169160239582e-11
C30_70 V30 V70 -1.3692898248351234e-20

R30_71 V30 V71 39348.564802528155
L30_71 V30 V71 1.0088840064067648e-10
C30_71 V30 V71 -1.0098274097803906e-20

R30_72 V30 V72 -99103.1302107159
L30_72 V30 V72 -4.759555456516866e-11
C30_72 V30 V72 -1.368397942860639e-21

R30_73 V30 V73 -729706.967691446
L30_73 V30 V73 -2.475208504268984e-11
C30_73 V30 V73 1.1454618667450625e-20

R30_74 V30 V74 -171127.49473864108
L30_74 V30 V74 -6.151444750536985e-12
C30_74 V30 V74 -1.1983620336123777e-20

R30_75 V30 V75 125013.83182454662
L30_75 V30 V75 9.242011998240828e-12
C30_75 V30 V75 1.9115604338141884e-20

R30_76 V30 V76 93161.73120513788
L30_76 V30 V76 -4.6007274252406866e-12
C30_76 V30 V76 -6.034348676521448e-21

R30_77 V30 V77 96686.76104821086
L30_77 V30 V77 -1.905341856093513e-11
C30_77 V30 V77 8.190647679034051e-22

R30_78 V30 V78 -29762543.753910623
L30_78 V30 V78 -1.284637521051552e-11
C30_78 V30 V78 -2.362057332969277e-21

R30_79 V30 V79 -753473.275849818
L30_79 V30 V79 -2.8605996883672427e-12
C30_79 V30 V79 -3.2327919869889095e-20

R30_80 V30 V80 107995.6016289426
L30_80 V30 V80 4.430206214703973e-12
C30_80 V30 V80 3.3927225365214525e-20

R30_81 V30 V81 -666320.1096496875
L30_81 V30 V81 1.0813849011915915e-11
C30_81 V30 V81 3.6127047348112486e-21

R30_82 V30 V82 181266.42245265679
L30_82 V30 V82 1.8423729174696238e-11
C30_82 V30 V82 3.286936364139087e-20

R30_83 V30 V83 67461.2791986384
L30_83 V30 V83 5.0544819365843426e-12
C30_83 V30 V83 3.1821160772305517e-20

R30_84 V30 V84 -213094.80350864725
L30_84 V30 V84 -5.841131687167846e-12
C30_84 V30 V84 -9.558905308252434e-21

R30_85 V30 V85 -100484.82076358383
L30_85 V30 V85 -4.4203488305831625e-12
C30_85 V30 V85 -2.3865669545077664e-20

R30_86 V30 V86 -97553.82981178259
L30_86 V30 V86 -9.028859853388992e-11
C30_86 V30 V86 -1.2166707600810585e-20

R30_87 V30 V87 -99477.39993630277
L30_87 V30 V87 -5.03808967926413e-12
C30_87 V30 V87 -2.3877293383132248e-20

R30_88 V30 V88 -437851.71458817937
L30_88 V30 V88 3.3949101916057803e-11
C30_88 V30 V88 3.075616048504375e-21

R30_89 V30 V89 220017.81684356363
L30_89 V30 V89 -8.816942748667125e-11
C30_89 V30 V89 1.6123227086198177e-20

R30_90 V30 V90 46257.25846776041
L30_90 V30 V90 2.465736343685218e-12
C30_90 V30 V90 3.2591007639164555e-20

R30_91 V30 V91 81454.41753534166
L30_91 V30 V91 1.197356013437339e-11
C30_91 V30 V91 2.5223463291935292e-20

R30_92 V30 V92 129681.70422530593
L30_92 V30 V92 2.4876037652297453e-11
C30_92 V30 V92 1.7926178725080937e-20

R30_93 V30 V93 252279.93473525517
L30_93 V30 V93 -1.1139842911509937e-11
C30_93 V30 V93 -5.9433478551137226e-21

R30_94 V30 V94 -57332.6559016524
L30_94 V30 V94 2.4012790931712355e-11
C30_94 V30 V94 -3.290186859072209e-21

R30_95 V30 V95 60504.81231121559
L30_95 V30 V95 2.092887145016254e-11
C30_95 V30 V95 1.5025780353548592e-20

R30_96 V30 V96 157657.58138744163
L30_96 V30 V96 2.3605032420542983e-11
C30_96 V30 V96 6.703412107732213e-21

R30_97 V30 V97 109539.53808272963
L30_97 V30 V97 3.892168151108144e-12
C30_97 V30 V97 1.0754022039204254e-20

R30_98 V30 V98 59462.787644390184
L30_98 V30 V98 5.983510501327025e-12
C30_98 V30 V98 2.3798912105239688e-20

R30_99 V30 V99 -39374.88771932962
L30_99 V30 V99 -5.248574513244718e-12
C30_99 V30 V99 -8.500282387995349e-21

R30_100 V30 V100 -1905242.1571750168
L30_100 V30 V100 2.4797676497400143e-11
C30_100 V30 V100 2.4514339099892428e-21

R30_101 V30 V101 944480.9609968049
L30_101 V30 V101 3.989155446209828e-11
C30_101 V30 V101 1.8273576864941975e-20

R30_102 V30 V102 23322.23942351135
L30_102 V30 V102 1.2408547119633543e-12
C30_102 V30 V102 7.653961839558823e-20

R30_103 V30 V103 -62050.04230976977
L30_103 V30 V103 -2.2206229427922333e-12
C30_103 V30 V103 -3.26623872001157e-20

R30_104 V30 V104 -266652.24008829205
L30_104 V30 V104 -2.1681609218773657e-11
C30_104 V30 V104 -2.9724207093429768e-21

R30_105 V30 V105 -97767.08996944307
L30_105 V30 V105 -3.6344674347135364e-12
C30_105 V30 V105 -2.9438759602149176e-20

R30_106 V30 V106 57686.07611436919
L30_106 V30 V106 2.3962927500051602e-12
C30_106 V30 V106 5.523423241220482e-20

R30_107 V30 V107 63243.4446058361
L30_107 V30 V107 1.4281986506433615e-12
C30_107 V30 V107 6.701521334679303e-20

R30_108 V30 V108 -152864.6462720215
L30_108 V30 V108 -1.9377137139745387e-12
C30_108 V30 V108 -5.951769777154249e-20

R30_109 V30 V109 -65665.21846351918
L30_109 V30 V109 -3.248196274543831e-12
C30_109 V30 V109 -3.186337086265933e-20

R30_110 V30 V110 47158.40391384817
L30_110 V30 V110 -8.964433370069457e-12
C30_110 V30 V110 -4.3168919105678895e-20

R30_111 V30 V111 -23720.545195388353
L30_111 V30 V111 -2.4648764196334948e-12
C30_111 V30 V111 -3.0998515292730804e-20

R30_112 V30 V112 25094.808187575974
L30_112 V30 V112 2.003655183823237e-12
C30_112 V30 V112 4.535233862296957e-20

R30_113 V30 V113 38204.135156551216
L30_113 V30 V113 4.143772896175452e-12
C30_113 V30 V113 2.1850606817800147e-20

R30_114 V30 V114 44949.147708499935
L30_114 V30 V114 4.798570367299428e-12
C30_114 V30 V114 2.157868313319494e-20

R30_115 V30 V115 30005.72633199544
L30_115 V30 V115 2.748515911728309e-12
C30_115 V30 V115 3.58300972230818e-20

R30_116 V30 V116 -40360.398534962755
L30_116 V30 V116 -3.5110472903877462e-12
C30_116 V30 V116 -3.5067162280260217e-20

R30_117 V30 V117 188451.71585572712
L30_117 V30 V117 -6.100553040740257e-12
C30_117 V30 V117 -3.0254323759697785e-20

R30_118 V30 V118 -66362.20646224408
L30_118 V30 V118 -5.110009545154678e-12
C30_118 V30 V118 -2.5470355059327075e-20

R30_119 V30 V119 -27668.853362429258
L30_119 V30 V119 -4.133794828801039e-12
C30_119 V30 V119 -2.6819196395981235e-20

R30_120 V30 V120 10292.98164304747
L30_120 V30 V120 3.3725043684329086e-12
C30_120 V30 V120 -7.709564926399781e-21

R30_121 V30 V121 -1022256.5444976554
L30_121 V30 V121 1.1969774002532558e-11
C30_121 V30 V121 5.8087044535560566e-21

R30_122 V30 V122 8774.99227364869
L30_122 V30 V122 2.239233461132405e-12
C30_122 V30 V122 -5.787360093704257e-21

R30_123 V30 V123 37492.97836414337
L30_123 V30 V123 1.0177814299453438e-11
C30_123 V30 V123 -4.836876300786814e-21

R30_124 V30 V124 -161309.25708956362
L30_124 V30 V124 -1.7193337939301214e-11
C30_124 V30 V124 -5.19773456742998e-21

R30_125 V30 V125 28810.041809066493
L30_125 V30 V125 2.1788793300350315e-11
C30_125 V30 V125 -1.0582044813911527e-20

R30_126 V30 V126 -6327.196905488674
L30_126 V30 V126 -1.7184875908920049e-12
C30_126 V30 V126 2.644546713089035e-22

R30_127 V30 V127 8190.179496415823
L30_127 V30 V127 2.023549216286794e-12
C30_127 V30 V127 3.942378971111094e-21

R30_128 V30 V128 124231.18430407673
L30_128 V30 V128 3.56303744516163e-11
C30_128 V30 V128 5.403169324874962e-22

R30_129 V30 V129 20932.908653296854
L30_129 V30 V129 5.115167087583386e-12
C30_129 V30 V129 3.0505494890523546e-21

R30_130 V30 V130 -23230.80762733394
L30_130 V30 V130 -2.817516648581308e-12
C30_130 V30 V130 -1.588080312946844e-20

R30_131 V30 V131 -26305.49607873186
L30_131 V30 V131 4.713221244971879e-10
C30_131 V30 V131 1.1536337226757149e-20

R30_132 V30 V132 -32944.74147077296
L30_132 V30 V132 -8.456428410074199e-12
C30_132 V30 V132 -6.317531237028837e-22

R30_133 V30 V133 -3614820.621521011
L30_133 V30 V133 1.3047545336575745e-11
C30_133 V30 V133 1.3799012422332848e-20

R30_134 V30 V134 -56083.95737305254
L30_134 V30 V134 -1.865090030836978e-11
C30_134 V30 V134 5.583723457421294e-21

R30_135 V30 V135 12239.157757425459
L30_135 V30 V135 3.523377082275401e-12
C30_135 V30 V135 -1.083776865788425e-20

R30_136 V30 V136 483154.1237776017
L30_136 V30 V136 7.146285028211068e-11
C30_136 V30 V136 -1.4192736889735745e-21

R30_137 V30 V137 72410.78297068244
L30_137 V30 V137 -3.244119410789875e-11
C30_137 V30 V137 -4.9068092780539756e-21

R30_138 V30 V138 -7370.49305361446
L30_138 V30 V138 -1.835586459747377e-12
C30_138 V30 V138 5.2826352983472e-21

R30_139 V30 V139 6172.066391202941
L30_139 V30 V139 1.4700922705971138e-12
C30_139 V30 V139 5.539240635837538e-21

R30_140 V30 V140 -22609.38330768265
L30_140 V30 V140 -3.668582990889301e-12
C30_140 V30 V140 -9.157488172707004e-21

R30_141 V30 V141 -30570.970239363138
L30_141 V30 V141 -6.706435162502513e-12
C30_141 V30 V141 -2.0160756825401997e-21

R30_142 V30 V142 -22189.232474007975
L30_142 V30 V142 -3.4265045154557314e-12
C30_142 V30 V142 -9.589867953255266e-21

R30_143 V30 V143 -19440.278220832075
L30_143 V30 V143 -4.992546137446755e-12
C30_143 V30 V143 -3.0185226436513212e-21

R30_144 V30 V144 48467.76700781865
L30_144 V30 V144 7.028381187646855e-12
C30_144 V30 V144 1.0680049182394217e-20

R31_31 V31 0 -677.2463739830906
L31_31 V31 0 -4.630836577809894e-13
C31_31 V31 0 -7.635512709707457e-19

R31_32 V31 V32 -150347.71433733366
L31_32 V31 V32 3.9449958420135514e-11
C31_32 V31 V32 -1.0564306725592786e-20

R31_33 V31 V33 16689.702677706126
L31_33 V31 V33 1.2483517990597067e-11
C31_33 V31 V33 2.5839435883683874e-20

R31_34 V31 V34 -62390.16178844936
L31_34 V31 V34 -5.859479100211915e-11
C31_34 V31 V34 -3.824639674032854e-21

R31_35 V31 V35 -109734.6400321361
L31_35 V31 V35 4.071794731534916e-12
C31_35 V31 V35 3.914756270893458e-20

R31_36 V31 V36 86046.15968872033
L31_36 V31 V36 -1.9813547729646308e-11
C31_36 V31 V36 -2.853524738162792e-22

R31_37 V31 V37 80208.38883151529
L31_37 V31 V37 -4.331027731773891e-12
C31_37 V31 V37 -9.096507174070752e-20

R31_38 V31 V38 -291187.12980830256
L31_38 V31 V38 6.702496633699585e-12
C31_38 V31 V38 2.3054400249954753e-20

R31_39 V31 V39 -9215.004243383115
L31_39 V31 V39 -2.560484509222458e-12
C31_39 V31 V39 -1.6562949452824915e-19

R31_40 V31 V40 -221141.91247046884
L31_40 V31 V40 1.6776544475730803e-11
C31_40 V31 V40 1.0458185320517849e-20

R31_41 V31 V41 4346.778975260577
L31_41 V31 V41 7.273002095885339e-12
C31_41 V31 V41 1.8116783443547262e-19

R31_42 V31 V42 6543.511791270724
L31_42 V31 V42 -7.343071124071814e-11
C31_42 V31 V42 1.5920496580313199e-19

R31_43 V31 V43 9841.867240044803
L31_43 V31 V43 3.368163373989162e-12
C31_43 V31 V43 1.7173636690835537e-19

R31_44 V31 V44 -103591.96279363312
L31_44 V31 V44 -2.5156067180965353e-12
C31_44 V31 V44 -1.3302300679899986e-19

R31_45 V31 V45 -81759.52607364352
L31_45 V31 V45 -1.2408736747810779e-12
C31_45 V31 V45 -3.894275801377738e-19

R31_46 V31 V46 8406.116594585053
L31_46 V31 V46 1.5644474821542143e-12
C31_46 V31 V46 1.7194833977211023e-19

R31_47 V31 V47 -124792.1185668988
L31_47 V31 V47 2.349517499742834e-12
C31_47 V31 V47 6.753389596089412e-20

R31_48 V31 V48 14675.07359020893
L31_48 V31 V48 -2.6700518094437075e-11
C31_48 V31 V48 3.915369183684737e-20

R31_49 V31 V49 8629.814343190339
L31_49 V31 V49 -3.616981308215365e-11
C31_49 V31 V49 1.379589313663367e-19

R31_50 V31 V50 -10806.665022509114
L31_50 V31 V50 6.710551111049107e-12
C31_50 V31 V50 -6.26557033746246e-20

R31_51 V31 V51 -20814.186648838873
L31_51 V31 V51 -4.007588646210346e-11
C31_51 V31 V51 -4.3424812626102735e-20

R31_52 V31 V52 90578.21694518896
L31_52 V31 V52 7.724911738550848e-12
C31_52 V31 V52 1.13771001602409e-19

R31_53 V31 V53 38942.89021070281
L31_53 V31 V53 9.138483752786475e-12
C31_53 V31 V53 5.464868473272182e-20

R31_54 V31 V54 21065.641334453663
L31_54 V31 V54 3.201707647895196e-11
C31_54 V31 V54 3.001516830306952e-20

R31_55 V31 V55 6634.993640691342
L31_55 V31 V55 6.0255190657824185e-12
C31_55 V31 V55 1.5669294219676447e-19

R31_56 V31 V56 72941.72954814375
L31_56 V31 V56 9.53369805636538e-12
C31_56 V31 V56 4.8051000854094794e-20

R31_57 V31 V57 2129.7399840796284
L31_57 V31 V57 3.914110437354869e-12
C31_57 V31 V57 -2.2723714165054136e-20

R31_58 V31 V58 6346.88027750515
L31_58 V31 V58 -7.619153305500128e-12
C31_58 V31 V58 1.6530049488919997e-22

R31_59 V31 V59 -5717.924170671477
L31_59 V31 V59 1.9119798411224885e-12
C31_59 V31 V59 -3.2999513373380715e-20

R31_60 V31 V60 7024.037421368009
L31_60 V31 V60 2.1399290685112047e-11
C31_60 V31 V60 3.2245483466640558e-21

R31_61 V31 V61 -9943.168604089162
L31_61 V31 V61 -3.528168937311123e-11
C31_61 V31 V61 7.295510148913137e-20

R31_62 V31 V62 -5901.710374315386
L31_62 V31 V62 8.99761673246018e-12
C31_62 V31 V62 5.575131641652888e-20

R31_63 V31 V63 48890.6548090538
L31_63 V31 V63 2.457015861586224e-10
C31_63 V31 V63 4.4135183916419306e-20

R31_64 V31 V64 -41449.423404387526
L31_64 V31 V64 1.1783385463135203e-11
C31_64 V31 V64 -9.993140501855125e-21

R31_65 V31 V65 5716.350501938123
L31_65 V31 V65 7.149188485040803e-12
C31_65 V31 V65 -1.497620970818684e-20

R31_66 V31 V66 4144.118152800058
L31_66 V31 V66 1.0750815703739788e-11
C31_66 V31 V66 6.747639166508188e-20

R31_67 V31 V67 85394.51609036155
L31_67 V31 V67 5.30317538367657e-12
C31_67 V31 V67 6.03619337744521e-20

R31_68 V31 V68 15784.376834895937
L31_68 V31 V68 -2.2671711291261228e-11
C31_68 V31 V68 2.8559005108956695e-21

R31_69 V31 V69 51413.48539965964
L31_69 V31 V69 -9.152967045949908e-12
C31_69 V31 V69 -2.815563598593372e-20

R31_70 V31 V70 -16466.52395934062
L31_70 V31 V70 1.8960939884764052e-10
C31_70 V31 V70 1.8107213961773287e-20

R31_71 V31 V71 34520.87692417017
L31_71 V31 V71 8.350150243207937e-11
C31_71 V31 V71 1.862959435782515e-21

R31_72 V31 V72 -11141.585641966094
L31_72 V31 V72 -1.0410603881654369e-11
C31_72 V31 V72 8.151568368817983e-21

R31_73 V31 V73 -328149.19832226576
L31_73 V31 V73 2.981713562293898e-11
C31_73 V31 V73 5.9491859419361195e-21

R31_74 V31 V74 -67675.27259556449
L31_74 V31 V74 1.6995914667813158e-11
C31_74 V31 V74 -2.2324631855316627e-20

R31_75 V31 V75 17842.626838314456
L31_75 V31 V75 5.4991099951494546e-11
C31_75 V31 V75 4.685679192304165e-21

R31_76 V31 V76 29041.631574761985
L31_76 V31 V76 9.108913995723185e-12
C31_76 V31 V76 2.872193641740813e-21

R31_77 V31 V77 66937.80557477374
L31_77 V31 V77 4.137317228064289e-11
C31_77 V31 V77 3.4954759535761985e-21

R31_78 V31 V78 137686.8675904633
L31_78 V31 V78 -4.180752445109613e-09
C31_78 V31 V78 3.4377940045177054e-20

R31_79 V31 V79 -107609.78490581845
L31_79 V31 V79 7.094140464777227e-12
C31_79 V31 V79 1.953174451305291e-21

R31_80 V31 V80 -71757.97613668175
L31_80 V31 V80 -5.588065000445004e-12
C31_80 V31 V80 1.0945349853841092e-20

R31_81 V31 V81 -94441.85807133593
L31_81 V31 V81 1.1545497470518496e-11
C31_81 V31 V81 -1.3270292248052825e-20

R31_82 V31 V82 -126690.39897710316
L31_82 V31 V82 3.0890443065253867e-12
C31_82 V31 V82 -1.0262146208550718e-20

R31_83 V31 V83 150229.89332780708
L31_83 V31 V83 6.985950266916288e-12
C31_83 V31 V83 -7.670515347074252e-21

R31_84 V31 V84 -74688.39680808887
L31_84 V31 V84 8.556046785871324e-12
C31_84 V31 V84 5.194955887356842e-22

R31_85 V31 V85 -57366.82494348403
L31_85 V31 V85 1.851419436849713e-11
C31_85 V31 V85 4.518536296988092e-22

R31_86 V31 V86 -238694.9428759523
L31_86 V31 V86 -6.767173313581188e-12
C31_86 V31 V86 -5.095903806317752e-22

R31_87 V31 V87 72000.65377148842
L31_87 V31 V87 -1.8744089417102512e-11
C31_87 V31 V87 -3.0393077208190662e-21

R31_88 V31 V88 -138130.91260445683
L31_88 V31 V88 -2.3285409805859852e-11
C31_88 V31 V88 1.5447076615915766e-21

R31_89 V31 V89 88770.88034245178
L31_89 V31 V89 -5.3795913059151663e-11
C31_89 V31 V89 1.1771433539455588e-20

R31_90 V31 V90 107743.02950144581
L31_90 V31 V90 -4.842055844108678e-12
C31_90 V31 V90 -7.176788051338148e-21

R31_91 V31 V91 -108739.5280895551
L31_91 V31 V91 2.6999089772627192e-12
C31_91 V31 V91 -9.147841524433764e-21

R31_92 V31 V92 322446.2455792067
L31_92 V31 V92 1.4222173122701416e-10
C31_92 V31 V92 4.570432502203001e-21

R31_93 V31 V93 -20757.15928320952
L31_93 V31 V93 -5.918812559222754e-10
C31_93 V31 V93 6.446512144249096e-21

R31_94 V31 V94 -30352.351245241112
L31_94 V31 V94 -1.470844496118981e-11
C31_94 V31 V94 -1.626405477894528e-21

R31_95 V31 V95 -175735.95770856406
L31_95 V31 V95 5.638007549548972e-12
C31_95 V31 V95 -4.764931788189694e-21

R31_96 V31 V96 314318.0197543303
L31_96 V31 V96 -7.299656379017081e-12
C31_96 V31 V96 1.523256904178313e-20

R31_97 V31 V97 356736.55996845214
L31_97 V31 V97 -4.092088497197696e-12
C31_97 V31 V97 3.726503117421267e-21

R31_98 V31 V98 48391.886165276796
L31_98 V31 V98 -2.7177332965556576e-11
C31_98 V31 V98 6.391361659431262e-21

R31_99 V31 V99 -55009.41809088717
L31_99 V31 V99 1.3711033590913483e-11
C31_99 V31 V99 -4.116241373982278e-21

R31_100 V31 V100 879620.6941634978
L31_100 V31 V100 -7.334919170982276e-11
C31_100 V31 V100 1.2485955844969662e-21

R31_101 V31 V101 -104016.16188739626
L31_101 V31 V101 5.7694205041343515e-11
C31_101 V31 V101 1.1860414389259697e-20

R31_102 V31 V102 242087.765598022
L31_102 V31 V102 -3.290762552318113e-12
C31_102 V31 V102 -8.166386262863106e-21

R31_103 V31 V103 1289204.6867623993
L31_103 V31 V103 5.060726925629105e-12
C31_103 V31 V103 6.878979592366106e-21

R31_104 V31 V104 -300874.95762474195
L31_104 V31 V104 -6.0531667634801936e-12
C31_104 V31 V104 2.865926562245853e-21

R31_105 V31 V105 87242.74984718833
L31_105 V31 V105 -3.621060272154682e-11
C31_105 V31 V105 5.8860917555390106e-21

R31_106 V31 V106 -75277.7976832654
L31_106 V31 V106 4.802133294222227e-12
C31_106 V31 V106 -3.0732861904518178e-21

R31_107 V31 V107 -451185.0153793596
L31_107 V31 V107 -4.646624401139266e-12
C31_107 V31 V107 -2.9877772533767427e-21

R31_108 V31 V108 47221.36911637509
L31_108 V31 V108 4.7827040090781445e-12
C31_108 V31 V108 -1.0982902857524414e-20

R31_109 V31 V109 76645.91551832341
L31_109 V31 V109 5.473101102157148e-10
C31_109 V31 V109 -3.429380965304984e-21

R31_110 V31 V110 50610.742755581414
L31_110 V31 V110 -4.8376091664209584e-12
C31_110 V31 V110 -6.371210804774589e-22

R31_111 V31 V111 69992.13939569733
L31_111 V31 V111 1.6556353105537706e-11
C31_111 V31 V111 2.507683708569339e-21

R31_112 V31 V112 18340.49958332575
L31_112 V31 V112 -5.217582905457347e-12
C31_112 V31 V112 6.69924500221316e-21

R31_113 V31 V113 34410.187589183144
L31_113 V31 V113 -3.1911554332409284e-11
C31_113 V31 V113 2.1009267453819766e-21

R31_114 V31 V114 -253915.1879154117
L31_114 V31 V114 2.065472717297492e-11
C31_114 V31 V114 4.9851892732735416e-21

R31_115 V31 V115 -291979.6273552763
L31_115 V31 V115 -1.0518168719766286e-11
C31_115 V31 V115 -7.241642464510281e-21

R31_116 V31 V116 -81322.86833356606
L31_116 V31 V116 8.540290406248844e-12
C31_116 V31 V116 -6.136837020065655e-22

R31_117 V31 V117 -108255.32858119057
L31_117 V31 V117 4.319300060439454e-11
C31_117 V31 V117 2.120033426510267e-21

R31_118 V31 V118 -32904337.711664047
L31_118 V31 V118 -1.1296774695402532e-11
C31_118 V31 V118 -8.633256889973424e-22

R31_119 V31 V119 36378.837712638284
L31_119 V31 V119 -1.6025530616061218e-11
C31_119 V31 V119 -2.6762118494751225e-22

R31_120 V31 V120 -118229.97536923303
L31_120 V31 V120 -1.8861423134371265e-11
C31_120 V31 V120 -4.099833338400129e-21

R31_121 V31 V121 14743.049594242553
L31_121 V31 V121 -1.757827339475626e-11
C31_121 V31 V121 -8.811528842520897e-21

R31_122 V31 V122 8112.234490284131
L31_122 V31 V122 -3.923935718222947e-12
C31_122 V31 V122 -2.7662051016116063e-22

R31_123 V31 V123 105806.66740451475
L31_123 V31 V123 -1.1634132732509567e-11
C31_123 V31 V123 4.35309171088035e-21

R31_124 V31 V124 193702.19312611734
L31_124 V31 V124 -1.7453258060274033e-10
C31_124 V31 V124 -1.9515941954294626e-22

R31_125 V31 V125 -13450.666482774308
L31_125 V31 V125 1.6935920251878218e-11
C31_125 V31 V125 -2.1492465984276898e-21

R31_126 V31 V126 -10017.75410592847
L31_126 V31 V126 3.912423073975181e-12
C31_126 V31 V126 1.1974808864259857e-21

R31_127 V31 V127 19172.025021137033
L31_127 V31 V127 -6.368610006816272e-12
C31_127 V31 V127 2.6453325871076026e-22

R31_128 V31 V128 -581173.5814737482
L31_128 V31 V128 1.2719985968899313e-10
C31_128 V31 V128 4.002156092426721e-21

R31_129 V31 V129 90563.76563479204
L31_129 V31 V129 -1.471408545987105e-11
C31_129 V31 V129 3.2096704505392096e-21

R31_130 V31 V130 -97539.64328962982
L31_130 V31 V130 6.012443720567078e-12
C31_130 V31 V130 -4.771563571947427e-21

R31_131 V31 V131 -35710.10020673438
L31_131 V31 V131 2.5953457039833868e-11
C31_131 V31 V131 -5.797231217166874e-21

R31_132 V31 V132 -54094.55966520116
L31_132 V31 V132 8.856491298602722e-12
C31_132 V31 V132 6.586513505343531e-22

R31_133 V31 V133 -59780.555873695506
L31_133 V31 V133 7.036996376780072e-12
C31_133 V31 V133 5.4093391406949534e-21

R31_134 V31 V134 -163677.70873274902
L31_134 V31 V134 1.3978669813760199e-11
C31_134 V31 V134 -1.976782805815592e-21

R31_135 V31 V135 24666.48906290097
L31_135 V31 V135 -8.922691395685441e-12
C31_135 V31 V135 -1.040599088817814e-23

R31_136 V31 V136 -146983.21768768318
L31_136 V31 V136 -5.420777010371411e-11
C31_136 V31 V136 -4.017001333674164e-21

R31_137 V31 V137 -21061.243669839056
L31_137 V31 V137 7.579149206312157e-11
C31_137 V31 V137 -6.636966313504474e-21

R31_138 V31 V138 -11404.052740542342
L31_138 V31 V138 3.1361549951636977e-12
C31_138 V31 V138 7.327739784136988e-21

R31_139 V31 V139 18848.94192724134
L31_139 V31 V139 -4.2647554625354095e-12
C31_139 V31 V139 -9.40575967321806e-22

R31_140 V31 V140 -57708.774604985294
L31_140 V31 V140 1.0610221723852557e-11
C31_140 V31 V140 -6.1517691502457265e-21

R31_141 V31 V141 -34809.67602848026
L31_141 V31 V141 2.2438922488991034e-11
C31_141 V31 V141 -1.1991166179981222e-21

R31_142 V31 V142 -778983.5328123191
L31_142 V31 V142 7.788753078102675e-12
C31_142 V31 V142 8.045157623645257e-21

R31_143 V31 V143 -74055.0435505763
L31_143 V31 V143 1.097985691703291e-11
C31_143 V31 V143 4.313490740752235e-21

R31_144 V31 V144 32539.04132785272
L31_144 V31 V144 -1.7299348304430505e-11
C31_144 V31 V144 7.966575937567916e-21

R32_32 V32 0 -1105.2358881112461
L32_32 V32 0 -5.223414870202502e-13
C32_32 V32 0 -4.982657575370658e-19

R32_33 V32 V33 38698.978543209276
L32_33 V32 V33 9.807398748991883e-11
C32_33 V32 V33 1.1310943632338316e-20

R32_34 V32 V34 -122510.46635220794
L32_34 V32 V34 -7.98621655852453e-11
C32_34 V32 V34 -1.9030028251393264e-21

R32_35 V32 V35 187333.74971116602
L32_35 V32 V35 -2.1621464105712045e-11
C32_35 V32 V35 1.3597996814844536e-20

R32_36 V32 V36 20319.048430313196
L32_36 V32 V36 8.211083588706447e-12
C32_36 V32 V36 9.799073684555515e-21

R32_37 V32 V37 -43327.53916506156
L32_37 V32 V37 -1.8701839923592364e-11
C32_37 V32 V37 -4.3334671204410215e-20

R32_38 V32 V38 109667.64371153597
L32_38 V32 V38 1.529642148930149e-11
C32_38 V32 V38 1.6545253954669153e-20

R32_39 V32 V39 -65193.60850907545
L32_39 V32 V39 -5.622463633402293e-11
C32_39 V32 V39 -3.504088397721702e-20

R32_40 V32 V40 -18091.924654660103
L32_40 V32 V40 -1.985614019313521e-12
C32_40 V32 V40 -1.206827407941505e-19

R32_41 V32 V41 10309.756520203753
L32_41 V32 V41 3.3261306028966133e-12
C32_41 V32 V41 1.5004359574102194e-19

R32_42 V32 V42 46438.53864185797
L32_42 V32 V42 -4.284822783695625e-11
C32_42 V32 V42 7.517693314315971e-20

R32_43 V32 V43 26802.428264325816
L32_43 V32 V43 1.3685428954925131e-11
C32_43 V32 V43 5.93143627032448e-20

R32_44 V32 V44 6043.08130947077
L32_44 V32 V44 1.1191647183754273e-12
C32_44 V32 V44 2.017315189781762e-19

R32_45 V32 V45 -11494.229515924335
L32_45 V32 V45 -2.6424983852743457e-12
C32_45 V32 V45 -1.8777578078526097e-19

R32_46 V32 V46 98853.16483291936
L32_46 V32 V46 3.897415373442395e-12
C32_46 V32 V46 2.6183921049740386e-20

R32_47 V32 V47 21035.086361023066
L32_47 V32 V47 9.745177035431197e-12
C32_47 V32 V47 -1.0534787697577256e-20

R32_48 V32 V48 15779.303473494907
L32_48 V32 V48 7.561778220155852e-12
C32_48 V32 V48 -5.291584587585839e-20

R32_49 V32 V49 100882.39016250632
L32_49 V32 V49 -3.9997927267033553e-10
C32_49 V32 V49 4.5286381415129e-20

R32_50 V32 V50 107879.33234662579
L32_50 V32 V50 1.804600848259368e-11
C32_50 V32 V50 1.339819855783472e-20

R32_51 V32 V51 124625.37742699868
L32_51 V32 V51 2.4814613344115684e-11
C32_51 V32 V51 -1.4806561150163232e-20

R32_52 V32 V52 268359.0183195676
L32_52 V32 V52 1.0232638126028785e-11
C32_52 V32 V52 9.219241258433568e-20

R32_53 V32 V53 42326.11496472192
L32_53 V32 V53 -8.390148360894744e-11
C32_53 V32 V53 -1.653193881208386e-20

R32_54 V32 V54 102513.6928567462
L32_54 V32 V54 -6.658217569933508e-11
C32_54 V32 V54 -1.5364249585151276e-20

R32_55 V32 V55 156513.14257878537
L32_55 V32 V55 1.3251571786319138e-11
C32_55 V32 V55 2.926247354861319e-20

R32_56 V32 V56 285580.5154429179
L32_56 V32 V56 5.0282064042548745e-12
C32_56 V32 V56 1.24784260932734e-19

R32_57 V32 V57 15382.601520892851
L32_57 V32 V57 5.8450772332139935e-12
C32_57 V32 V57 -5.5217198863131245e-21

R32_58 V32 V58 -17411.43603549072
L32_58 V32 V58 -4.732342165775092e-12
C32_58 V32 V58 -1.3265713609262079e-20

R32_59 V32 V59 92590.25024389864
L32_59 V32 V59 -3.374657084332211e-10
C32_59 V32 V59 -1.2058338895872612e-20

R32_60 V32 V60 3284.130351833501
L32_60 V32 V60 1.272507696461516e-12
C32_60 V32 V60 -8.824277443077825e-21

R32_61 V32 V61 -78283.65232264785
L32_61 V32 V61 -1.3011157377918812e-11
C32_61 V32 V61 3.4731617433014244e-20

R32_62 V32 V62 17253.874037565987
L32_62 V32 V62 1.0533368012731879e-11
C32_62 V32 V62 3.8167536030198954e-20

R32_63 V32 V63 190218.25102222513
L32_63 V32 V63 1.169190562525761e-11
C32_63 V32 V63 2.830109465400757e-20

R32_64 V32 V64 120950.52800356742
L32_64 V32 V64 1.8445721711250103e-11
C32_64 V32 V64 5.813647957313433e-20

R32_65 V32 V65 25426.972631277105
L32_65 V32 V65 1.6212879579658623e-11
C32_65 V32 V65 1.099592274120939e-20

R32_66 V32 V66 169342.27277293443
L32_66 V32 V66 -2.841065919247657e-11
C32_66 V32 V66 1.5240178772295805e-20

R32_67 V32 V67 35065.62093949705
L32_67 V32 V67 9.650051684421227e-12
C32_67 V32 V67 2.215566306953831e-20

R32_68 V32 V68 9394.87785993857
L32_68 V32 V68 3.061204132386726e-12
C32_68 V32 V68 1.4505686005156993e-20

R32_69 V32 V69 -19376.030654962302
L32_69 V32 V69 -5.862229660454392e-12
C32_69 V32 V69 -1.3586568228485683e-20

R32_70 V32 V70 55163.96370448885
L32_70 V32 V70 -2.3245017391171243e-11
C32_70 V32 V70 -1.2756820584497042e-20

R32_71 V32 V71 -1454190.6497142687
L32_71 V32 V71 6.903952099002212e-11
C32_71 V32 V71 4.1829118983499073e-22

R32_72 V32 V72 -104936.68604911078
L32_72 V32 V72 -3.43211485691045e-11
C32_72 V32 V72 -3.66305582341869e-21

R32_73 V32 V73 34946.540092420786
L32_73 V32 V73 -4.220107759927269e-11
C32_73 V32 V73 -4.01538855470614e-21

R32_74 V32 V74 -102751.63428060434
L32_74 V32 V74 -4.561674027600934e-11
C32_74 V32 V74 -8.746111887169062e-21

R32_75 V32 V75 5299749.748942424
L32_75 V32 V75 5.786293788101585e-11
C32_75 V32 V75 1.848501614309313e-20

R32_76 V32 V76 -217774.96571894197
L32_76 V32 V76 -4.141084922183272e-11
C32_76 V32 V76 -2.727244479803449e-21

R32_77 V32 V77 -192443.69052965965
L32_77 V32 V77 1.1722539258858298e-11
C32_77 V32 V77 6.254679173143696e-21

R32_78 V32 V78 -168726.32391670175
L32_78 V32 V78 -1.0661833341566969e-10
C32_78 V32 V78 -9.59767582235399e-21

R32_79 V32 V79 -585962.4222894075
L32_79 V32 V79 -2.772461906794509e-10
C32_79 V32 V79 -6.359074165705269e-21

R32_80 V32 V80 93647.35578638664
L32_80 V32 V80 4.916159026358753e-12
C32_80 V32 V80 4.238505923575161e-20

R32_81 V32 V81 -60860.65713772832
L32_81 V32 V81 -2.038385146879801e-12
C32_81 V32 V81 -6.778940357032276e-20

R32_82 V32 V82 75872.48836331106
L32_82 V32 V82 1.0390359495626003e-11
C32_82 V32 V82 4.533846429032276e-20

R32_83 V32 V83 54487.41408793054
L32_83 V32 V83 3.95467291548546e-12
C32_83 V32 V83 6.017768022362444e-20

R32_84 V32 V84 -384537.5404173457
L32_84 V32 V84 1.189113507234971e-11
C32_84 V32 V84 4.653229204461226e-21

R32_85 V32 V85 -421522.27954259154
L32_85 V32 V85 -1.621128289051528e-11
C32_85 V32 V85 -1.6471967394163006e-20

R32_86 V32 V86 159700.707750512
L32_86 V32 V86 -3.527039594845293e-11
C32_86 V32 V86 -3.726724142507433e-21

R32_87 V32 V87 -70808.01184911467
L32_87 V32 V87 -1.0076318681519094e-11
C32_87 V32 V87 -3.367136984620722e-20

R32_88 V32 V88 -93185.63635243678
L32_88 V32 V88 -8.497954280195939e-12
C32_88 V32 V88 -2.1701438300013867e-20

R32_89 V32 V89 134981.91813530843
L32_89 V32 V89 1.3456981093710624e-11
C32_89 V32 V89 2.8014036185226414e-20

R32_90 V32 V90 441479.875228644
L32_90 V32 V90 -1.496172968968571e-11
C32_90 V32 V90 3.0052460079431217e-21

R32_91 V32 V91 127325.59991709594
L32_91 V32 V91 -3.124676600350739e-11
C32_91 V32 V91 2.5146605656475646e-20

R32_92 V32 V92 37225.10367580149
L32_92 V32 V92 2.316303878197001e-12
C32_92 V32 V92 8.534968057702247e-20

R32_93 V32 V93 -384280.5636858739
L32_93 V32 V93 -2.3434168671000113e-11
C32_93 V32 V93 -8.073682631305967e-21

R32_94 V32 V94 -63497.94364142523
L32_94 V32 V94 -5.269235972809239e-12
C32_94 V32 V94 -4.244643896104521e-20

R32_95 V32 V95 181586.35122089574
L32_95 V32 V95 2.2405062713858018e-11
C32_95 V32 V95 2.031253345778033e-20

R32_96 V32 V96 46028.44077999984
L32_96 V32 V96 1.9881163680753505e-12
C32_96 V32 V96 7.752102429111473e-20

R32_97 V32 V97 -111222.28603556826
L32_97 V32 V97 -4.766229328533989e-12
C32_97 V32 V97 -2.7230638371049096e-20

R32_98 V32 V98 123758.26190440565
L32_98 V32 V98 7.27870232140893e-12
C32_98 V32 V98 3.7530499718329386e-20

R32_99 V32 V99 -148958.3064598652
L32_99 V32 V99 -3.983126426691041e-11
C32_99 V32 V99 -1.2296403260363226e-20

R32_100 V32 V100 -62749.322542203474
L32_100 V32 V100 -5.476345111206745e-12
C32_100 V32 V100 -3.181324074957569e-20

R32_101 V32 V101 65192.62137187692
L32_101 V32 V101 6.210256410720698e-12
C32_101 V32 V101 3.913891580031056e-20

R32_102 V32 V102 -571819.0377357663
L32_102 V32 V102 -1.4032621005460482e-11
C32_102 V32 V102 1.231265693488152e-20

R32_103 V32 V103 -4059979.624982065
L32_103 V32 V103 5.417122456956572e-11
C32_103 V32 V103 2.534023679243233e-21

R32_104 V32 V104 49758.497242978236
L32_104 V32 V104 3.0240971511732672e-12
C32_104 V32 V104 5.1417731567660766e-20

R32_105 V32 V105 -47349.388317644996
L32_105 V32 V105 -5.896544598374769e-12
C32_105 V32 V105 -5.18400140171789e-20

R32_106 V32 V106 47694.85970301921
L32_106 V32 V106 5.934699342935417e-12
C32_106 V32 V106 6.232925244553066e-20

R32_107 V32 V107 434588.6643205142
L32_107 V32 V107 -4.097833352669128e-11
C32_107 V32 V107 1.4240977864449163e-20

R32_108 V32 V108 -42194.34388052657
L32_108 V32 V108 -6.347491024307931e-12
C32_108 V32 V108 -4.839135995318971e-20

R32_109 V32 V109 44906.058206943104
L32_109 V32 V109 3.4320373303127937e-12
C32_109 V32 V109 4.93277886822208e-20

R32_110 V32 V110 -56675.61204124184
L32_110 V32 V110 -4.92189388007928e-12
C32_110 V32 V110 -5.651320915622969e-20

R32_111 V32 V111 -112158.17512161589
L32_111 V32 V111 -1.2801012914623925e-11
C32_111 V32 V111 -2.6164807295126606e-20

R32_112 V32 V112 120852.05983498294
L32_112 V32 V112 2.0009743954974722e-11
C32_112 V32 V112 3.1850732292834346e-20

R32_113 V32 V113 -117207.17038084463
L32_113 V32 V113 -9.357422401820974e-12
C32_113 V32 V113 -1.3555814788433466e-20

R32_114 V32 V114 402257.0634609164
L32_114 V32 V114 1.0695583852007786e-11
C32_114 V32 V114 3.755199732226838e-20

R32_115 V32 V115 -1604722.9522732755
L32_115 V32 V115 9.0280838746024e-09
C32_115 V32 V115 9.523466020846722e-21

R32_116 V32 V116 -82041.50724767226
L32_116 V32 V116 -8.434377064936308e-12
C32_116 V32 V116 -3.2961047908778483e-20

R32_117 V32 V117 299044.1041793458
L32_117 V32 V117 1.9261786647548452e-11
C32_117 V32 V117 6.095865489580261e-21

R32_118 V32 V118 1543644.9212333881
L32_118 V32 V118 2.2621677417620447e-11
C32_118 V32 V118 -7.470709876172874e-21

R32_119 V32 V119 -61890.58956824637
L32_119 V32 V119 -5.2840319602577226e-12
C32_119 V32 V119 -5.762611282138846e-20

R32_120 V32 V120 -844285.3746290075
L32_120 V32 V120 -6.054856623384948e-12
C32_120 V32 V120 -2.9121190977207544e-20

R32_121 V32 V121 -1015355.7498906408
L32_121 V32 V121 -2.9093279640778123e-11
C32_121 V32 V121 2.4396404480545585e-21

R32_122 V32 V122 -164137.66419404873
L32_122 V32 V122 -6.916839671731963e-12
C32_122 V32 V122 -7.692693696973236e-22

R32_123 V32 V123 -128336.1220156753
L32_123 V32 V123 -1.8994635553821806e-11
C32_123 V32 V123 -5.102654836563113e-21

R32_124 V32 V124 -55530.61203863228
L32_124 V32 V124 -7.382936711485542e-12
C32_124 V32 V124 -3.5559711628114954e-20

R32_125 V32 V125 443705.8979610468
L32_125 V32 V125 -5.1974813968400314e-11
C32_125 V32 V125 -4.6666385114819285e-21

R32_126 V32 V126 -339509.4445023999
L32_126 V32 V126 6.417485099696443e-12
C32_126 V32 V126 4.1521717032773764e-22

R32_127 V32 V127 -3240923.186098627
L32_127 V32 V127 -7.678754593491854e-12
C32_127 V32 V127 -9.77897869096568e-21

R32_128 V32 V128 -803286.8632421978
L32_128 V32 V128 2.6704455863887533e-11
C32_128 V32 V128 5.859058299731874e-22

R32_129 V32 V129 -76438.12826181881
L32_129 V32 V129 -9.962611554335658e-12
C32_129 V32 V129 -9.480543599066344e-21

R32_130 V32 V130 146820.6456874146
L32_130 V32 V130 1.0020214807383811e-11
C32_130 V32 V130 -4.729420247545584e-21

R32_131 V32 V131 87084.8101253671
L32_131 V32 V131 1.1425444194441685e-11
C32_131 V32 V131 6.591291193486208e-21

R32_132 V32 V132 -1652909.8557646805
L32_132 V32 V132 -1.7735089812738304e-11
C32_132 V32 V132 -7.923662586134155e-21

R32_133 V32 V133 136359.73340179338
L32_133 V32 V133 1.446651131499798e-11
C32_133 V32 V133 1.818032409293622e-20

R32_134 V32 V134 520599.359158146
L32_134 V32 V134 4.315378864338731e-11
C32_134 V32 V134 -2.3371449160117203e-21

R32_135 V32 V135 611631.6072932151
L32_135 V32 V135 -1.3799457764791488e-11
C32_135 V32 V135 -3.8389778505992144e-21

R32_136 V32 V136 417699.94641490735
L32_136 V32 V136 1.4226811518164477e-10
C32_136 V32 V136 -5.600431491045973e-21

R32_137 V32 V137 -145836.01007305307
L32_137 V32 V137 -4.7192655817406086e-11
C32_137 V32 V137 -1.809573448120974e-20

R32_138 V32 V138 136987.43740353972
L32_138 V32 V138 6.708009473293033e-12
C32_138 V32 V138 -1.1855113135976076e-20

R32_139 V32 V139 204030.96385597214
L32_139 V32 V139 -6.7697238622755495e-12
C32_139 V32 V139 1.1306312897962357e-21

R32_140 V32 V140 -168618.26214116786
L32_140 V32 V140 6.023443269231434e-11
C32_140 V32 V140 -5.978330078786067e-21

R32_141 V32 V141 -221461.13563750382
L32_141 V32 V141 -8.596137726701337e-11
C32_141 V32 V141 -2.0912768530648074e-21

R32_142 V32 V142 9275748.781922258
L32_142 V32 V142 1.383635478407061e-11
C32_142 V32 V142 -1.3403982251914027e-20

R32_143 V32 V143 -2880960.9946731655
L32_143 V32 V143 1.6072134678749572e-11
C32_143 V32 V143 -3.145429079523971e-21

R32_144 V32 V144 1228523.3369362184
L32_144 V32 V144 1.9934749122302848e-11
C32_144 V32 V144 5.30425171355282e-22

R33_33 V33 0 72.6778665758794
L33_33 V33 0 6.224772943227566e-14
C33_33 V33 0 1.6375240215721183e-18

R33_34 V33 V34 2965.048974451275
L33_34 V33 V34 3.1111204897093995e-12
C33_34 V33 V34 4.841212948093656e-20

R33_35 V33 V35 -2081.5806336120295
L33_35 V33 V35 -2.3273194345672827e-12
C33_35 V33 V35 -7.261415861888334e-20

R33_36 V33 V36 7480.65589650531
L33_36 V33 V36 8.455679954859465e-12
C33_36 V33 V36 1.160822253841362e-20

R33_37 V33 V37 5489.834398861078
L33_37 V33 V37 1.0315690243026513e-12
C33_37 V33 V37 1.6316473722478752e-19

R33_38 V33 V38 -25438.490562707804
L33_38 V33 V38 -4.1379467637145004e-11
C33_38 V33 V38 1.803038689222859e-20

R33_39 V33 V39 2930.1810686851272
L33_39 V33 V39 1.2205366584160298e-12
C33_39 V33 V39 1.5005034847371008e-19

R33_40 V33 V40 -19518.12276065673
L33_40 V33 V40 6.344576182343642e-11
C33_40 V33 V40 1.5464182458189038e-20

R33_41 V33 V41 -574.6831016529187
L33_41 V33 V41 -2.710305044367209e-13
C33_41 V33 V41 -5.161506665390357e-19

R33_42 V33 V42 -1029.7763921786252
L33_42 V33 V42 -3.933540736833115e-13
C33_42 V33 V42 -4.348236134511906e-19

R33_43 V33 V43 -2097.6427425477755
L33_43 V33 V43 -8.158784991174289e-13
C33_43 V33 V43 -1.6239565235930617e-19

R33_44 V33 V44 22339.648213595083
L33_44 V33 V44 -1.0765169806305038e-11
C33_44 V33 V44 -7.017360203637038e-20

R33_45 V33 V45 -1396.3649169268283
L33_45 V33 V45 7.427244598165516e-13
C33_45 V33 V45 2.774721429810524e-19

R33_46 V33 V46 -1119.3716093581854
L33_46 V33 V46 4.331040036005797e-12
C33_46 V33 V46 2.2230640288516192e-19

R33_47 V33 V47 -1335.869416198952
L33_47 V33 V47 -1.0431819232951174e-11
C33_47 V33 V47 6.481561374852758e-20

R33_48 V33 V48 3903.167540364774
L33_48 V33 V48 4.8907371702279185e-12
C33_48 V33 V48 3.0998935241924335e-20

R33_49 V33 V49 1697.313292602418
L33_49 V33 V49 -3.0377163711627306e-12
C33_49 V33 V49 -8.751485467998761e-20

R33_50 V33 V50 -1794.7665059199105
L33_50 V33 V50 -1.3860019356383626e-12
C33_50 V33 V50 -1.0605727110725663e-19

R33_51 V33 V51 2447.7364532442957
L33_51 V33 V51 1.641636983120994e-12
C33_51 V33 V51 8.297226312998084e-20

R33_52 V33 V52 7885.479369979831
L33_52 V33 V52 -7.229151972305563e-13
C33_52 V33 V52 -2.534940869361732e-19

R33_53 V33 V53 -21655.625360989114
L33_53 V33 V53 -1.0017100122411623e-12
C33_53 V33 V53 -1.2419718635859218e-19

R33_54 V33 V54 -1879.6333644488288
L33_54 V33 V54 -2.1168683649601837e-12
C33_54 V33 V54 -1.172259723754232e-20

R33_55 V33 V55 -1855.5496315453079
L33_55 V33 V55 -1.3092317910968369e-12
C33_55 V33 V55 -3.634986130924901e-20

R33_56 V33 V56 -2557.5790252368306
L33_56 V33 V56 -1.7633022172796827e-12
C33_56 V33 V56 -4.27747805624295e-20

R33_57 V33 V57 -180.31425859075017
L33_57 V33 V57 -3.113877270975599e-13
C33_57 V33 V57 8.858025460308748e-20

R33_58 V33 V58 -872.3616650644694
L33_58 V33 V58 -1.342573809455931e-12
C33_58 V33 V58 4.3697550204603504e-20

R33_59 V33 V59 -1798.2511403205096
L33_59 V33 V59 -1.6603319695054003e-11
C33_59 V33 V59 3.3002639058574634e-20

R33_60 V33 V60 -1283.6122373238882
L33_60 V33 V60 -1.9255034239038183e-12
C33_60 V33 V60 1.9173934204236054e-20

R33_61 V33 V61 625.0664715997376
L33_61 V33 V61 -1.0916652920680852e-09
C33_61 V33 V61 -2.26312164150244e-19

R33_62 V33 V62 699.7355513071516
L33_62 V33 V62 4.681137187813941e-12
C33_62 V33 V62 -1.963703007083193e-19

R33_63 V33 V63 6970.242953664399
L33_63 V33 V63 -9.313074178090899e-10
C33_63 V33 V63 -1.4023240589660024e-20

R33_64 V33 V64 -12873.135368277042
L33_64 V33 V64 -4.5616702117430385e-12
C33_64 V33 V64 -2.0890516423933402e-20

R33_65 V33 V65 -496.40501986296863
L33_65 V33 V65 -5.346845594222371e-13
C33_65 V33 V65 -1.1406772859009288e-19

R33_66 V33 V66 -631.1745212973865
L33_66 V33 V66 -5.489196283446669e-13
C33_66 V33 V66 -5.738654292425049e-20

R33_67 V33 V67 -2276.5521474769266
L33_67 V33 V67 -2.5494518218789838e-12
C33_67 V33 V67 -1.613597793647898e-20

R33_68 V33 V68 -8224.712556207138
L33_68 V33 V68 -4.779633666604484e-12
C33_68 V33 V68 -2.1474249975723185e-20

R33_69 V33 V69 3659.5717975769185
L33_69 V33 V69 2.73601003031872e-12
C33_69 V33 V69 1.4342537077894793e-20

R33_70 V33 V70 3632.2867047366085
L33_70 V33 V70 5.357441086580394e-12
C33_70 V33 V70 3.357917000897724e-20

R33_71 V33 V71 27430.920309428668
L33_71 V33 V71 6.614657752086014e-12
C33_71 V33 V71 1.3449254245538708e-20

R33_72 V33 V72 2900.896517079657
L33_72 V33 V72 1.9214156606868234e-12
C33_72 V33 V72 5.453512229259675e-20

R33_73 V33 V73 -21832.695079520137
L33_73 V33 V73 -7.478411322081244e-11
C33_73 V33 V73 -9.268740584394099e-21

R33_74 V33 V74 3487.7379475623334
L33_74 V33 V74 2.3369886835728027e-12
C33_74 V33 V74 3.8109221006009735e-20

R33_75 V33 V75 -3676.121435226469
L33_75 V33 V75 -2.7895137932472792e-12
C33_75 V33 V75 -4.995633820412075e-20

R33_76 V33 V76 -4129.074996066117
L33_76 V33 V76 -1.641489629049302e-12
C33_76 V33 V76 -5.365715965203082e-20

R33_77 V33 V77 -12663.838135367145
L33_77 V33 V77 -4.8355607286566925e-12
C33_77 V33 V77 -2.276623089083245e-20

R33_78 V33 V78 20095.78345274829
L33_78 V33 V78 -4.7916428626991995e-12
C33_78 V33 V78 2.0055784907200225e-21

R33_79 V33 V79 16302.080996232122
L33_79 V33 V79 4.28031160973787e-11
C33_79 V33 V79 -1.4007456004938714e-20

R33_80 V33 V80 11133.555589365766
L33_80 V33 V80 5.549781265340319e-12
C33_80 V33 V80 -1.0710991051472551e-20

R33_81 V33 V81 134338.01344844856
L33_81 V33 V81 1.305138642996718e-11
C33_81 V33 V81 9.496635436185272e-21

R33_82 V33 V82 19071.5709889699
L33_82 V33 V82 1.3107206907493397e-11
C33_82 V33 V82 -8.603322094174648e-20

R33_83 V33 V83 -26248.5612340294
L33_83 V33 V83 5.674542130303207e-12
C33_83 V33 V83 -2.449959033920416e-20

R33_84 V33 V84 -12488.289618447077
L33_84 V33 V84 2.1558036682979155e-11
C33_84 V33 V84 3.6535321902971475e-20

R33_85 V33 V85 21588.973584022893
L33_85 V33 V85 2.246187877068399e-10
C33_85 V33 V85 3.7782189830021905e-20

R33_86 V33 V86 23138.447267527627
L33_86 V33 V86 -2.2325907404620745e-11
C33_86 V33 V86 4.384310075257647e-20

R33_87 V33 V87 254747.69676752773
L33_87 V33 V87 -7.663155606100266e-12
C33_87 V33 V87 3.374080505937755e-20

R33_88 V33 V88 16221.047966374612
L33_88 V33 V88 -1.477163796972836e-11
C33_88 V33 V88 -7.936741295559149e-21

R33_89 V33 V89 -14589.180562829515
L33_89 V33 V89 -1.764700267715409e-11
C33_89 V33 V89 -9.493591403930156e-20

R33_90 V33 V90 55189.95673697543
L33_90 V33 V90 1.8841075543266012e-11
C33_90 V33 V90 3.34619109875233e-22

R33_91 V33 V91 -173710.15609999906
L33_91 V33 V91 8.926505925848747e-12
C33_91 V33 V91 -7.953707174323468e-20

R33_92 V33 V92 -81643.30139267225
L33_92 V33 V92 1.7713667722895216e-11
C33_92 V33 V92 -2.8922719421694246e-20

R33_93 V33 V93 2794.849657982805
L33_93 V33 V93 -1.189384764836425e-10
C33_93 V33 V93 -3.087963547070087e-20

R33_94 V33 V94 6471.359582996318
L33_94 V33 V94 -7.327335146069956e-11
C33_94 V33 V94 3.412498383679478e-20

R33_95 V33 V95 64029.9838937919
L33_95 V33 V95 1.48947034330836e-11
C33_95 V33 V95 -3.7565149512297166e-20

R33_96 V33 V96 -15009.429539698083
L33_96 V33 V96 3.2182140228834204e-11
C33_96 V33 V96 1.186403610829485e-20

R33_97 V33 V97 11881.842346054444
L33_97 V33 V97 -3.618342431978672e-10
C33_97 V33 V97 1.171945126162491e-20

R33_98 V33 V98 20237.877553740975
L33_98 V33 V98 1.457544065826527e-11
C33_98 V33 V98 -4.188220875747287e-20

R33_99 V33 V99 12952.835435115416
L33_99 V33 V99 -2.5691700567975195e-11
C33_99 V33 V99 1.991237764573505e-21

R33_100 V33 V100 -29801.38130535814
L33_100 V33 V100 -5.55155297646623e-11
C33_100 V33 V100 3.654281787450984e-21

R33_101 V33 V101 11677.785349487265
L33_101 V33 V101 4.300751784842902e-11
C33_101 V33 V101 -8.822229080221676e-20

R33_102 V33 V102 10618.41661717047
L33_102 V33 V102 6.840620014641906e-12
C33_102 V33 V102 -4.3526917397586114e-20

R33_103 V33 V103 27541.054860418215
L33_103 V33 V103 -1.100330922188427e-11
C33_103 V33 V103 -4.4011505204314075e-20

R33_104 V33 V104 173574.72716869295
L33_104 V33 V104 -3.9237717773440135e-11
C33_104 V33 V104 1.568325116281069e-20

R33_105 V33 V105 -9672.118066672772
L33_105 V33 V105 -8.184040185634426e-12
C33_105 V33 V105 3.136072859108614e-20

R33_106 V33 V106 -10855.20665113219
L33_106 V33 V106 4.931525351363769e-12
C33_106 V33 V106 -6.184453916446427e-20

R33_107 V33 V107 83883.61583192719
L33_107 V33 V107 6.250637253487353e-12
C33_107 V33 V107 1.7435459207172722e-20

R33_108 V33 V108 -15222.503173834379
L33_108 V33 V108 -9.985954261867243e-12
C33_108 V33 V108 5.229413804389e-20

R33_109 V33 V109 -37697.95648451304
L33_109 V33 V109 -2.063066768331559e-11
C33_109 V33 V109 2.724882979909259e-20

R33_110 V33 V110 31996.40207863062
L33_110 V33 V110 -8.101006103896037e-12
C33_110 V33 V110 6.303462119464052e-20

R33_111 V33 V111 -7400.735794774523
L33_111 V33 V111 -7.29562672303986e-12
C33_111 V33 V111 -1.0205661496878806e-20

R33_112 V33 V112 -6204.678554058241
L33_112 V33 V112 1.2167545342763239e-11
C33_112 V33 V112 -5.743288229297931e-20

R33_113 V33 V113 -7296.221305030417
L33_113 V33 V113 2.743036631561926e-11
C33_113 V33 V113 -2.6640656528122405e-20

R33_114 V33 V114 50924.44763826083
L33_114 V33 V114 8.798768722691697e-12
C33_114 V33 V114 -3.3633824608381364e-20

R33_115 V33 V115 11102.811910589757
L33_115 V33 V115 1.3088332799464005e-11
C33_115 V33 V115 5.991458003987137e-21

R33_116 V33 V116 58242.6080406773
L33_116 V33 V116 -1.3322689703638067e-11
C33_116 V33 V116 1.94495351552483e-20

R33_117 V33 V117 7216.816897815734
L33_117 V33 V117 -1.1578809908066883e-10
C33_117 V33 V117 3.9108306225366953e-20

R33_118 V33 V118 -19206.850278558406
L33_118 V33 V118 -1.0598318785805718e-11
C33_118 V33 V118 3.143482693547233e-20

R33_119 V33 V119 -5128.470781517021
L33_119 V33 V119 -8.671990090803496e-12
C33_119 V33 V119 3.7101474488793667e-20

R33_120 V33 V120 3368.8031175279566
L33_120 V33 V120 1.516117008641877e-11
C33_120 V33 V120 5.7476129794792566e-21

R33_121 V33 V121 -3453.845932048321
L33_121 V33 V121 1.1492858918015462e-10
C33_121 V33 V121 5.30093263470196e-22

R33_122 V33 V122 -3414.118092270135
L33_122 V33 V122 2.0995227554804754e-11
C33_122 V33 V122 -6.819082580321968e-21

R33_123 V33 V123 33339.39487932598
L33_123 V33 V123 2.911693455268801e-11
C33_123 V33 V123 8.78640092743096e-21

R33_124 V33 V124 124147.1851703754
L33_124 V33 V124 -8.28207031660066e-11
C33_124 V33 V124 -2.5243916086334677e-21

R33_125 V33 V125 2310.0415831733762
L33_125 V33 V125 8.964845836586997e-11
C33_125 V33 V125 -1.0690275281177819e-21

R33_126 V33 V126 9196.605691963528
L33_126 V33 V126 -1.0668418149637e-11
C33_126 V33 V126 -1.111741528095003e-20

R33_127 V33 V127 11237.430880120757
L33_127 V33 V127 9.93189337642933e-12
C33_127 V33 V127 -5.641916706095774e-21

R33_128 V33 V128 18954.80770542815
L33_128 V33 V128 5.592578165427064e-11
C33_128 V33 V128 -4.496357304642017e-22

R33_129 V33 V129 8874.296806416725
L33_129 V33 V129 1.2872645819510721e-11
C33_129 V33 V129 1.22247700993246e-20

R33_130 V33 V130 58156.558874779636
L33_130 V33 V130 -1.4318198226436263e-11
C33_130 V33 V130 1.0926946646837896e-20

R33_131 V33 V131 17075.505433802868
L33_131 V33 V131 3.6640783164303896e-10
C33_131 V33 V131 2.7544268495803966e-21

R33_132 V33 V132 -215041.98550407306
L33_132 V33 V132 -1.0214602539069042e-10
C33_132 V33 V132 -3.561404378183456e-21

R33_133 V33 V133 76341.00508908479
L33_133 V33 V133 2.5799186513156227e-11
C33_133 V33 V133 -3.869593618184052e-20

R33_134 V33 V134 -11256.929074476106
L33_134 V33 V134 -3.13830004876917e-11
C33_134 V33 V134 -1.2482387196158152e-20

R33_135 V33 V135 -117382.41211043237
L33_135 V33 V135 2.3857024236384874e-11
C33_135 V33 V135 -3.895295330797742e-21

R33_136 V33 V136 22298.66975652808
L33_136 V33 V136 -6.066108823143118e-10
C33_136 V33 V136 3.8074463424052786e-21

R33_137 V33 V137 2963.898565684639
L33_137 V33 V137 2.9846888670616925e-11
C33_137 V33 V137 2.304914485310662e-20

R33_138 V33 V138 9494.79360079531
L33_138 V33 V138 -1.2652054516148763e-11
C33_138 V33 V138 -7.58685889487084e-21

R33_139 V33 V139 5798.1164249255935
L33_139 V33 V139 6.8062319921002035e-12
C33_139 V33 V139 7.257608401815136e-21

R33_140 V33 V140 -9518.226521769848
L33_140 V33 V140 -2.6589840086721848e-11
C33_140 V33 V140 1.641969638020614e-20

R33_141 V33 V141 8754.819780716254
L33_141 V33 V141 -7.588047901041852e-11
C33_141 V33 V141 -5.0916526158060905e-21

R33_142 V33 V142 -6184.20007130281
L33_142 V33 V142 -1.7170146912463e-11
C33_142 V33 V142 1.4701460852118094e-20

R33_143 V33 V143 -14671.494601651715
L33_143 V33 V143 -1.6179451837699076e-11
C33_143 V33 V143 -1.1845319361194019e-20

R33_144 V33 V144 -6966.238014317405
L33_144 V33 V144 -9.646878522421483e-11
C33_144 V33 V144 -2.2668681738925217e-20

R34_34 V34 0 -155.76251015303035
L34_34 V34 0 -1.556123802783228e-13
C34_34 V34 0 -6.536724560149204e-19

R34_35 V34 V35 4155.921566349996
L34_35 V34 V35 5.169882545171307e-12
C34_35 V34 V35 1.9716463167467302e-20

R34_36 V34 V36 -19555.933298189502
L34_36 V34 V36 -1.8657599316003015e-11
C34_36 V34 V36 -6.075311565311023e-21

R34_37 V34 V37 -10592.912094489684
L34_37 V34 V37 -2.3003121184947584e-12
C34_37 V34 V37 -5.944244053612526e-20

R34_38 V34 V38 19926.704982452244
L34_38 V34 V38 9.266828726012485e-12
C34_38 V34 V38 1.4439987111458727e-20

R34_39 V34 V39 -5839.740786206837
L34_39 V34 V39 -2.3143542855652663e-12
C34_39 V34 V39 -6.354841198830844e-20

R34_40 V34 V40 30048.56426535234
L34_40 V34 V40 1.834405169682359e-10
C34_40 V34 V40 1.9206241332304678e-20

R34_41 V34 V41 1216.206279842737
L34_41 V34 V41 6.263396602947512e-13
C34_41 V34 V41 1.801700836805542e-19

R34_42 V34 V42 3676.9340373815485
L34_42 V34 V42 1.3818857950454665e-12
C34_42 V34 V42 5.547355998836803e-20

R34_43 V34 V43 3646.146495777524
L34_43 V34 V43 1.3610411505599644e-12
C34_43 V34 V43 8.83443538690629e-20

R34_44 V34 V44 -30801.42922076684
L34_44 V34 V44 -3.577812957235758e-11
C34_44 V34 V44 -2.263385438764634e-20

R34_45 V34 V45 2756.752958906312
L34_45 V34 V45 -1.5523233152343892e-12
C34_45 V34 V45 -7.101858235529564e-20

R34_46 V34 V46 2518.7519882884208
L34_46 V34 V46 1.657644486535378e-11
C34_46 V34 V46 -2.970921136370748e-20

R34_47 V34 V47 1794.6361742093727
L34_47 V34 V47 8.149432876757371e-12
C34_47 V34 V47 -3.6948800379972115e-20

R34_48 V34 V48 -30760.51429064262
L34_48 V34 V48 -1.8013692353608936e-11
C34_48 V34 V48 3.65824562473403e-21

R34_49 V34 V49 -3206.3171377709614
L34_49 V34 V49 9.454035011799525e-12
C34_49 V34 V49 3.2041663662385935e-20

R34_50 V34 V50 3798.3848397248826
L34_50 V34 V50 3.3714723810509447e-12
C34_50 V34 V50 1.4411764844124085e-20

R34_51 V34 V51 -5553.658882162931
L34_51 V34 V51 -7.230012871135514e-12
C34_51 V34 V51 3.1717084184536855e-20

R34_52 V34 V52 -8148.894883919062
L34_52 V34 V52 1.8355687484477747e-12
C34_52 V34 V52 7.273062198034058e-20

R34_53 V34 V53 8894.311734657518
L34_53 V34 V53 2.0420226131677223e-12
C34_53 V34 V53 5.723623388541595e-20

R34_54 V34 V54 3720.1480231011515
L34_54 V34 V54 7.285519277451722e-12
C34_54 V34 V54 -7.833839642534854e-21

R34_55 V34 V55 4281.174508270399
L34_55 V34 V55 3.213011936742637e-12
C34_55 V34 V55 2.6143805082847408e-20

R34_56 V34 V56 4663.9315141529405
L34_56 V34 V56 4.021016890848984e-12
C34_56 V34 V56 2.5830663999568292e-21

R34_57 V34 V57 381.1018044351391
L34_57 V34 V57 7.53158861651488e-13
C34_57 V34 V57 -3.60009276634227e-20

R34_58 V34 V58 7532.0982955487025
L34_58 V34 V58 -1.9587574510289166e-11
C34_58 V34 V58 3.839226632858031e-21

R34_59 V34 V59 3357.5551146883204
L34_59 V34 V59 8.69404862886243e-12
C34_59 V34 V59 1.4234880630353761e-21

R34_60 V34 V60 2254.5542738299323
L34_60 V34 V60 5.21053386663285e-12
C34_60 V34 V60 -2.350500098164163e-21

R34_61 V34 V61 -1356.0727591668874
L34_61 V34 V61 9.465704977787727e-11
C34_61 V34 V61 9.3804765496907e-20

R34_62 V34 V62 -1511.839885608607
L34_62 V34 V62 -1.587216831641462e-11
C34_62 V34 V62 5.559253428320699e-20

R34_63 V34 V63 -7555.135535674093
L34_63 V34 V63 -1.3922913281717427e-11
C34_63 V34 V63 2.256136282121965e-20

R34_64 V34 V64 17844.722028832824
L34_64 V34 V64 1.0405483100557317e-11
C34_64 V34 V64 1.1866989358544855e-20

R34_65 V34 V65 1062.8409908996
L34_65 V34 V65 1.3472545882232383e-12
C34_65 V34 V65 2.858472056173739e-20

R34_66 V34 V66 1403.8614523727701
L34_66 V34 V66 1.3978241464817225e-12
C34_66 V34 V66 4.073636198720156e-20

R34_67 V34 V67 3328.8997092826767
L34_67 V34 V67 3.455713922122403e-12
C34_67 V34 V67 3.241257979481652e-20

R34_68 V34 V68 15585.381696316284
L34_68 V34 V68 1.538661223889355e-11
C34_68 V34 V68 9.420421514521046e-21

R34_69 V34 V69 -7318.760999483705
L34_69 V34 V69 -9.417114392421035e-12
C34_69 V34 V69 2.005237126861629e-20

R34_70 V34 V70 -9719.807298409774
L34_70 V34 V70 -1.2168706275550263e-11
C34_70 V34 V70 4.5290790869346135e-21

R34_71 V34 V71 84156.39427978867
L34_71 V34 V71 -3.5160822894343e-11
C34_71 V34 V71 2.631897847819005e-21

R34_72 V34 V72 -5920.501332089174
L34_72 V34 V72 -4.209432284884929e-12
C34_72 V34 V72 -1.880617915679609e-20

R34_73 V34 V73 -350372.19742829737
L34_73 V34 V73 -4.242333843203868e-11
C34_73 V34 V73 7.894594424514133e-21

R34_74 V34 V74 -6227.24398227546
L34_74 V34 V74 -4.583916412271292e-12
C34_74 V34 V74 -4.1138483420857605e-20

R34_75 V34 V75 6946.381429100335
L34_75 V34 V75 6.301235151493243e-12
C34_75 V34 V75 -8.197158002149039e-21

R34_76 V34 V76 11035.257941300113
L34_76 V34 V76 5.1428728797292e-12
C34_76 V34 V76 1.5821413284912178e-20

R34_77 V34 V77 74995.58558522638
L34_77 V34 V77 1.77819633338477e-11
C34_77 V34 V77 -9.917643971493846e-21

R34_78 V34 V78 -44189.14666644535
L34_78 V34 V78 7.584113987906037e-12
C34_78 V34 V78 4.646082131306168e-20

R34_79 V34 V79 -20143.2318133938
L34_79 V34 V79 -1.4799126949947346e-11
C34_79 V34 V79 -3.0556312547748993e-21

R34_80 V34 V80 -26243.495146951253
L34_80 V34 V80 -2.866531121277818e-11
C34_80 V34 V80 2.0050151002691542e-21

R34_81 V34 V81 91501.66604676889
L34_81 V34 V81 -2.3589898506735443e-10
C34_81 V34 V81 2.69515666123516e-20

R34_82 V34 V82 -21593.194848607534
L34_82 V34 V82 -4.357616682897565e-11
C34_82 V34 V82 -4.8596313601795335e-21

R34_83 V34 V83 56185.655704754674
L34_83 V34 V83 -2.2021814072106092e-11
C34_83 V34 V83 -3.3777796463228904e-20

R34_84 V34 V84 75627.44742382
L34_84 V34 V84 -2.2279590771261092e-11
C34_84 V34 V84 -8.013656704094757e-21

R34_85 V34 V85 -34701.17435786033
L34_85 V34 V85 -5.521921738779743e-11
C34_85 V34 V85 1.3564967162884975e-20

R34_86 V34 V86 -35688.17527137024
L34_86 V34 V86 2.164348348031244e-09
C34_86 V34 V86 -1.5832845209070268e-21

R34_87 V34 V87 123781.72631079708
L34_87 V34 V87 3.4747326849379074e-11
C34_87 V34 V87 4.402434149952234e-21

R34_88 V34 V88 -63741.09008484065
L34_88 V34 V88 2.041354867017114e-11
C34_88 V34 V88 2.2670368352742324e-20

R34_89 V34 V89 38818.23726848818
L34_89 V34 V89 4.280999972899305e-11
C34_89 V34 V89 2.518148229073738e-20

R34_90 V34 V90 344705.2077661354
L34_90 V34 V90 8.686824672585157e-11
C34_90 V34 V90 -1.3387853315073218e-20

R34_91 V34 V91 -98787.33153561257
L34_91 V34 V91 -2.4953502265028698e-11
C34_91 V34 V91 -9.150876986664776e-21

R34_92 V34 V92 -93271.54320423702
L34_92 V34 V92 -3.967038948004211e-11
C34_92 V34 V92 -2.4575218395246405e-20

R34_93 V34 V93 -6101.034793191509
L34_93 V34 V93 4.538578052864083e-10
C34_93 V34 V93 2.1094985173788308e-20

R34_94 V34 V94 -17284.597782296423
L34_94 V34 V94 7.538859017715705e-11
C34_94 V34 V94 6.194180241822516e-21

R34_95 V34 V95 -59382.45196724221
L34_95 V34 V95 -3.3951303775619814e-11
C34_95 V34 V95 -1.1209086482458605e-20

R34_96 V34 V96 43164.483729155334
L34_96 V34 V96 -5.2114788884223685e-11
C34_96 V34 V96 -3.149953440580137e-20

R34_97 V34 V97 -28056.011627939846
L34_97 V34 V97 3.0718377854986494e-11
C34_97 V34 V97 1.7513983744952928e-20

R34_98 V34 V98 -22590.017875858703
L34_98 V34 V98 -1.067136821639993e-10
C34_98 V34 V98 -2.307617076231554e-21

R34_99 V34 V99 -23852.06916325378
L34_99 V34 V99 -6.854068472454028e-11
C34_99 V34 V99 -6.55165623859175e-21

R34_100 V34 V100 47898.82748070527
L34_100 V34 V100 1.1807808228231898e-10
C34_100 V34 V100 1.0056687726236914e-20

R34_101 V34 V101 -20760.014023297957
L34_101 V34 V101 -8.389975822281657e-11
C34_101 V34 V101 5.458381213698354e-21

R34_102 V34 V102 -18938.22981938908
L34_102 V34 V102 2.7526211957405345e-10
C34_102 V34 V102 -1.9453153605047488e-20

R34_103 V34 V103 -45160.380160584
L34_103 V34 V103 5.360882440283173e-11
C34_103 V34 V103 4.0652195639917944e-20

R34_104 V34 V104 -97644.05474321923
L34_104 V34 V104 -3.834337697387106e-11
C34_104 V34 V104 -3.1421174085702134e-20

R34_105 V34 V105 16600.009516968217
L34_105 V34 V105 2.6125056922891345e-11
C34_105 V34 V105 3.3652359827395143e-20

R34_106 V34 V106 32432.088891179854
L34_106 V34 V106 -2.1119930860459635e-11
C34_106 V34 V106 -3.335664803205744e-20

R34_107 V34 V107 -88639.52707423059
L34_107 V34 V107 7.032384025301493e-11
C34_107 V34 V107 -1.0930674766369098e-20

R34_108 V34 V108 41767.68022750162
L34_108 V34 V108 -3.557176089567593e-11
C34_108 V34 V108 -1.0571872646949863e-20

R34_109 V34 V109 -13166276.222408537
L34_109 V34 V109 -3.5187755806911224e-11
C34_109 V34 V109 -2.7378440240825716e-20

R34_110 V34 V110 -8745185.436357822
L34_110 V34 V110 2.1677293952632703e-11
C34_110 V34 V110 3.0509125830930414e-20

R34_111 V34 V111 16685.645639573624
L34_111 V34 V111 1.2534330340750841e-10
C34_111 V34 V111 1.6478824982531474e-20

R34_112 V34 V112 19632.135035253883
L34_112 V34 V112 3.8214358890237274e-11
C34_112 V34 V112 8.084651071531757e-21

R34_113 V34 V113 16177.11360506191
L34_113 V34 V113 4.5905043660920523e-10
C34_113 V34 V113 2.3955535107765847e-21

R34_114 V34 V114 -40526.09292044511
L34_114 V34 V114 -5.278153831085497e-11
C34_114 V34 V114 -8.93495779534791e-21

R34_115 V34 V115 -18015.850817517927
L34_115 V34 V115 1.6875588842185177e-10
C34_115 V34 V115 -9.400465925120473e-21

R34_116 V34 V116 -372787.15332426975
L34_116 V34 V116 7.212667010758372e-11
C34_116 V34 V116 1.8757253954787702e-20

R34_117 V34 V117 -17239.54956836932
L34_117 V34 V117 2.591420686445979e-10
C34_117 V34 V117 2.5974849617556045e-21

R34_118 V34 V118 31856.287587463255
L34_118 V34 V118 1.0614329049056488e-10
C34_118 V34 V118 3.5644568032165086e-21

R34_119 V34 V119 9911.128899327874
L34_119 V34 V119 5.575243676499338e-11
C34_119 V34 V119 1.6476300825748246e-20

R34_120 V34 V120 -8855.457312503097
L34_120 V34 V120 -1.4627466104023458e-10
C34_120 V34 V120 4.589339706632363e-22

R34_121 V34 V121 9047.96992147607
L34_121 V34 V121 -2.3215781205698435e-10
C34_121 V34 V121 -1.5329529408999624e-20

R34_122 V34 V122 8367.823737569555
L34_122 V34 V122 1.4607094045260957e-10
C34_122 V34 V122 -4.287757291188664e-21

R34_123 V34 V123 -45280.80428443227
L34_123 V34 V123 -9.620935425854318e-11
C34_123 V34 V123 1.079146645008532e-21

R34_124 V34 V124 -56186.94969517174
L34_124 V34 V124 -2.1056840431854915e-10
C34_124 V34 V124 4.11826578138817e-21

R34_125 V34 V125 -5660.07838621441
L34_125 V34 V125 -1.6309015011975647e-10
C34_125 V34 V125 2.821634144875813e-21

R34_126 V34 V126 -17044.84820573858
L34_126 V34 V126 -2.7546110351030547e-11
C34_126 V34 V126 -1.4195714144236222e-20

R34_127 V34 V127 -33901.740163669085
L34_127 V34 V127 5.922765598098653e-11
C34_127 V34 V127 6.491253209434017e-21

R34_128 V34 V128 -87700.42257976283
L34_128 V34 V128 8.991549408511033e-11
C34_128 V34 V128 1.065022807235741e-20

R34_129 V34 V129 -15464.96071274692
L34_129 V34 V129 1.1849982367178433e-10
C34_129 V34 V129 1.3748423785881717e-20

R34_130 V34 V130 118862.06980083199
L34_130 V34 V130 6.4822558866675e-11
C34_130 V34 V130 6.951167625876942e-23

R34_131 V34 V131 -58571.98775948724
L34_131 V34 V131 -8.71984663269886e-11
C34_131 V34 V131 -1.8390919976766673e-20

R34_132 V34 V132 223875.6358130691
L34_132 V34 V132 8.23452199628855e-11
C34_132 V34 V132 1.4395249778961837e-20

R34_133 V34 V133 -369123.7091256891
L34_133 V34 V133 8.824886833047145e-11
C34_133 V34 V133 7.179309092312631e-21

R34_134 V34 V134 20825.224333414695
L34_134 V34 V134 7.243850433329582e-11
C34_134 V34 V134 6.831476659949532e-21

R34_135 V34 V135 64793.44633286939
L34_135 V34 V135 -1.0924189944383282e-10
C34_135 V34 V135 -1.2634997919422779e-20

R34_136 V34 V136 -76506.2170545493
L34_136 V34 V136 -4.4241630426837046e-11
C34_136 V34 V136 -1.6654930182549392e-20

R34_137 V34 V137 -6900.9878598791165
L34_137 V34 V137 -2.611652217236833e-11
C34_137 V34 V137 -1.9551246540713338e-20

R34_138 V34 V138 -27805.527990358456
L34_138 V34 V138 5.183775029782012e-11
C34_138 V34 V138 2.2796335182564784e-20

R34_139 V34 V139 -14056.42404552167
L34_139 V34 V139 8.013570620002989e-10
C34_139 V34 V139 -1.9705505269019312e-21

R34_140 V34 V140 20057.839830742392
L34_140 V34 V140 -4.0542600022564044e-11
C34_140 V34 V140 -1.1917391985960138e-20

R34_141 V34 V141 -15403.88920189703
L34_141 V34 V141 -1.9752913994914978e-10
C34_141 V34 V141 2.8060436533386207e-21

R34_142 V34 V142 10850.217761911426
L34_142 V34 V142 7.599710404904309e-11
C34_142 V34 V142 5.0212858244856e-21

R34_143 V34 V143 33066.71286459452
L34_143 V34 V143 6.277747722180211e-11
C34_143 V34 V143 1.0457499392613082e-20

R34_144 V34 V144 14096.001622372076
L34_144 V34 V144 2.816142389364858e-11
C34_144 V34 V144 1.558098885663229e-20

R35_35 V35 0 120.06805879681744
L35_35 V35 0 9.787113760556132e-14
C35_35 V35 0 1.1560447358536636e-18

R35_36 V35 V36 6561.364417064848
L35_36 V35 V36 6.5035845477688635e-12
C35_36 V35 V36 8.730353044273261e-21

R35_37 V35 V37 3632.213457480202
L35_37 V35 V37 1.1968192926816483e-12
C35_37 V35 V37 1.0177221417983623e-19

R35_38 V35 V38 -10461.589099460705
L35_38 V35 V38 -5.0835755052519945e-12
C35_38 V35 V38 -2.179394285796665e-20

R35_39 V35 V39 3904.146336600454
L35_39 V35 V39 9.9663496807123e-13
C35_39 V35 V39 2.0388747694457912e-19

R35_40 V35 V40 -10909.938901335587
L35_40 V35 V40 -5.366874333296034e-12
C35_40 V35 V40 1.7172392247481568e-20

R35_41 V35 V41 -1077.551694647915
L35_41 V35 V41 -5.506577652429838e-13
C35_41 V35 V41 -2.307077902604583e-19

R35_42 V35 V42 -2225.14895555297
L35_42 V35 V42 -7.249842205306734e-13
C35_42 V35 V42 -2.2347147064093673e-19

R35_43 V35 V43 -2713.12503177362
L35_43 V35 V43 -8.985665463925868e-13
C35_43 V35 V43 -2.1823829284084187e-19

R35_44 V35 V44 4130.4278684004885
L35_44 V35 V44 1.3621711395383129e-12
C35_44 V35 V44 6.066281931603479e-20

R35_45 V35 V45 -8836.155778297925
L35_45 V35 V45 4.949025528095046e-13
C35_45 V35 V45 3.739652586179549e-19

R35_46 V35 V46 -1244.0417430782031
L35_46 V35 V46 -9.898625445308212e-13
C35_46 V35 V46 -1.551191532057725e-19

R35_47 V35 V47 -1252.249469260893
L35_47 V35 V47 -1.325479755666562e-12
C35_47 V35 V47 -2.344011604218845e-20

R35_48 V35 V48 2583.3278959867803
L35_48 V35 V48 3.799225320109121e-12
C35_48 V35 V48 -1.897285434157529e-20

R35_49 V35 V49 1345.0066004996909
L35_49 V35 V49 -1.779452712617782e-11
C35_49 V35 V49 -1.589049573260461e-19

R35_50 V35 V50 -1395.4727886925004
L35_50 V35 V50 -1.5818698645051954e-12
C35_50 V35 V50 5.606725963328584e-20

R35_51 V35 V51 4121.885379049718
L35_51 V35 V51 2.2045098412429197e-12
C35_51 V35 V51 6.998167779380949e-20

R35_52 V35 V52 34383.236171957135
L35_52 V35 V52 -1.1346599747349071e-12
C35_52 V35 V52 -1.4408678331238583e-19

R35_53 V35 V53 -26051.570916535376
L35_53 V35 V53 -1.8703469938625088e-12
C35_53 V35 V53 -4.8636343040802684e-20

R35_54 V35 V54 -3058.3794497638078
L35_54 V35 V54 -3.3975687304377736e-12
C35_54 V35 V54 -3.643769976148294e-21

R35_55 V35 V55 -8547.600374361336
L35_55 V35 V55 -1.707666388466707e-12
C35_55 V35 V55 -1.0241600836289809e-19

R35_56 V35 V56 -3355.9142112247864
L35_56 V35 V56 -2.3901598200220896e-12
C35_56 V35 V56 -4.2394864359290987e-20

R35_57 V35 V57 -299.09329736325594
L35_57 V35 V57 -5.154377675536621e-13
C35_57 V35 V57 4.8959644525576594e-20

R35_58 V35 V58 -1911.5234255607654
L35_58 V35 V58 -3.1054715666873355e-12
C35_58 V35 V58 2.901742847605131e-20

R35_59 V35 V59 -894.739222381029
L35_59 V35 V59 -9.508205069190702e-13
C35_59 V35 V59 2.405534871201015e-20

R35_60 V35 V60 -3220.393891635347
L35_60 V35 V60 -4.2333701881669405e-12
C35_60 V35 V60 1.2572134715546523e-20

R35_61 V35 V61 959.7002368043206
L35_61 V35 V61 5.5863131618285435e-12
C35_61 V35 V61 -1.13762192498964e-19

R35_62 V35 V62 1653.9389109808762
L35_62 V35 V62 -5.5121412592725564e-12
C35_62 V35 V62 -1.2313692671988427e-19

R35_63 V35 V63 7588.4228317632715
L35_63 V35 V63 -3.1973957923856775e-11
C35_63 V35 V63 -1.3322032462249704e-20

R35_64 V35 V64 -8884.288788492586
L35_64 V35 V64 -7.091541067222446e-12
C35_64 V35 V64 7.32384867028293e-22

R35_65 V35 V65 -827.0111591942493
L35_65 V35 V65 -8.848867284453083e-13
C35_65 V35 V65 -8.294594647813029e-20

R35_66 V35 V66 -1371.7202856410474
L35_66 V35 V66 -1.1743556405541964e-12
C35_66 V35 V66 -3.095136863526986e-20

R35_67 V35 V67 -2436.689685042113
L35_67 V35 V67 -2.488500715022404e-12
C35_67 V35 V67 -9.443263433757167e-21

R35_68 V35 V68 15669.163952669209
L35_68 V35 V68 3.4962447184875635e-11
C35_68 V35 V68 -1.5907446772257706e-20

R35_69 V35 V69 2884.734047205127
L35_69 V35 V69 1.629238797161429e-12
C35_69 V35 V69 5.098153218267986e-20

R35_70 V35 V70 19492.20442818118
L35_70 V35 V70 5.604806966146162e-11
C35_70 V35 V70 4.99098507072936e-20

R35_71 V35 V71 8560.049635319723
L35_71 V35 V71 8.54161161600572e-12
C35_71 V35 V71 1.7757522826768805e-20

R35_72 V35 V72 19254.993233497295
L35_72 V35 V72 3.5632570841955127e-12
C35_72 V35 V72 5.371371248365306e-20

R35_73 V35 V73 -20638.09831428076
L35_73 V35 V73 -2.564848998019252e-11
C35_73 V35 V73 4.073124396585216e-21

R35_74 V35 V74 4957.03530112305
L35_74 V35 V74 4.075286149109319e-12
C35_74 V35 V74 -5.715658610328177e-21

R35_75 V35 V75 -10016.675539646647
L35_75 V35 V75 -3.918096695040837e-12
C35_75 V35 V75 -7.445479678467702e-20

R35_76 V35 V76 -8846.75487966453
L35_76 V35 V76 -4.179083292600481e-12
C35_76 V35 V76 -3.466898038183263e-20

R35_77 V35 V77 -27989.095593673155
L35_77 V35 V77 -1.0797456450169916e-11
C35_77 V35 V77 -2.2097003161510127e-20

R35_78 V35 V78 33443.344989785845
L35_78 V35 V78 -7.96293711877759e-11
C35_78 V35 V78 5.984270200388548e-20

R35_79 V35 V79 45849.548025861346
L35_79 V35 V79 3.986250931425691e-11
C35_79 V35 V79 -1.4258195334078883e-20

R35_80 V35 V80 23138.862608266303
L35_80 V35 V80 8.323163929908729e-12
C35_80 V35 V80 9.061115856294184e-22

R35_81 V35 V81 -251950.87568790157
L35_81 V35 V81 -9.472052634556525e-12
C35_81 V35 V81 5.762286600647661e-21

R35_82 V35 V82 714811.1257568762
L35_82 V35 V82 -2.504812727039338e-12
C35_82 V35 V82 -1.903669080747309e-19

R35_83 V35 V83 -29378.189886834283
L35_83 V35 V83 -4.98133105054157e-12
C35_83 V35 V83 -1.2202042531311212e-19

R35_84 V35 V84 -10365.065910331725
L35_84 V35 V84 4.210431127230943e-11
C35_84 V35 V84 1.6687460452105446e-20

R35_85 V35 V85 290401.3326346767
L35_85 V35 V85 9.98482624030591e-12
C35_85 V35 V85 5.85748421078929e-20

R35_86 V35 V86 31353.36760663355
L35_86 V35 V86 5.738205761137012e-12
C35_86 V35 V86 8.632933744662109e-20

R35_87 V35 V87 18666.930850675217
L35_87 V35 V87 7.1148745705480386e-12
C35_87 V35 V87 7.759181220466085e-20

R35_88 V35 V88 23674.83590350843
L35_88 V35 V88 6.847004554237023e-11
C35_88 V35 V88 1.5746194258614475e-20

R35_89 V35 V89 -21405.577784907604
L35_89 V35 V89 -8.045495869018162e-12
C35_89 V35 V89 -9.590681810522184e-20

R35_90 V35 V90 25752.141758279886
L35_90 V35 V90 -5.967407334882334e-11
C35_90 V35 V90 -4.321075944624007e-21

R35_91 V35 V91 -16148.978066150845
L35_91 V35 V91 -2.163688144280504e-12
C35_91 V35 V91 -2.0784151129434207e-19

R35_92 V35 V92 -74127.30020276183
L35_92 V35 V92 -3.813237089322192e-11
C35_92 V35 V92 -6.134228887653621e-20

R35_93 V35 V93 5443.8047467011575
L35_93 V35 V93 2.4079904663762706e-11
C35_93 V35 V93 -3.2572106321852315e-21

R35_94 V35 V94 12217.480362546272
L35_94 V35 V94 1.1255291598634765e-11
C35_94 V35 V94 7.208983394146778e-20

R35_95 V35 V95 -70106.38959853986
L35_95 V35 V95 -4.926081449676795e-12
C35_95 V35 V95 -1.0117787975528619e-19

R35_96 V35 V96 -14197.305103743758
L35_96 V35 V96 7.0960374007317635e-12
C35_96 V35 V96 -6.196006568767703e-21

R35_97 V35 V97 16586.99437834284
L35_97 V35 V97 1.441265149515406e-11
C35_97 V35 V97 4.556519335339563e-20

R35_98 V35 V98 21447.04177643082
L35_98 V35 V98 -8.887103625632685e-12
C35_98 V35 V98 -7.159208800759658e-20

R35_99 V35 V99 25085.7905304341
L35_99 V35 V99 -1.29933966464615e-10
C35_99 V35 V99 3.326286015103723e-21

R35_100 V35 V100 -34875.74900712844
L35_100 V35 V100 -5.0179623907812185e-11
C35_100 V35 V100 2.845601916015723e-21

R35_101 V35 V101 43829.265397121075
L35_101 V35 V101 -7.010870236352727e-12
C35_101 V35 V101 -1.064083047341537e-19

R35_102 V35 V102 11172.069590949217
L35_102 V35 V102 -6.489717406332048e-12
C35_102 V35 V102 -6.610692222693299e-20

R35_103 V35 V103 58079.38563725639
L35_103 V35 V103 -2.130223038769203e-11
C35_103 V35 V103 -3.3665586547119464e-20

R35_104 V35 V104 208772.62284403306
L35_104 V35 V104 5.601395533678063e-12
C35_104 V35 V104 2.5340988881607986e-20

R35_105 V35 V105 -25042.136157432513
L35_105 V35 V105 5.577321909521281e-12
C35_105 V35 V105 9.353738985782685e-20

R35_106 V35 V106 -7661.921573838693
L35_106 V35 V106 -2.858134852403279e-12
C35_106 V35 V106 -1.8034913612624808e-19

R35_107 V35 V107 -159766.35379495958
L35_107 V35 V107 -1.844146375100016e-11
C35_107 V35 V107 -1.3311124380636915e-20

R35_108 V35 V108 -63747.03206296888
L35_108 V35 V108 9.947288698196901e-11
C35_108 V35 V108 3.2034509293371003e-20

R35_109 V35 V109 89018.85535385687
L35_109 V35 V109 6.909875101429727e-12
C35_109 V35 V109 3.4556166491853795e-20

R35_110 V35 V110 8986.273766800556
L35_110 V35 V110 3.121006080274714e-12
C35_110 V35 V110 1.7971498334694666e-19

R35_111 V35 V111 -13889.010068527941
L35_111 V35 V111 2.445498824782956e-11
C35_111 V35 V111 2.1173641125380674e-20

R35_112 V35 V112 -30640.26953291691
L35_112 V35 V112 -8.010096300892971e-12
C35_112 V35 V112 -5.795658321553277e-20

R35_113 V35 V113 -13891.559940964207
L35_113 V35 V113 -6.683523463376195e-12
C35_113 V35 V113 -5.589637247513755e-20

R35_114 V35 V114 -29329.09981053838
L35_114 V35 V114 -7.109854153077093e-12
C35_114 V35 V114 -9.41358449458186e-20

R35_115 V35 V115 13516.443177254598
L35_115 V35 V115 -2.966177747730628e-11
C35_115 V35 V115 -2.902389537944321e-21

R35_116 V35 V116 -64304.84294198016
L35_116 V35 V116 3.908133343512311e-11
C35_116 V35 V116 2.4383359782053824e-20

R35_117 V35 V117 11643.673633093966
L35_117 V35 V117 7.735450551021175e-12
C35_117 V35 V117 5.705323049529886e-20

R35_118 V35 V118 -709082.3604433228
L35_118 V35 V118 4.753422954815298e-12
C35_118 V35 V118 9.654865034372255e-20

R35_119 V35 V119 -13737.602243593843
L35_119 V35 V119 6.5514482557536035e-12
C35_119 V35 V119 9.891269661000947e-20

R35_120 V35 V120 4820.699664034406
L35_120 V35 V120 -9.00375978113495e-11
C35_120 V35 V120 8.840294357986636e-21

R35_121 V35 V121 -9674.771465811906
L35_121 V35 V121 -1.056654323879335e-11
C35_121 V35 V121 -2.3167545473489957e-20

R35_122 V35 V122 -39496.641246905034
L35_122 V35 V122 -1.9102937592125628e-11
C35_122 V35 V122 -9.217980662568288e-21

R35_123 V35 V123 29212.062717932942
L35_123 V35 V123 1.2353628167884589e-11
C35_123 V35 V123 3.234702491665501e-20

R35_124 V35 V124 39136.78127987955
L35_124 V35 V124 9.663204256839058e-11
C35_124 V35 V124 1.1392348767736933e-20

R35_125 V35 V125 4897.684170851137
L35_125 V35 V125 2.0032196245837686e-11
C35_125 V35 V125 8.060895799702879e-21

R35_126 V35 V126 -11993.22563854212
L35_126 V35 V126 1.5613450016134478e-10
C35_126 V35 V126 -2.3697535570645185e-20

R35_127 V35 V127 6585.392035687092
L35_127 V35 V127 -2.521089426594821e-11
C35_127 V35 V127 3.509618264063735e-22

R35_128 V35 V128 26718.97266809866
L35_128 V35 V128 3.541499174572001e-11
C35_128 V35 V128 2.0385451859061824e-20

R35_129 V35 V129 9362.927303828861
L35_129 V35 V129 2.180016607680745e-11
C35_129 V35 V129 3.165404583897659e-20

R35_130 V35 V130 50478.4155767438
L35_130 V35 V130 2.5612866920636404e-10
C35_130 V35 V130 2.586722550916276e-20

R35_131 V35 V131 163302.13368448906
L35_131 V35 V131 -3.027481996686656e-11
C35_131 V35 V131 -7.369024267148173e-21

R35_132 V35 V132 -31292.784867425056
L35_132 V35 V132 -2.878646072684231e-11
C35_132 V35 V132 -1.207286534277485e-21

R35_133 V35 V133 -28558.41090541144
L35_133 V35 V133 -7.1903892674897364e-12
C35_133 V35 V133 -7.1931043704385e-20

R35_134 V35 V134 -18045.648220173876
L35_134 V35 V134 1.2672850325339053e-10
C35_134 V35 V134 5.616810219294602e-21

R35_135 V35 V135 19906.14269969323
L35_135 V35 V135 -3.6475111474333844e-11
C35_135 V35 V135 -1.1354799255619889e-20

R35_136 V35 V136 53232.68407915445
L35_136 V35 V136 -8.759388809125083e-11
C35_136 V35 V136 -1.0076313326446524e-20

R35_137 V35 V137 5394.288981993675
L35_137 V35 V137 1.580363065616466e-11
C35_137 V35 V137 2.0714244561071957e-20

R35_138 V35 V138 -17387.172487440053
L35_138 V35 V138 1.3374193182253023e-10
C35_138 V35 V138 6.450262239752688e-21

R35_139 V35 V139 4888.798273070887
L35_139 V35 V139 -2.5291358274903883e-11
C35_139 V35 V139 -1.72512174187889e-22

R35_140 V35 V140 -10140.476584444616
L35_140 V35 V140 3.714061996297311e-11
C35_140 V35 V140 5.487193026096635e-21

R35_141 V35 V141 20912.00703646955
L35_141 V35 V141 4.410300092641006e-11
C35_141 V35 V141 2.248647161881543e-21

R35_142 V35 V142 -8063.582372028328
L35_142 V35 V142 2.0243107122694983e-11
C35_142 V35 V142 2.276702978892006e-20

R35_143 V35 V143 -14326.055048526714
L35_143 V35 V143 -4.387399633667388e-11
C35_143 V35 V143 -3.9250910087163194e-21

R35_144 V35 V144 -13851.439267376167
L35_144 V35 V144 -4.0958349905275086e-11
C35_144 V35 V144 -2.1609339555210676e-20

R36_36 V36 0 -3331.393208396566
L36_36 V36 0 -2.3946772199329958e-12
C36_36 V36 0 -4.870141201547591e-20

R36_37 V36 V37 -18259.90401838387
L36_37 V36 V37 -5.788917190617562e-12
C36_37 V36 V37 1.8074705068748452e-21

R36_38 V36 V38 30581.758547778016
L36_38 V36 V38 -4.608784746344943e-11
C36_38 V36 V38 -5.244116993647597e-21

R36_39 V36 V39 -13188.65539565363
L36_39 V36 V39 -4.622802885098657e-12
C36_39 V36 V39 -1.2259472566424827e-20

R36_40 V36 V40 18337.568200801506
L36_40 V36 V40 2.120259899101845e-12
C36_40 V36 V40 7.316213646634365e-20

R36_41 V36 V41 4334.434482863044
L36_41 V36 V41 2.4320480214880064e-12
C36_41 V36 V41 -1.71217349180184e-20

R36_42 V36 V42 4635.917496437755
L36_42 V36 V42 2.0379211981672955e-12
C36_42 V36 V42 8.00444710744663e-21

R36_43 V36 V43 14150.82853249078
L36_43 V36 V43 4.4752410988248426e-12
C36_43 V36 V43 2.2972435104903077e-21

R36_44 V36 V44 -2294.684588026703
L36_44 V36 V44 -1.0443160613527781e-12
C36_44 V36 V44 -1.1813070853121324e-19

R36_45 V36 V45 4189.393138192901
L36_45 V36 V45 -3.062510007872727e-11
C36_45 V36 V45 5.76228784699209e-20

R36_46 V36 V46 3668.890707513822
L36_46 V36 V46 -9.583639714415386e-12
C36_46 V36 V46 -1.7834874472236432e-20

R36_47 V36 V47 333130.0810326606
L36_47 V36 V47 -3.514790558770543e-10
C36_47 V36 V47 -2.193296817789406e-21

R36_48 V36 V48 -2078.5286497611783
L36_48 V36 V48 -6.84056823430094e-12
C36_48 V36 V48 4.558282127849221e-20

R36_49 V36 V49 -4609.504499622074
L36_49 V36 V49 8.226420991133332e-11
C36_49 V36 V49 -7.427084535920738e-21

R36_50 V36 V50 4674.740186312312
L36_50 V36 V50 7.231588214279072e-12
C36_50 V36 V50 7.347337056571234e-23

R36_51 V36 V51 -6315.777338678028
L36_51 V36 V51 -6.421492766468737e-12
C36_51 V36 V51 1.6374077682419626e-21

R36_52 V36 V52 9550.086425803769
L36_52 V36 V52 5.292497686280279e-12
C36_52 V36 V52 -1.760232055405227e-20

R36_53 V36 V53 -7711.585158884601
L36_53 V36 V53 4.284976230255878e-12
C36_53 V36 V53 2.73519659278717e-20

R36_54 V36 V54 17966.765698938965
L36_54 V36 V54 1.0261835819958634e-11
C36_54 V36 V54 8.93354004389352e-21

R36_55 V36 V55 9678.817657676755
L36_55 V36 V55 8.691969456879909e-12
C36_55 V36 V55 -6.136534455857658e-21

R36_56 V36 V56 3256.7017203800865
L36_56 V36 V56 -6.99509209278622e-12
C36_56 V36 V56 -5.98706038675423e-20

R36_57 V36 V57 936.6626449662278
L36_57 V36 V57 2.2075184599452456e-12
C36_57 V36 V57 -1.0764192071885346e-20

R36_58 V36 V58 2042.8154220580063
L36_58 V36 V58 4.056834032786701e-12
C36_58 V36 V58 5.241323891581702e-21

R36_59 V36 V59 4219.796811701852
L36_59 V36 V59 8.333826962691884e-12
C36_59 V36 V59 7.003945992081673e-21

R36_60 V36 V60 -808.8758395958588
L36_60 V36 V60 -1.3726849655431369e-12
C36_60 V36 V60 -2.5745948368386103e-21

R36_61 V36 V61 -3546.999946332965
L36_61 V36 V61 3.0711332389150366e-11
C36_61 V36 V61 1.8449541916037293e-20

R36_62 V36 V62 -2001.5465099322607
L36_62 V36 V62 -8.044411185634193e-12
C36_62 V36 V62 4.156825567852386e-21

R36_63 V36 V63 -83214.28734672976
L36_63 V36 V63 -2.1262044225810258e-11
C36_63 V36 V63 -1.3640929774696632e-20

R36_64 V36 V64 8335.65853548507
L36_64 V36 V64 -1.5116268260863174e-11
C36_64 V36 V64 1.6005443505597844e-21

R36_65 V36 V65 3031.30897644775
L36_65 V36 V65 3.4396768137781014e-12
C36_65 V36 V65 5.8959248444009284e-21

R36_66 V36 V66 2888.9645207670887
L36_66 V36 V66 3.722655595281345e-12
C36_66 V36 V66 1.1344878651023742e-20

R36_67 V36 V67 42329.529447351626
L36_67 V36 V67 6.989805516220559e-11
C36_67 V36 V67 -6.875032336559804e-21

R36_68 V36 V68 -2159.548551695769
L36_68 V36 V68 -2.8690661346792174e-12
C36_68 V36 V68 -4.336375515374468e-21

R36_69 V36 V69 9823.112934390952
L36_69 V36 V69 1.296779150774412e-11
C36_69 V36 V69 1.8037121934283156e-20

R36_70 V36 V70 -8269.436688147112
L36_70 V36 V70 -1.1036826140514288e-11
C36_70 V36 V70 8.139879280370716e-21

R36_71 V36 V71 48794.885928132804
L36_71 V36 V71 -3.079870728364419e-11
C36_71 V36 V71 -5.289501081992549e-22

R36_72 V36 V72 -87813.81318398628
L36_72 V36 V72 -1.1496866392747194e-11
C36_72 V36 V72 -1.5083968614203818e-20

R36_73 V36 V73 -7603.834105149405
L36_73 V36 V73 -1.604218290290143e-11
C36_73 V36 V73 2.7564593884619603e-20

R36_74 V36 V74 -18950.07675773508
L36_74 V36 V74 -1.5368490935090364e-11
C36_74 V36 V74 -1.3223580870263642e-21

R36_75 V36 V75 12311.497897017838
L36_75 V36 V75 1.3761809323874026e-11
C36_75 V36 V75 -1.804205578475385e-20

R36_76 V36 V76 12596.50095747908
L36_76 V36 V76 1.4016251539202168e-11
C36_76 V36 V76 2.5010866918133533e-20

R36_77 V36 V77 27183.737162244168
L36_77 V36 V77 1.6098565050481156e-11
C36_77 V36 V77 -3.469265002167724e-20

R36_78 V36 V78 -695652.5014309759
L36_78 V36 V78 6.33388218157231e-11
C36_78 V36 V78 1.4644372920619584e-20

R36_79 V36 V79 -163252.13791023017
L36_79 V36 V79 -5.7200474380290324e-11
C36_79 V36 V79 1.7560331709864995e-20

R36_80 V36 V80 -31894.269872096047
L36_80 V36 V80 -1.8252165102249364e-11
C36_80 V36 V80 -6.655316871747125e-20

R36_81 V36 V81 39881.013100374614
L36_81 V36 V81 1.6536458108351166e-11
C36_81 V36 V81 1.2993978173549625e-19

R36_82 V36 V82 -37788.75617775046
L36_82 V36 V82 1.6381493265200313e-11
C36_82 V36 V82 -8.53078667360191e-21

R36_83 V36 V83 -121237.40088734945
L36_83 V36 V83 -5.41598669966653e-11
C36_83 V36 V83 -6.430924459917407e-20

R36_84 V36 V84 28514.35247750972
L36_84 V36 V84 -2.1850872169301004e-11
C36_84 V36 V84 -1.880295293804926e-20

R36_85 V36 V85 -64163.55155000339
L36_85 V36 V85 -3.632789542179993e-11
C36_85 V36 V85 2.1256168227120188e-20

R36_86 V36 V86 -17916.226528778272
L36_86 V36 V86 -4.3144608214337234e-11
C36_86 V36 V86 -5.696412409771288e-21

R36_87 V36 V87 46802.88688363948
L36_87 V36 V87 -4.3518487635577065e-11
C36_87 V36 V87 2.1021236145213877e-20

R36_88 V36 V88 113899.0661408571
L36_88 V36 V88 5.86598129306981e-11
C36_88 V36 V88 3.192308770888354e-20

R36_89 V36 V89 81935.64724228841
L36_89 V36 V89 4.5062921899273814e-11
C36_89 V36 V89 -9.492012248887202e-21

R36_90 V36 V90 -96883.7761725964
L36_90 V36 V90 2.9842919068357997e-10
C36_90 V36 V90 -9.032315617998347e-21

R36_91 V36 V91 165899.3106374229
L36_91 V36 V91 1.8892354697089673e-11
C36_91 V36 V91 1.7473703501645047e-20

R36_92 V36 V92 -21427.30543486567
L36_92 V36 V92 -1.97337847880496e-11
C36_92 V36 V92 -1.1198036789919236e-19

R36_93 V36 V93 -14165.893698302803
L36_93 V36 V93 -4.70895768777352e-10
C36_93 V36 V93 1.8561500377159962e-20

R36_94 V36 V94 -56348.63751089534
L36_94 V36 V94 6.493476895688389e-11
C36_94 V36 V94 5.025909071648718e-20

R36_95 V36 V95 264176.03326874046
L36_95 V36 V95 4.610099520182721e-11
C36_95 V36 V95 -1.411948195571936e-21

R36_96 V36 V96 -85626.3888162328
L36_96 V36 V96 -1.4359448485331003e-11
C36_96 V36 V96 -1.282311297639598e-19

R36_97 V36 V97 -135766.38408228647
L36_97 V36 V97 6.807387231619419e-11
C36_97 V36 V97 3.083988103357905e-20

R36_98 V36 V98 -56747.38131242537
L36_98 V36 V98 1.0679909764751944e-10
C36_98 V36 V98 -3.7306186359916855e-20

R36_99 V36 V99 -87603.88538507947
L36_99 V36 V99 1.549085899830651e-10
C36_99 V36 V99 1.8625526054932577e-20

R36_100 V36 V100 22423.92730047387
L36_100 V36 V100 8.32181373880827e-11
C36_100 V36 V100 5.0956330805334216e-20

R36_101 V36 V101 -25789.553603374057
L36_101 V36 V101 5.881615218226229e-11
C36_101 V36 V101 -3.023634334566566e-20

R36_102 V36 V102 -57223.60447046775
L36_102 V36 V102 2.7695171663496675e-11
C36_102 V36 V102 -1.0045566598760637e-20

R36_103 V36 V103 -72753.01252866194
L36_103 V36 V103 -4.1093929744173294e-10
C36_103 V36 V103 1.838501364527905e-20

R36_104 V36 V104 -23274.57205015646
L36_104 V36 V104 -1.0983009953889833e-11
C36_104 V36 V104 -1.0980472525892984e-19

R36_105 V36 V105 14514.194403764353
L36_105 V36 V105 7.213684232727108e-11
C36_105 V36 V105 6.835110866421561e-20

R36_106 V36 V106 -4173174.432272364
L36_106 V36 V106 6.038350509162893e-11
C36_106 V36 V106 -5.732146121981014e-20

R36_107 V36 V107 -219787.86600033642
L36_107 V36 V107 5.796128012768295e-11
C36_107 V36 V107 -2.0812368890553836e-20

R36_108 V36 V108 14442.687669518924
L36_108 V36 V108 -1.0526445233955291e-09
C36_108 V36 V108 5.977395468462479e-20

R36_109 V36 V109 -20427.28773837399
L36_109 V36 V109 -1.2923270631842723e-11
C36_109 V36 V109 -9.858917937918791e-20

R36_110 V36 V110 78358.86081313231
L36_110 V36 V110 -4.4763740092813306e-11
C36_110 V36 V110 4.277969199359637e-20

R36_111 V36 V111 32430.40517737213
L36_111 V36 V111 -1.1492468112543766e-09
C36_111 V36 V111 3.4995753007881696e-20

R36_112 V36 V112 39082.830841946445
L36_112 V36 V112 2.0342861866928668e-11
C36_112 V36 V112 -2.346372022309029e-20

R36_113 V36 V113 14535.21417306269
L36_113 V36 V113 3.256611833803346e-11
C36_113 V36 V113 2.8770867447319234e-20

R36_114 V36 V114 488305.41155266727
L36_114 V36 V114 3.6099510044707643e-11
C36_114 V36 V114 -2.2961852433041696e-20

R36_115 V36 V115 -72704.87385977976
L36_115 V36 V115 1.0999258496656652e-10
C36_115 V36 V115 -1.4993415893147615e-20

R36_116 V36 V116 48775.67361468114
L36_116 V36 V116 -7.282400848849632e-10
C36_116 V36 V116 4.1090401568499113e-20

R36_117 V36 V117 -23068.104754919976
L36_117 V36 V117 -8.51746102253269e-11
C36_117 V36 V117 -1.1939367845916637e-20

R36_118 V36 V118 -489549.6170924603
L36_118 V36 V118 -2.757579365023506e-11
C36_118 V36 V118 -9.09464138701308e-21

R36_119 V36 V119 16242.72125701284
L36_119 V36 V119 -1.1971843120616366e-10
C36_119 V36 V119 4.8703704596030385e-20

R36_120 V36 V120 -27623.680193617598
L36_120 V36 V120 1.2324765980133917e-10
C36_120 V36 V120 3.196600647323135e-20

R36_121 V36 V121 17766.753418633707
L36_121 V36 V121 4.374020139838278e-11
C36_121 V36 V121 -3.548617154289135e-21

R36_122 V36 V122 10640.000183803046
L36_122 V36 V122 2.793581175299901e-11
C36_122 V36 V122 -3.6011542422470224e-21

R36_123 V36 V123 716493.2929164806
L36_123 V36 V123 -1.1915496807530192e-10
C36_123 V36 V123 -4.64082362363795e-21

R36_124 V36 V124 47949.71581176025
L36_124 V36 V124 3.3401215197655046e-11
C36_124 V36 V124 4.1881358278611236e-20

R36_125 V36 V125 -11106.612861091311
L36_125 V36 V125 -6.473769861469389e-11
C36_125 V36 V125 4.935321454980324e-21

R36_126 V36 V126 -20969.60439236406
L36_126 V36 V126 -3.8790034135769726e-11
C36_126 V36 V126 1.33994674262219e-22

R36_127 V36 V127 148041.7037718201
L36_127 V36 V127 3.9666392450807665e-11
C36_127 V36 V127 6.468059158366513e-21

R36_128 V36 V128 -139354.80312886392
L36_128 V36 V128 8.976444207935283e-11
C36_128 V36 V128 3.879814419302784e-21

R36_129 V36 V129 -155165.68427445498
L36_129 V36 V129 7.71933772711893e-11
C36_129 V36 V129 8.717286288865016e-21

R36_130 V36 V130 -55599.35796357718
L36_130 V36 V130 7.359422363691017e-11
C36_130 V36 V130 1.4748636657302702e-20

R36_131 V36 V131 -30056.154878700203
L36_131 V36 V131 2.466077341512367e-10
C36_131 V36 V131 -4.710151056207934e-21

R36_132 V36 V132 759196.3137613162
L36_132 V36 V132 4.7710305449757716e-11
C36_132 V36 V132 2.856526429326821e-20

R36_133 V36 V133 -112723.13755787486
L36_133 V36 V133 -1.6689316551829022e-10
C36_133 V36 V133 -2.0251766563470432e-20

R36_134 V36 V134 115130.48976867854
L36_134 V36 V134 4.64795369772767e-10
C36_134 V36 V134 3.2850030275202186e-21

R36_135 V36 V135 54839.38045629415
L36_135 V36 V135 6.60901265180941e-11
C36_135 V36 V135 7.506959421316966e-21

R36_136 V36 V136 -118882.31799937779
L36_136 V36 V136 -3.7427561649533476e-11
C36_136 V36 V136 -1.2838315228524124e-20

R36_137 V36 V137 -17130.37621931863
L36_137 V36 V137 -6.033093765563119e-11
C36_137 V36 V137 1.4998910769699193e-20

R36_138 V36 V138 -19374.47235887821
L36_138 V36 V138 -2.2695903565637793e-11
C36_138 V36 V138 2.355405029437537e-21

R36_139 V36 V139 -149197.73326612488
L36_139 V36 V139 4.330657425849599e-11
C36_139 V36 V139 -8.0199270647771e-21

R36_140 V36 V140 33863.657580706946
L36_140 V36 V140 -2.0536629840193415e-10
C36_140 V36 V140 2.3669337483346622e-21

R36_141 V36 V141 -24134.869091240787
L36_141 V36 V141 -5.396296064008705e-11
C36_141 V36 V141 -1.0720305557983154e-20

R36_142 V36 V142 19170.208530596927
L36_142 V36 V142 -2.0826628700729338e-10
C36_142 V36 V142 1.0920586191429477e-20

R36_143 V36 V143 69590.1764082093
L36_143 V36 V143 -2.965343129818138e-10
C36_143 V36 V143 6.0442967345428115e-21

R36_144 V36 V144 24131.112044474474
L36_144 V36 V144 3.9542777009624673e-11
C36_144 V36 V144 1.2439326120115268e-20

R37_37 V37 0 -349.0490472136228
L37_37 V37 0 -4.4774741571089503e-14
C37_37 V37 0 -5.46974073774562e-18

R37_38 V37 V38 14381.823408533255
L37_38 V37 V38 6.615774295072415e-12
C37_38 V37 V38 -8.492524985342332e-21

R37_39 V37 V39 -3337.1622556426373
L37_39 V37 V39 -6.318680690081844e-13
C37_39 V37 V39 -5.603917693176921e-19

R37_40 V37 V40 22172.940603736555
L37_40 V37 V40 2.1466779717409005e-11
C37_40 V37 V40 -2.380739292984748e-20

R37_41 V37 V41 1023.5697311658813
L37_41 V37 V41 1.8557493516331813e-13
C37_41 V37 V41 2.197738616476753e-18

R37_42 V37 V42 1627.2138179181488
L37_42 V37 V42 2.7007078525048766e-13
C37_42 V37 V42 1.5657731206066262e-18

R37_43 V37 V43 2205.002789105791
L37_43 V37 V43 4.627761543211613e-13
C37_43 V37 V43 8.331590914656555e-19

R37_44 V37 V44 -7823.430316169315
L37_44 V37 V44 -3.5401586131897856e-12
C37_44 V37 V44 -7.605049144679943e-21

R37_45 V37 V45 -1003.4717067562169
L37_45 V37 V45 -3.7420869282714485e-13
C37_45 V37 V45 -1.6785686418916669e-18

R37_46 V37 V46 -5186.883544121982
L37_46 V37 V46 2.765161565531983e-12
C37_46 V37 V46 -6.517896374602867e-19

R37_47 V37 V47 3669.6786823425446
L37_47 V37 V47 1.7768697607017196e-12
C37_47 V37 V47 -2.309931213226353e-19

R37_48 V37 V48 -4495.808397131187
L37_48 V37 V48 -2.7155830404591564e-12
C37_48 V37 V48 -4.4388581219977e-20

R37_49 V37 V49 -4399.614331955292
L37_49 V37 V49 5.191837400758334e-12
C37_49 V37 V49 4.448531777895532e-19

R37_50 V37 V50 1706.1737474759132
L37_50 V37 V50 9.34963628224649e-13
C37_50 V37 V50 2.9072329514397155e-19

R37_51 V37 V51 -6664.4904891608485
L37_51 V37 V51 -1.1025962991961184e-12
C37_51 V37 V51 -2.9311140676406274e-19

R37_52 V37 V52 1942.5270960960963
L37_52 V37 V52 5.983641307588767e-13
C37_52 V37 V52 1.0265106405327717e-18

R37_53 V37 V53 3159.114294498699
L37_53 V37 V53 9.56790665352369e-13
C37_53 V37 V53 5.280431623777851e-19

R37_54 V37 V54 19131.497947344633
L37_54 V37 V54 1.7252584561300495e-12
C37_54 V37 V54 7.620497472205643e-20

R37_55 V37 V55 -12504.82636047174
L37_55 V37 V55 8.694610393588018e-13
C37_55 V37 V55 3.1854766226750876e-19

R37_56 V37 V56 6539.639355129991
L37_56 V37 V56 1.1955431495311546e-12
C37_56 V37 V56 2.564737402443451e-19

R37_57 V37 V57 -5984.579935220864
L37_57 V37 V57 1.985645338948189e-13
C37_57 V37 V57 -1.8976008933883238e-19

R37_58 V37 V58 -2580.669997425738
L37_58 V37 V58 1.1107921784001639e-12
C37_58 V37 V58 -1.1395989587237105e-19

R37_59 V37 V59 1453.314972259544
L37_59 V37 V59 1.6437890172152117e-12
C37_59 V37 V59 -1.307437765694991e-19

R37_60 V37 V60 -10042.627844305754
L37_60 V37 V60 1.3893311575092453e-12
C37_60 V37 V60 -4.808053373555467e-20

R37_61 V37 V61 2995.1035988022236
L37_61 V37 V61 -2.691762750920643e-12
C37_61 V37 V61 6.748793004918333e-19

R37_62 V37 V62 1674.1324606492894
L37_62 V37 V62 -3.9129329337924025e-12
C37_62 V37 V62 5.886755392154589e-19

R37_63 V37 V63 196692.46379742504
L37_63 V37 V63 5.06869928069253e-12
C37_63 V37 V63 1.330295642544826e-19

R37_64 V37 V64 9308.94448483986
L37_64 V37 V64 5.583619922581317e-12
C37_64 V37 V64 7.076289435202696e-20

R37_65 V37 V65 9973.169275035078
L37_65 V37 V65 4.654717523809194e-13
C37_65 V37 V65 2.5310134289053127e-19

R37_66 V37 V66 -6487.263024692882
L37_66 V37 V66 6.030349137783931e-13
C37_66 V37 V66 1.1963164856442034e-19

R37_67 V37 V67 5544.682462510143
L37_67 V37 V67 1.809152856863701e-12
C37_67 V37 V67 1.0030798818212872e-19

R37_68 V37 V68 -10366.148922359847
L37_68 V37 V68 3.884457115553824e-12
C37_68 V37 V68 8.359778083220822e-20

R37_69 V37 V69 -4377.725819564655
L37_69 V37 V69 -1.9761482890890572e-12
C37_69 V37 V69 -4.631813980960696e-20

R37_70 V37 V70 5905.677383822921
L37_70 V37 V70 1.0521761367814382e-11
C37_70 V37 V70 3.7008921015452485e-20

R37_71 V37 V71 -95888.18418356293
L37_71 V37 V71 8.549222544387958e-12
C37_71 V37 V71 2.843322717990365e-20

R37_72 V37 V72 7881.951246413082
L37_72 V37 V72 -3.6550854177593546e-12
C37_72 V37 V72 -1.639091248515716e-20

R37_73 V37 V73 28459.624838918007
L37_73 V37 V73 4.3498514678409535e-12
C37_73 V37 V73 9.374900777295584e-20

R37_74 V37 V74 -9048.242524716869
L37_74 V37 V74 -2.5423085485315923e-12
C37_74 V37 V74 -7.154090368661989e-20

R37_75 V37 V75 -101166.36201920341
L37_75 V37 V75 3.005178890681342e-12
C37_75 V37 V75 1.0214288038764894e-19

R37_76 V37 V76 36242.938708730544
L37_76 V37 V76 2.2779758678557667e-12
C37_76 V37 V76 1.0895556418414194e-19

R37_77 V37 V77 -986790.7770013578
L37_77 V37 V77 5.972750738861899e-12
C37_77 V37 V77 2.2566720057545992e-20

R37_78 V37 V78 72352.35081282162
L37_78 V37 V78 1.04470352723369e-11
C37_78 V37 V78 7.058331593298598e-21

R37_79 V37 V79 67821.65036382739
L37_79 V37 V79 2.7253160382419027e-11
C37_79 V37 V79 2.4366292479283446e-20

R37_80 V37 V80 228169.05535271493
L37_80 V37 V80 -1.54978502397546e-11
C37_80 V37 V80 -8.757177027253379e-21

R37_81 V37 V81 93268.98237256709
L37_81 V37 V81 5.829782168374157e-11
C37_81 V37 V81 1.493925599029277e-20

R37_82 V37 V82 45051.03057746985
L37_82 V37 V82 7.362172034460118e-12
C37_82 V37 V82 1.2745873643725956e-19

R37_83 V37 V83 34884.547956664086
L37_83 V37 V83 5.2803739183865685e-12
C37_83 V37 V83 1.0625167684804435e-19

R37_84 V37 V84 54076.602545535556
L37_84 V37 V84 1.6027143346276113e-11
C37_84 V37 V84 7.216652033834422e-21

R37_85 V37 V85 81023.13212592626
L37_85 V37 V85 2.655773236140646e-11
C37_85 V37 V85 -9.179964208928314e-21

R37_86 V37 V86 -29217.458153304422
L37_86 V37 V86 -1.2344120796629732e-11
C37_86 V37 V86 -7.39919045109643e-20

R37_87 V37 V87 -22768.27073039102
L37_87 V37 V87 -1.063911867060757e-11
C37_87 V37 V87 -5.229390218033096e-20

R37_88 V37 V88 104736.98830110338
L37_88 V37 V88 -2.545453867550922e-11
C37_88 V37 V88 6.81494383155874e-21

R37_89 V37 V89 56741.75260215957
L37_89 V37 V89 8.399308711813267e-12
C37_89 V37 V89 6.164108942914226e-20

R37_90 V37 V90 -108653.5157110656
L37_90 V37 V90 -6.212665467710353e-11
C37_90 V37 V90 -8.211618325153387e-21

R37_91 V37 V91 15750.161669243205
L37_91 V37 V91 3.814813601224676e-12
C37_91 V37 V91 1.71251006702604e-19

R37_92 V37 V92 2614919.318199618
L37_92 V37 V92 1.1340122764282622e-11
C37_92 V37 V92 4.109593760667899e-20

R37_93 V37 V93 27202.758358611736
L37_93 V37 V93 -3.056614081048928e-11
C37_93 V37 V93 -7.607527822516373e-21

R37_94 V37 V94 -713927.9300494984
L37_94 V37 V94 -8.595057201184999e-12
C37_94 V37 V94 -4.591771809382158e-20

R37_95 V37 V95 45197.41580292975
L37_95 V37 V95 1.0390241250031946e-11
C37_95 V37 V95 6.413580922960185e-20

R37_96 V37 V96 129018.63465410365
L37_96 V37 V96 -4.714940890062119e-11
C37_96 V37 V96 -3.0546960342042033e-20

R37_97 V37 V97 976605.3376623632
L37_97 V37 V97 -1.0921180516161613e-10
C37_97 V37 V97 -3.4553697611605803e-20

R37_98 V37 V98 145326.0874779199
L37_98 V37 V98 5.897834316116657e-12
C37_98 V37 V98 5.324515539485508e-20

R37_99 V37 V99 -117681.61749673498
L37_99 V37 V99 5.626760398900678e-11
C37_99 V37 V99 -4.617276156315268e-21

R37_100 V37 V100 195383.89798933777
L37_100 V37 V100 -3.52253686623211e-11
C37_100 V37 V100 1.577053932493239e-21

R37_101 V37 V101 20230.394554469647
L37_101 V37 V101 5.496663645110492e-12
C37_101 V37 V101 8.343814452415242e-20

R37_102 V37 V102 -226472.9345628602
L37_102 V37 V102 1.292323953589069e-11
C37_102 V37 V102 5.588281824140147e-20

R37_103 V37 V103 47364.23854295944
L37_103 V37 V103 9.504085009953912e-12
C37_103 V37 V103 7.28941635630182e-20

R37_104 V37 V104 -37612.0882737754
L37_104 V37 V104 -1.5967632998771725e-11
C37_104 V37 V104 -5.966123307709148e-20

R37_105 V37 V105 -36948.48634955079
L37_105 V37 V105 -8.280874180222764e-12
C37_105 V37 V105 -7.746767737238797e-20

R37_106 V37 V106 19388.08903973755
L37_106 V37 V106 6.7997633290529766e-12
C37_106 V37 V106 1.1854159943388435e-19

R37_107 V37 V107 251146.68202604502
L37_107 V37 V107 8.762253987681123e-11
C37_107 V37 V107 1.601287151025912e-20

R37_108 V37 V108 -24695.974404512966
L37_108 V37 V108 -2.1369885650416828e-11
C37_108 V37 V108 -5.171349735252417e-20

R37_109 V37 V109 -21838.881245235978
L37_109 V37 V109 -1.2111754629407143e-10
C37_109 V37 V109 -5.820660869466069e-20

R37_110 V37 V110 -14239.881389745768
L37_110 V37 V110 -4.283797053276894e-12
C37_110 V37 V110 -1.2272919981415345e-19

R37_111 V37 V111 -58140.86701507894
L37_111 V37 V111 2.668311698814768e-11
C37_111 V37 V111 -7.637738574863047e-21

R37_112 V37 V112 -31592.29459783605
L37_112 V37 V112 5.357493208174159e-12
C37_112 V37 V112 4.475484814112665e-20

R37_113 V37 V113 60364.582120474384
L37_113 V37 V113 1.0885632185493488e-11
C37_113 V37 V113 3.6102460250350967e-20

R37_114 V37 V114 35058.098486611045
L37_114 V37 V114 9.61901882310417e-12
C37_114 V37 V114 6.053694575323812e-20

R37_115 V37 V115 -35410.80084714287
L37_115 V37 V115 -5.894945031463974e-11
C37_115 V37 V115 -1.3334535728739232e-20

R37_116 V37 V116 -562386.4832352505
L37_116 V37 V116 -1.4391307579670386e-11
C37_116 V37 V116 -2.9302599391646756e-20

R37_117 V37 V117 -167047.55681429864
L37_117 V37 V117 -1.094984701550487e-11
C37_117 V37 V117 -4.56818465002931e-20

R37_118 V37 V118 -23721.45859374701
L37_118 V37 V118 -6.205788640510538e-12
C37_118 V37 V118 -8.327340680811669e-20

R37_119 V37 V119 -24522.109856107567
L37_119 V37 V119 -1.1289623839401393e-11
C37_119 V37 V119 -7.04131160197669e-20

R37_120 V37 V120 22670.19382983824
L37_120 V37 V120 -7.467471323107037e-12
C37_120 V37 V120 5.3885292605096516e-21

R37_121 V37 V121 -16458.639247474865
L37_121 V37 V121 5.966147257842515e-12
C37_121 V37 V121 2.087944425928585e-20

R37_122 V37 V122 -13951.167642782195
L37_122 V37 V122 1.0413602890751298e-11
C37_122 V37 V122 -2.0301651829188632e-20

R37_123 V37 V123 -63445.511481225745
L37_123 V37 V123 -1.7983588141772226e-11
C37_123 V37 V123 -2.3049074463002627e-20

R37_124 V37 V124 -29529.407396588187
L37_124 V37 V124 -9.854010508177222e-11
C37_124 V37 V124 9.725831588295509e-21

R37_125 V37 V125 16758.690184886837
L37_125 V37 V125 -5.187028428264265e-12
C37_125 V37 V125 -1.8692862997907792e-20

R37_126 V37 V126 26978.826876340634
L37_126 V37 V126 1.1250409707111906e-10
C37_126 V37 V126 1.1691656861853013e-20

R37_127 V37 V127 371693.3179820729
L37_127 V37 V127 -3.3843368509541605e-11
C37_127 V37 V127 1.5917170451903644e-20

R37_128 V37 V128 30272.281780454534
L37_128 V37 V128 -1.0508747447015538e-10
C37_128 V37 V128 4.894644304515872e-21

R37_129 V37 V129 -36081.78898938638
L37_129 V37 V129 -1.621274711338988e-11
C37_129 V37 V129 -5.109226623705233e-22

R37_130 V37 V130 121972.61925129431
L37_130 V37 V130 5.914772307643625e-11
C37_130 V37 V130 -9.850638216560157e-21

R37_131 V37 V131 38733.21027157663
L37_131 V37 V131 -2.4028376621520813e-10
C37_131 V37 V131 -5.199673293835133e-21

R37_132 V37 V132 115593.76427858368
L37_132 V37 V132 5.743816417045328e-11
C37_132 V37 V132 1.2653006984602021e-20

R37_133 V37 V133 23877.227479592726
L37_133 V37 V133 1.912074986163927e-11
C37_133 V37 V133 6.352721284032765e-20

R37_134 V37 V134 -863089.9746432342
L37_134 V37 V134 -3.731937594526379e-11
C37_134 V37 V134 1.1771932102041555e-20

R37_135 V37 V135 124088.19157947619
L37_135 V37 V135 -2.915715311455184e-11
C37_135 V37 V135 1.270200201612457e-21

R37_136 V37 V136 45310.055079377504
L37_136 V37 V136 -5.4687919436527e-11
C37_136 V37 V136 -2.893516912376423e-21

R37_137 V37 V137 36400.58384103726
L37_137 V37 V137 -7.295328110431926e-12
C37_137 V37 V137 -2.0172436468654856e-21

R37_138 V37 V138 16583.617928106047
L37_138 V37 V138 -7.217685818831121e-11
C37_138 V37 V138 4.67705276717049e-20

R37_139 V37 V139 763926.018322333
L37_139 V37 V139 -3.1218137260923e-11
C37_139 V37 V139 -1.448045124910273e-20

R37_140 V37 V140 273348.8617701351
L37_140 V37 V140 -3.992375652213318e-11
C37_140 V37 V140 -3.250575371004936e-20

R37_141 V37 V141 -94571.2944654177
L37_141 V37 V141 4.108732763987791e-10
C37_141 V37 V141 1.4467883693953822e-20

R37_142 V37 V142 78979.64329916061
L37_142 V37 V142 -3.774511159875586e-11
C37_142 V37 V142 -3.939012628975546e-20

R37_143 V37 V143 3827316.679352134
L37_143 V37 V143 2.193123008396158e-11
C37_143 V37 V143 1.4198234463723994e-20

R37_144 V37 V144 164329.8613896334
L37_144 V37 V144 3.675805495519519e-11
C37_144 V37 V144 4.3580845379360544e-20

R38_38 V38 0 1108.5553211180124
L38_38 V38 0 1.6713315360589603e-12
C38_38 V38 0 5.702363440511644e-20

R38_39 V38 V39 -1957513.0185570526
L38_39 V38 V39 5.159435654419098e-12
C38_39 V38 V39 4.119199897682823e-20

R38_40 V38 V40 -58901.92207840511
L38_40 V38 V40 1.6269502237633337e-11
C38_40 V38 V40 7.042122971829954e-20

R38_41 V38 V41 -16771.284861512588
L38_41 V38 V41 -4.256414665439973e-12
C38_41 V38 V41 -5.402156336546122e-20

R38_42 V38 V42 2755.561841824069
L38_42 V38 V42 8.005963869306785e-13
C38_42 V38 V42 5.1835798228856695e-19

R38_43 V38 V43 -9173.343606220065
L38_43 V38 V43 -1.4538794676487758e-12
C38_43 V38 V43 -2.537624084060778e-19

R38_44 V38 V44 15496.423546529424
L38_44 V38 V44 -4.6824394565656744e-11
C38_44 V38 V44 -1.0271099404920717e-19

R38_45 V38 V45 13204.610225857761
L38_45 V38 V45 2.4786439118063063e-12
C38_45 V38 V45 3.141456115229395e-20

R38_46 V38 V46 -4469.770468108673
L38_46 V38 V46 -1.5367772071966018e-12
C38_46 V38 V46 -3.604773208631924e-19

R38_47 V38 V47 -6022.616574905612
L38_47 V38 V47 -2.919283988327637e-12
C38_47 V38 V47 1.7114251884383524e-19

R38_48 V38 V48 8588.497111093959
L38_48 V38 V48 -1.1423697205585076e-11
C38_48 V38 V48 5.2002349470794414e-20

R38_49 V38 V49 5765.699877941959
L38_49 V38 V49 1.3104236838547003e-11
C38_49 V38 V49 -1.2789201466271833e-20

R38_50 V38 V50 -5960.297091537084
L38_50 V38 V50 -1.1449301253052677e-10
C38_50 V38 V50 8.001875916297152e-20

R38_51 V38 V51 -16662.184076957612
L38_51 V38 V51 -3.2378695358461517e-12
C38_51 V38 V51 -2.2454793073656346e-19

R38_52 V38 V52 -298474.43983768637
L38_52 V38 V52 1.1077952360884738e-11
C38_52 V38 V52 5.656131905129919e-20

R38_53 V38 V53 -12315.243005697885
L38_53 V38 V53 -2.9741972994944558e-12
C38_53 V38 V53 1.8672369223594558e-21

R38_54 V38 V54 221712.6708083363
L38_54 V38 V54 7.340025656987076e-12
C38_54 V38 V54 1.2625208945239727e-19

R38_55 V38 V55 24032.65577006817
L38_55 V38 V55 -5.3835250922943405e-11
C38_55 V38 V55 -1.8807749399397953e-20

R38_56 V38 V56 -6065.100732241424
L38_56 V38 V56 -3.5632388602077563e-12
C38_56 V38 V56 -7.667374804460848e-20

R38_57 V38 V57 -6494.430944395491
L38_57 V38 V57 1.3251934449706454e-11
C38_57 V38 V57 -3.724858205760615e-21

R38_58 V38 V58 13533.621440191495
L38_58 V38 V58 8.000238464471167e-13
C38_58 V38 V58 -1.4571047217634827e-20

R38_59 V38 V59 -2586.90836110795
L38_59 V38 V59 -2.7325853279808284e-12
C38_59 V38 V59 -8.545003700033949e-21

R38_60 V38 V60 17823.391537279058
L38_60 V38 V60 -4.129699496609677e-12
C38_60 V38 V60 -1.3662476747186494e-20

R38_61 V38 V61 21475.31813226012
L38_61 V38 V61 -9.482319506136472e-12
C38_61 V38 V61 2.601355895896622e-20

R38_62 V38 V62 38532.565039836954
L38_62 V38 V62 -8.233588491685053e-12
C38_62 V38 V62 6.20257728777747e-20

R38_63 V38 V63 -10298.683494350169
L38_63 V38 V63 4.684343906645981e-12
C38_63 V38 V63 -6.854638248887435e-20

R38_64 V38 V64 -8317.513512085465
L38_64 V38 V64 -6.498808834828146e-12
C38_64 V38 V64 -5.408122450795268e-20

R38_65 V38 V65 -9529.412823524808
L38_65 V38 V65 -6.458398125412211e-11
C38_65 V38 V65 5.621223795417025e-21

R38_66 V38 V66 -23179.336714084227
L38_66 V38 V66 2.577442376449608e-11
C38_66 V38 V66 1.648946625323577e-20

R38_67 V38 V67 -124823.33702624365
L38_67 V38 V67 -3.542421854586827e-12
C38_67 V38 V67 -3.431732862606236e-20

R38_68 V38 V68 11656.060275183512
L38_68 V38 V68 6.370891161078915e-11
C38_68 V38 V68 -6.227251784518689e-21

R38_69 V38 V69 5631.4834162964835
L38_69 V38 V69 5.022124778658164e-12
C38_69 V38 V69 1.2901946025601882e-21

R38_70 V38 V70 -10278.807231394045
L38_70 V38 V70 -6.6082742169002055e-12
C38_70 V38 V70 -2.8758180639465487e-21

R38_71 V38 V71 -6851.285370491508
L38_71 V38 V71 -4.0640449895876506e-12
C38_71 V38 V71 -1.8082654629238354e-20

R38_72 V38 V72 27664.00519589105
L38_72 V38 V72 9.116425539501462e-12
C38_72 V38 V72 1.1041342230322977e-20

R38_73 V38 V73 11039.77497930547
L38_73 V38 V73 7.855534244103947e-12
C38_73 V38 V73 2.1896622823109115e-20

R38_74 V38 V74 8597.982044499984
L38_74 V38 V74 1.9793191770484523e-11
C38_74 V38 V74 -1.0474701496650508e-20

R38_75 V38 V75 -87825.64755480226
L38_75 V38 V75 -1.0984272398030155e-10
C38_75 V38 V75 -1.1503835347948088e-20

R38_76 V38 V76 41427.72830044907
L38_76 V38 V76 -1.3560537456522506e-11
C38_76 V38 V76 4.259889857491049e-21

R38_77 V38 V77 54289.45026529985
L38_77 V38 V77 -1.1917812598125884e-10
C38_77 V38 V77 1.154399117009256e-21

R38_78 V38 V78 32966.29017367464
L38_78 V38 V78 -1.2466506528348682e-10
C38_78 V38 V78 3.6185403283534484e-20

R38_79 V38 V79 31701.004708198412
L38_79 V38 V79 -7.838379447729294e-12
C38_79 V38 V79 -4.035069373769264e-20

R38_80 V38 V80 -514936.5887312948
L38_80 V38 V80 8.43312375473473e-12
C38_80 V38 V80 3.414117555901408e-20

R38_81 V38 V81 -379677.82022742805
L38_81 V38 V81 2.7917948077283543e-11
C38_81 V38 V81 2.258375056927863e-20

R38_82 V38 V82 392593.045149989
L38_82 V38 V82 -7.871141324536845e-11
C38_82 V38 V82 -5.658073549416452e-20

R38_83 V38 V83 -17323.606358162004
L38_83 V38 V83 -4.136456574273264e-11
C38_83 V38 V83 -3.9117388406860917e-20

R38_84 V38 V84 40825.85597731477
L38_84 V38 V84 -1.934844783141659e-10
C38_84 V38 V84 -1.2289685090004779e-20

R38_85 V38 V85 101444.86235998463
L38_85 V38 V85 -2.2486587167113508e-11
C38_85 V38 V85 -2.752968490914791e-21

R38_86 V38 V86 18304.601238843676
L38_86 V38 V86 1.2669603247704005e-11
C38_86 V38 V86 1.3079736970449933e-20

R38_87 V38 V87 38414.894340870436
L38_87 V38 V87 -1.1776944630327625e-11
C38_87 V38 V87 1.9528313238649528e-20

R38_88 V38 V88 86381.2722613829
L38_88 V38 V88 -3.4092080856612913e-10
C38_88 V38 V88 1.926137427976296e-20

R38_89 V38 V89 2208392.0554271177
L38_89 V38 V89 -7.391702053682342e-11
C38_89 V38 V89 -1.3754279015637082e-20

R38_90 V38 V90 -38301.29965751775
L38_90 V38 V90 6.423487811830684e-12
C38_90 V38 V90 3.8706578368845607e-20

R38_91 V38 V91 -26112.638243780864
L38_91 V38 V91 -8.682640235316352e-11
C38_91 V38 V91 -5.074446833590789e-20

R38_92 V38 V92 -216305.5727225371
L38_92 V38 V92 4.999148384461409e-11
C38_92 V38 V92 -2.3455974305408205e-20

R38_93 V38 V93 44282.78359011122
L38_93 V38 V93 -2.936657629404597e-11
C38_93 V38 V93 2.719114023030737e-21

R38_94 V38 V94 20586.824901632343
L38_94 V38 V94 2.6795895865858165e-11
C38_94 V38 V94 4.1919747225206394e-20

R38_95 V38 V95 -53592.84882916482
L38_95 V38 V95 -1.0905152348403119e-10
C38_95 V38 V95 -3.0075888966231216e-20

R38_96 V38 V96 -43947.61418579142
L38_96 V38 V96 3.969770908368203e-11
C38_96 V38 V96 -2.447302216199877e-20

R38_97 V38 V97 -81148.96555463834
L38_97 V38 V97 6.893119251093554e-12
C38_97 V38 V97 3.86944930883117e-20

R38_98 V38 V98 -26958.11694484824
L38_98 V38 V98 1.489060090430891e-11
C38_98 V38 V98 -1.0282392830972103e-20

R38_99 V38 V99 19726.765592769825
L38_99 V38 V99 -1.164639504985603e-11
C38_99 V38 V99 5.308216575309676e-21

R38_100 V38 V100 295621.596614729
L38_100 V38 V100 4.832223290137194e-11
C38_100 V38 V100 2.0959874636036796e-20

R38_101 V38 V101 167388.27216256625
L38_101 V38 V101 -1.4325254341251923e-10
C38_101 V38 V101 -2.853006300602199e-20

R38_102 V38 V102 59686.63226735719
L38_102 V38 V102 3.001520618751049e-12
C38_102 V38 V102 6.537417599275062e-20

R38_103 V38 V103 -60606.88369855245
L38_103 V38 V103 -4.884725528231872e-12
C38_103 V38 V103 -4.7286420986690376e-20

R38_104 V38 V104 69314.22641221074
L38_104 V38 V104 -3.364159391898757e-09
C38_104 V38 V104 -8.061914292409957e-21

R38_105 V38 V105 106505.92074333929
L38_105 V38 V105 -1.0456464273226496e-11
C38_105 V38 V105 2.9241879796995236e-20

R38_106 V38 V106 239239.22168837013
L38_106 V38 V106 6.992498312528257e-12
C38_106 V38 V106 -3.266436315969698e-20

R38_107 V38 V107 38100.81891740029
L38_107 V38 V107 3.291047797663999e-12
C38_107 V38 V107 4.980398427605188e-20

R38_108 V38 V108 -16953.156645216797
L38_108 V38 V108 -4.155585130618493e-12
C38_108 V38 V108 -3.5259926023760994e-20

R38_109 V38 V109 -59057.93948656267
L38_109 V38 V109 -8.937842041815135e-12
C38_109 V38 V109 -3.7245815241163055e-20

R38_110 V38 V110 -26389.590287878753
L38_110 V38 V110 -7.807157414086971e-11
C38_110 V38 V110 4.96542284096812e-20

R38_111 V38 V111 40077.381403040796
L38_111 V38 V111 -6.1527282086877874e-12
C38_111 V38 V111 -9.179787350920877e-22

R38_112 V38 V112 -23907.529860812152
L38_112 V38 V112 4.372829222207796e-12
C38_112 V38 V112 2.3293729700186916e-20

R38_113 V38 V113 -24772.545986482754
L38_113 V38 V113 1.1019907581795283e-11
C38_113 V38 V113 1.0107779959879302e-20

R38_114 V38 V114 -26948.676591635372
L38_114 V38 V114 1.2127415727687408e-11
C38_114 V38 V114 -3.448580394369808e-20

R38_115 V38 V115 19009927.202831704
L38_115 V38 V115 5.483550144923399e-12
C38_115 V38 V115 3.9968453605463137e-20

R38_116 V38 V116 -1329589.038561195
L38_116 V38 V116 -6.904558634895917e-12
C38_116 V38 V116 -2.7815346130952854e-20

R38_117 V38 V117 -21721.961860310203
L38_117 V38 V117 -1.6649093374030243e-11
C38_117 V38 V117 -2.189361039426788e-20

R38_118 V38 V118 40333.13316654326
L38_118 V38 V118 -1.2120230586230255e-11
C38_118 V38 V118 1.0337670577282163e-20

R38_119 V38 V119 28380.0388848467
L38_119 V38 V119 -9.684386601883144e-12
C38_119 V38 V119 2.452519679614586e-20

R38_120 V38 V120 -6855.81975639067
L38_120 V38 V120 7.960093167783488e-12
C38_120 V38 V120 3.0498382382568707e-21

R38_121 V38 V121 -25820.166252029838
L38_121 V38 V121 3.907941330913427e-11
C38_121 V38 V121 -8.577236848940106e-21

R38_122 V38 V122 -3908.4968715160944
L38_122 V38 V122 4.205977263316563e-12
C38_122 V38 V122 1.1179430016183204e-21

R38_123 V38 V123 -17948.899206552025
L38_123 V38 V123 1.4400157615342574e-11
C38_123 V38 V123 7.892758008987418e-21

R38_124 V38 V124 55869.34241491755
L38_124 V38 V124 -2.9983518428261315e-11
C38_124 V38 V124 1.5122822056619427e-20

R38_125 V38 V125 -94229.62346622864
L38_125 V38 V125 6.449526479067377e-11
C38_125 V38 V125 -4.030422075264451e-21

R38_126 V38 V126 3247.0317482117503
L38_126 V38 V126 -3.4822261895017787e-12
C38_126 V38 V126 -2.1458175775996794e-22

R38_127 V38 V127 -4711.705157564303
L38_127 V38 V127 4.129412141989797e-12
C38_127 V38 V127 1.4742417732590784e-20

R38_128 V38 V128 -76053.70584914359
L38_128 V38 V128 3.3964885961390273e-11
C38_128 V38 V128 1.2078465462332491e-20

R38_129 V38 V129 -12361.814631027093
L38_129 V38 V129 9.517695386421768e-12
C38_129 V38 V129 1.8774176539736886e-20

R38_130 V38 V130 14564.869375780958
L38_130 V38 V130 -6.103160231276859e-12
C38_130 V38 V130 -3.19015777155517e-21

R38_131 V38 V131 9902.364112793155
L38_131 V38 V131 -3.842847494815698e-11
C38_131 V38 V131 4.476513724997361e-21

R38_132 V38 V132 17023.98128577274
L38_132 V38 V132 -1.739133493645035e-11
C38_132 V38 V132 -3.250190590520373e-22

R38_133 V38 V133 60141.98529533389
L38_133 V38 V133 3.333313138189638e-11
C38_133 V38 V133 -5.770256672736534e-21

R38_134 V38 V134 17308.47860337615
L38_134 V38 V134 -3.160559238563354e-11
C38_134 V38 V134 1.0818740809144662e-20

R38_135 V38 V135 -6223.077450286463
L38_135 V38 V135 7.256672833435367e-12
C38_135 V38 V135 -6.041879927373617e-21

R38_136 V38 V136 -478259.7619621074
L38_136 V38 V136 -9.593549090022678e-11
C38_136 V38 V136 -5.107699001112265e-21

R38_137 V38 V137 40996.750674258576
L38_137 V38 V137 -2.737588186719884e-11
C38_137 V38 V137 1.1931645254039164e-20

R38_138 V38 V138 3730.3630278632218
L38_138 V38 V138 -3.589994727485717e-12
C38_138 V38 V138 1.0897657847357969e-20

R38_139 V38 V139 -3483.0859549819584
L38_139 V38 V139 3.0704029782450183e-12
C38_139 V38 V139 1.606965275429383e-21

R38_140 V38 V140 14705.748161389785
L38_140 V38 V140 -8.290945935245595e-12
C38_140 V38 V140 -1.0716102063625969e-20

R38_141 V38 V141 16589.472572297916
L38_141 V38 V141 -1.6028816422025432e-11
C38_141 V38 V141 1.9187133447483593e-21

R38_142 V38 V142 13839.006081375363
L38_142 V38 V142 -9.855878571026916e-12
C38_142 V38 V142 1.2510295042406289e-20

R38_143 V38 V143 10921.012639964369
L38_143 V38 V143 -8.979056495574754e-12
C38_143 V38 V143 -4.5738757009609005e-21

R38_144 V38 V144 -21628.626816840977
L38_144 V38 V144 1.191035704545617e-11
C38_144 V38 V144 1.146442581328194e-20

R39_39 V39 0 -136.04859134349252
L39_39 V39 0 -5.0830143517789784e-14
C39_39 V39 0 -4.389535799547415e-18

R39_40 V39 V40 92367.1600345268
L39_40 V39 V40 5.582446235968725e-12
C39_40 V39 V40 1.994589400693773e-20

R39_41 V39 V41 686.9993937948228
L39_41 V39 V41 2.2277843374606845e-13
C39_41 V39 V41 1.5216344171425803e-18

R39_42 V39 V42 1029.7400784223576
L39_42 V39 V42 3.1145460659281924e-13
C39_42 V39 V42 1.204041060784447e-18

R39_43 V39 V43 1685.4583354831898
L39_43 V39 V43 4.863537440572014e-13
C39_43 V39 V43 8.419434116120186e-19

R39_44 V39 V44 -8412.252806977665
L39_44 V39 V44 -1.4190664171198743e-12
C39_44 V39 V44 -2.7731440619138717e-19

R39_45 V39 V45 -4397.11216222035
L39_45 V39 V45 -3.4123022536673977e-13
C39_45 V39 V45 -1.6614371257153128e-18

R39_46 V39 V46 2632.7383627993795
L39_46 V39 V46 1.213759836941066e-12
C39_46 V39 V46 2.019358435870642e-20

R39_47 V39 V47 4117.524913927744
L39_47 V39 V47 1.2260880760809413e-12
C39_47 V39 V47 -1.0027156553870148e-20

R39_48 V39 V48 -17059.794096406305
L39_48 V39 V48 -2.679987174386467e-12
C39_48 V39 V48 4.602562442758345e-20

R39_49 V39 V49 45184.64971410783
L39_49 V39 V49 5.672727261652678e-12
C39_49 V39 V49 5.270510937763e-19

R39_50 V39 V50 11003.518845548404
L39_50 V39 V50 1.001575157614891e-12
C39_50 V39 V50 2.4066733552302138e-20

R39_51 V39 V51 -4087.6536232527737
L39_51 V39 V51 -1.2017836026873113e-12
C39_51 V39 V51 -2.6109274236939187e-19

R39_52 V39 V52 6565.1799453819085
L39_52 V39 V52 6.469204901895074e-13
C39_52 V39 V52 7.77900081731494e-19

R39_53 V39 V53 17209.172119516385
L39_53 V39 V53 1.1004354186679747e-12
C39_53 V39 V53 3.835855428965798e-19

R39_54 V39 V54 4691.810577182877
L39_54 V39 V54 1.7517471671789898e-12
C39_54 V39 V54 7.934586857671246e-20

R39_55 V39 V55 2318.1844887612083
L39_55 V39 V55 8.265756341103196e-13
C39_55 V39 V55 4.5044315065869825e-19

R39_56 V39 V56 4373.078120207068
L39_56 V39 V56 1.3115627963234093e-12
C39_56 V39 V56 1.8775390621039539e-19

R39_57 V39 V57 430.1618835799758
L39_57 V39 V57 2.2850335984799257e-13
C39_57 V39 V57 -1.6933765833630663e-19

R39_58 V39 V58 2224.0810835790257
L39_58 V39 V58 1.329952937656031e-12
C39_58 V39 V58 -8.802526875247796e-20

R39_59 V39 V59 67836.83268167647
L39_59 V39 V59 1.0617728392272877e-12
C39_59 V39 V59 -1.4951489509809135e-19

R39_60 V39 V60 4545.440988871866
L39_60 V39 V60 1.8818165427475015e-12
C39_60 V39 V60 -2.906126080847203e-20

R39_61 V39 V61 -2256.2046613667685
L39_61 V39 V61 -2.725453651284102e-12
C39_61 V39 V61 5.227934158760057e-19

R39_62 V39 V62 -2199.1894339690743
L39_62 V39 V62 -1.0960173868915231e-11
C39_62 V39 V62 4.76674453177447e-19

R39_63 V39 V63 45315.13843157307
L39_63 V39 V63 5.859799352013952e-12
C39_63 V39 V63 1.2138366206010614e-19

R39_64 V39 V64 -419091.3052464173
L39_64 V39 V64 6.0533128882017806e-12
C39_64 V39 V64 -8.899617084126199e-21

R39_65 V39 V65 1290.1000243814822
L39_65 V39 V65 4.973206531429527e-13
C39_65 V39 V65 1.7725313184642155e-19

R39_66 V39 V66 2002.5258200978856
L39_66 V39 V66 7.366097551279295e-13
C39_66 V39 V66 1.7851650896218527e-19

R39_67 V39 V67 4244.240264304448
L39_67 V39 V67 1.675315024296086e-12
C39_67 V39 V67 1.3078303547775889e-19

R39_68 V39 V68 12526.071114063308
L39_68 V39 V68 1.1409393590995223e-11
C39_68 V39 V68 4.769153317639347e-20

R39_69 V39 V69 -295448.6984957587
L39_69 V39 V69 -1.3413561327337482e-12
C39_69 V39 V69 -1.2114950514112706e-19

R39_70 V39 V70 -14259.861433302207
L39_70 V39 V70 1.2817930275040625e-11
C39_70 V39 V70 -4.133561432125942e-21

R39_71 V39 V71 -89203.52966256905
L39_71 V39 V71 7.301680354669816e-10
C39_71 V39 V71 -1.4348356451157985e-20

R39_72 V39 V72 -44542.086672533726
L39_72 V39 V72 -4.108352815406536e-12
C39_72 V39 V72 -4.217470866040645e-20

R39_73 V39 V73 7405.110804708925
L39_73 V39 V73 6.107097719600426e-12
C39_73 V39 V73 5.108547220113851e-20

R39_74 V39 V74 -18107.101076031922
L39_74 V39 V74 -2.3247292980335755e-12
C39_74 V39 V74 -6.474103371335097e-20

R39_75 V39 V75 8380.871393865711
L39_75 V39 V75 3.001012088960485e-12
C39_75 V39 V75 1.322363926456217e-19

R39_76 V39 V76 11663.972816496846
L39_76 V39 V76 2.8378357521426336e-12
C39_76 V39 V76 8.244192645146786e-20

R39_77 V39 V77 41211.2333039502
L39_77 V39 V77 6.538627323138547e-12
C39_77 V39 V77 2.756494701385023e-20

R39_78 V39 V78 -18031.592809062084
L39_78 V39 V78 -1.8932305754319732e-11
C39_78 V39 V78 -3.371459520939337e-20

R39_79 V39 V79 33371.75938106164
L39_79 V39 V79 -3.172800404397702e-11
C39_79 V39 V79 1.493271993086132e-20

R39_80 V39 V80 -68270.39893761139
L39_80 V39 V80 -2.2975749130860557e-11
C39_80 V39 V80 1.5153446233464618e-20

R39_81 V39 V81 48619.87006242474
L39_81 V39 V81 7.66427592918568e-11
C39_81 V39 V81 1.059289574381645e-21

R39_82 V39 V82 58634.63346150736
L39_82 V39 V82 2.113622212248999e-12
C39_82 V39 V82 2.3928820513715234e-19

R39_83 V39 V83 14431.70426494559
L39_83 V39 V83 2.487184882154262e-12
C39_83 V39 V83 1.5836520751685425e-19

R39_84 V39 V84 14256.835159854669
L39_84 V39 V84 1.6471452815044736e-11
C39_84 V39 V84 -2.2835022554942208e-20

R39_85 V39 V85 346054.57968102786
L39_85 V39 V85 -1.222296467652552e-11
C39_85 V39 V85 -7.209956797300235e-20

R39_86 V39 V86 -46789.20231618418
L39_86 V39 V86 -5.679093144073475e-12
C39_86 V39 V86 -8.902683860963593e-20

R39_87 V39 V87 -31633.198672441642
L39_87 V39 V87 -4.750716651619544e-12
C39_87 V39 V87 -8.390050378208617e-20

R39_88 V39 V88 -30261.22870728056
L39_88 V39 V88 -1.198139400630215e-11
C39_88 V39 V88 5.33285880853707e-21

R39_89 V39 V89 20194.424988824205
L39_89 V39 V89 5.550529771663406e-12
C39_89 V39 V89 1.3923486323363502e-19

R39_90 V39 V90 -103101.23378406452
L39_90 V39 V90 2.713872236646076e-11
C39_90 V39 V90 1.815964972823215e-20

R39_91 V39 V91 14431.712886389114
L39_91 V39 V91 1.92599678121508e-12
C39_91 V39 V91 2.1636487238562973e-19

R39_92 V39 V92 28071.060676283367
L39_92 V39 V92 5.512960714818459e-12
C39_92 V39 V92 6.92375447800479e-20

R39_93 V39 V93 -9394.691681725724
L39_93 V39 V93 -1.237725832461874e-11
C39_93 V39 V93 1.3292395971962308e-20

R39_94 V39 V94 -12645.18861143009
L39_94 V39 V94 -4.3860911728221815e-12
C39_94 V39 V94 -9.386803259774339e-20

R39_95 V39 V95 28029.66696278062
L39_95 V39 V95 3.8702878720323e-12
C39_95 V39 V95 1.1580899468712193e-19

R39_96 V39 V96 47161.88945818394
L39_96 V39 V96 -5.415237905096686e-11
C39_96 V39 V96 3.7295402943842035e-22

R39_97 V39 V97 -20599.367642455112
L39_97 V39 V97 -1.0188037389339007e-11
C39_97 V39 V97 -3.811596860013234e-20

R39_98 V39 V98 -71416.79078374023
L39_98 V39 V98 3.4246943586826545e-12
C39_98 V39 V98 1.0785804510532847e-19

R39_99 V39 V99 -23495.730043022246
L39_99 V39 V99 -3.085295851982969e-11
C39_99 V39 V99 -2.1918655438883605e-20

R39_100 V39 V100 47728.39714171908
L39_100 V39 V100 -2.2526740566608497e-11
C39_100 V39 V100 4.286711435466204e-21

R39_101 V39 V101 250632.941506606
L39_101 V39 V101 3.688326518059669e-12
C39_101 V39 V101 1.4998142207991301e-19

R39_102 V39 V102 68808.72534467903
L39_102 V39 V102 3.785235215254622e-12
C39_102 V39 V102 1.3889533468648035e-19

R39_103 V39 V103 143404.93078404613
L39_103 V39 V103 1.3586183474631166e-11
C39_103 V39 V103 5.801694824688384e-20

R39_104 V39 V104 -537600.2902316836
L39_104 V39 V104 -8.768819578525368e-12
C39_104 V39 V104 -4.899540098588743e-20

R39_105 V39 V105 -297167.80296352913
L39_105 V39 V105 -3.3047486815853505e-12
C39_105 V39 V105 -1.2173969442956342e-19

R39_106 V39 V106 7933.96754921405
L39_106 V39 V106 2.2453047827480106e-12
C39_106 V39 V106 2.0642175291055247e-19

R39_107 V39 V107 650702.1303390859
L39_107 V39 V107 6.1539758643134215e-12
C39_107 V39 V107 6.418294589974059e-20

R39_108 V39 V108 -27839.112779447456
L39_108 V39 V108 -6.306782114708411e-12
C39_108 V39 V108 -1.0735689707687411e-19

R39_109 V39 V109 -33238.97440904525
L39_109 V39 V109 -1.1280652275116576e-11
C39_109 V39 V109 -9.76881701201773e-20

R39_110 V39 V110 -16125.349684663477
L39_110 V39 V110 -2.204332872662675e-12
C39_110 V39 V110 -2.435779652084526e-19

R39_111 V39 V111 62781.83792496182
L39_111 V39 V111 -1.2323817180639985e-11
C39_111 V39 V111 -4.783306495873904e-20

R39_112 V39 V112 12945.943544947479
L39_112 V39 V112 3.117217467497299e-12
C39_112 V39 V112 1.051915430590993e-19

R39_113 V39 V113 24865.53631329286
L39_113 V39 V113 5.770007253171171e-12
C39_113 V39 V113 7.679742793169478e-20

R39_114 V39 V114 14989.48861384286
L39_114 V39 V114 4.03386468339783e-12
C39_114 V39 V114 1.2962033049189008e-19

R39_115 V39 V115 -47104.10216646432
L39_115 V39 V115 1.253332086683022e-11
C39_115 V39 V115 7.32507090548882e-21

R39_116 V39 V116 -25471.071377340617
L39_116 V39 V116 -7.989454082210834e-12
C39_116 V39 V116 -6.228561193328003e-20

R39_117 V39 V117 -14627.088586909273
L39_117 V39 V117 -6.280409613514636e-12
C39_117 V39 V117 -8.563013553817646e-20

R39_118 V39 V118 -97478.13637886762
L39_118 V39 V118 -4.008691357264936e-12
C39_118 V39 V118 -1.170192729263338e-19

R39_119 V39 V119 -108233.66198331716
L39_119 V39 V119 -4.517446268437164e-12
C39_119 V39 V119 -1.1633985971965073e-19

R39_120 V39 V120 -20031.772352928612
L39_120 V39 V120 -9.331767614678213e-12
C39_120 V39 V120 -1.1956017678109805e-20

R39_121 V39 V121 16883.227947070314
L39_121 V39 V121 5.4149883560651334e-12
C39_121 V39 V121 2.6408230892755328e-20

R39_122 V39 V122 11417.582834041983
L39_122 V39 V122 6.697194777796448e-12
C39_122 V39 V122 -1.4771761111555086e-20

R39_123 V39 V123 44600.10892160847
L39_123 V39 V123 -1.8488173838061367e-11
C39_123 V39 V123 -4.6321882773186554e-20

R39_124 V39 V124 25084.0171143333
L39_124 V39 V124 -2.07680838711219e-11
C39_124 V39 V124 -9.586354946188994e-21

R39_125 V39 V125 -11093.329754660388
L39_125 V39 V125 -6.113949116479476e-12
C39_125 V39 V125 -2.1143084331018365e-20

R39_126 V39 V126 -15581.31637040969
L39_126 V39 V126 -2.3492242696396914e-11
C39_126 V39 V126 1.8856583206611567e-20

R39_127 V39 V127 1587317.3215841954
L39_127 V39 V127 2.4464628066756375e-11
C39_127 V39 V127 7.313425953976106e-21

R39_128 V39 V128 -17968.76204154779
L39_128 V39 V128 4.2897774737752575e-11
C39_128 V39 V128 -1.2147666881984307e-20

R39_129 V39 V129 55112.274629713735
L39_129 V39 V129 -3.4791976663332263e-11
C39_129 V39 V129 -3.0998836196775e-20

R39_130 V39 V130 -10923.428440728583
L39_130 V39 V130 -2.728437368830007e-11
C39_130 V39 V130 -3.124869614647732e-20

R39_131 V39 V131 -13501.634581397886
L39_131 V39 V131 4.23854655749958e-11
C39_131 V39 V131 1.5837890037161028e-20

R39_132 V39 V132 1160672.0294228955
L39_132 V39 V132 -1.0009656190322271e-10
C39_132 V39 V132 -4.892303445158593e-21

R39_133 V39 V133 45233.877193108216
L39_133 V39 V133 9.347729177223433e-12
C39_133 V39 V133 6.579045199431686e-20

R39_134 V39 V134 19422.175486913227
L39_134 V39 V134 -9.509156583003883e-11
C39_134 V39 V134 1.7823827262303475e-20

R39_135 V39 V135 33478.41122464454
L39_135 V39 V135 -1.6456665348833428e-10
C39_135 V39 V135 -4.86876316586384e-21

R39_136 V39 V136 -26136.929705745177
L39_136 V39 V136 3.5625457794092077e-10
C39_136 V39 V136 8.93062520706216e-21

R39_137 V39 V137 -13345.314281241714
L39_137 V39 V137 -6.800107479684703e-12
C39_137 V39 V137 -1.661564132835892e-20

R39_138 V39 V138 -13297.642358578338
L39_138 V39 V138 -1.0520425476321588e-11
C39_138 V39 V138 1.0342612667777062e-20

R39_139 V39 V139 -31617.44153638176
L39_139 V39 V139 1.9901082025846885e-11
C39_139 V39 V139 -1.3782731547408987e-20

R39_140 V39 V140 178806.82257775567
L39_140 V39 V140 -2.980936834339524e-11
C39_140 V39 V140 -2.0907101567639018e-20

R39_141 V39 V141 -84983.13716694893
L39_141 V39 V141 -2.5549014521847208e-11
C39_141 V39 V141 -2.9041983205803393e-21

R39_142 V39 V142 -38133.80499500371
L39_142 V39 V142 -7.720536194572763e-12
C39_142 V39 V142 -5.903781419312766e-20

R39_143 V39 V143 -87040.26786434613
L39_143 V39 V143 4.442570053829891e-11
C39_143 V39 V143 7.100290860461377e-21

R39_144 V39 V144 14505.692155326378
L39_144 V39 V144 1.3882424145526244e-11
C39_144 V39 V144 4.8982716242102097e-20

R40_40 V40 0 -5800.180042767919
L40_40 V40 0 -1.5406236242993928e-13
C40_40 V40 0 -1.4737472059869668e-18

R40_41 V40 V41 16022.2005594443
L40_41 V40 V41 2.3467613039548474e-12
C40_41 V40 V41 1.9819145447399237e-19

R40_42 V40 V42 665191.4334489903
L40_42 V40 V42 -1.1932357837754448e-11
C40_42 V40 V42 1.447576738332968e-20

R40_43 V40 V43 -213209.7845403652
L40_43 V40 V43 -1.5647818603194907e-11
C40_43 V40 V43 3.2515805851880033e-20

R40_44 V40 V44 1505.0363234178212
L40_44 V40 V44 3.743032128922804e-13
C40_44 V40 V44 1.1476987155430463e-18

R40_45 V40 V45 -5775.356074411326
L40_45 V40 V45 -1.4385237573856933e-12
C40_45 V40 V45 -4.839936407865203e-19

R40_46 V40 V46 -432275.01170136756
L40_46 V40 V46 3.302643223376246e-12
C40_46 V40 V46 2.2425955702885103e-19

R40_47 V40 V47 -7865.1505772694
L40_47 V40 V47 7.434442898063943e-12
C40_47 V40 V47 -6.49150339485341e-21

R40_48 V40 V48 220614.34445299255
L40_48 V40 V48 3.935456729361886e-12
C40_48 V40 V48 -2.561456812956195e-19

R40_49 V40 V49 5190.309159118118
L40_49 V40 V49 7.605345938113192e-12
C40_49 V40 V49 7.773665558036033e-20

R40_50 V40 V50 -5530.4423298567135
L40_50 V40 V50 -5.061455062744043e-11
C40_50 V40 V50 4.0433911724387777e-20

R40_51 V40 V51 15836.778614677263
L40_51 V40 V51 8.576135488984938e-12
C40_51 V40 V51 -3.186500990234949e-20

R40_52 V40 V52 33008.58327378795
L40_52 V40 V52 5.1848375828893984e-12
C40_52 V40 V52 2.450310154178558e-19

R40_53 V40 V53 -6929.1205552646625
L40_53 V40 V53 -3.312020230823929e-12
C40_53 V40 V53 -2.522688163092518e-19

R40_54 V40 V54 -11203.435874573
L40_54 V40 V54 -1.7092060824420785e-11
C40_54 V40 V54 -8.832778953962605e-20

R40_55 V40 V55 62471.00407154338
L40_55 V40 V55 1.6036159973698012e-11
C40_55 V40 V55 4.5103665451598745e-20

R40_56 V40 V56 5735.54919789663
L40_56 V40 V56 1.1603212335015539e-12
C40_56 V40 V56 6.555307026977717e-19

R40_57 V40 V57 -3771.8211253651016
L40_57 V40 V57 5.120170503290402e-12
C40_57 V40 V57 1.6847572929400122e-20

R40_58 V40 V58 -17423.71147171301
L40_58 V40 V58 -3.953648976636459e-12
C40_58 V40 V58 -4.1451221934923986e-20

R40_59 V40 V59 -3426.740630830508
L40_59 V40 V59 -5.768511388593374e-12
C40_59 V40 V59 -2.4534778247608833e-20

R40_60 V40 V60 3838.657194498179
L40_60 V40 V60 4.2851018939103804e-13
C40_60 V40 V60 -5.552333064695602e-20

R40_61 V40 V61 11103.648818763928
L40_61 V40 V61 -7.458111116059125e-12
C40_61 V40 V61 1.9390536021103074e-20

R40_62 V40 V62 11390.65809896976
L40_62 V40 V62 3.336402771286397e-12
C40_62 V40 V62 3.4193222959805926e-20

R40_63 V40 V63 22165.124579864332
L40_63 V40 V63 4.826143166640497e-12
C40_63 V40 V63 7.076423806496399e-20

R40_64 V40 V64 16890.36033926734
L40_64 V40 V64 5.322874491795573e-12
C40_64 V40 V64 2.9779822911882714e-19

R40_65 V40 V65 -5964.224884322025
L40_65 V40 V65 1.2618636169843895e-11
C40_65 V40 V65 -1.6636048635374326e-20

R40_66 V40 V66 -9328.92914520108
L40_66 V40 V66 -1.942832646348343e-11
C40_66 V40 V66 7.838634777838914e-20

R40_67 V40 V67 40626.59671817842
L40_67 V40 V67 7.204187628669873e-12
C40_67 V40 V67 7.214528617725261e-20

R40_68 V40 V68 5213.004598142344
L40_68 V40 V68 8.251778273004187e-13
C40_68 V40 V68 1.0998256549140076e-19

R40_69 V40 V69 11538.776935752354
L40_69 V40 V69 -2.033154489793223e-12
C40_69 V40 V69 -8.605959712117425e-20

R40_70 V40 V70 -100572.73073345497
L40_70 V40 V70 7.716609283333205e-12
C40_70 V40 V70 -4.719922756959615e-21

R40_71 V40 V71 -18155.79533312503
L40_71 V40 V71 -1.9014222708921307e-11
C40_71 V40 V71 -1.874000827826544e-20

R40_72 V40 V72 20633.68324589205
L40_72 V40 V72 -2.640231995238902e-11
C40_72 V40 V72 2.779074004159212e-20

R40_73 V40 V73 11578.99937292804
L40_73 V40 V73 3.952691660082184e-12
C40_73 V40 V73 -3.366662783178202e-20

R40_74 V40 V74 12351.131609020704
L40_74 V40 V74 2.4543034707976585e-08
C40_74 V40 V74 -3.989209783939919e-21

R40_75 V40 V75 -126407.36555747096
L40_75 V40 V75 -4.500147508418185e-11
C40_75 V40 V75 7.912342813159051e-20

R40_76 V40 V76 -33229.99666541368
L40_76 V40 V76 -1.6477416705990806e-11
C40_76 V40 V76 -1.8310209579571178e-20

R40_77 V40 V77 -106952.67929729822
L40_77 V40 V77 -6.049288055125434e-11
C40_77 V40 V77 2.6435747336135636e-20

R40_78 V40 V78 -209345.50439610318
L40_78 V40 V78 -2.4422755198393507e-11
C40_78 V40 V78 -3.354267840887423e-20

R40_79 V40 V79 48220.92767104246
L40_79 V40 V79 -3.875447356587761e-11
C40_79 V40 V79 -4.145273694542193e-20

R40_80 V40 V80 24979.95186638899
L40_80 V40 V80 5.289941532245184e-12
C40_80 V40 V80 1.2380622277854472e-19

R40_81 V40 V81 -23081.443235384857
L40_81 V40 V81 -3.2577972533870834e-12
C40_81 V40 V81 -1.5822604359817195e-19

R40_82 V40 V82 72487.61961529891
L40_82 V40 V82 2.2530702757310508e-11
C40_82 V40 V82 4.253629148728022e-20

R40_83 V40 V83 60894.319591442814
L40_83 V40 V83 6.500666130266354e-12
C40_83 V40 V83 9.81570024329237e-20

R40_84 V40 V84 89536.43493658304
L40_84 V40 V84 1.28317533836249e-11
C40_84 V40 V84 2.0369346858400716e-20

R40_85 V40 V85 119213.62739291103
L40_85 V40 V85 -2.4778790682223715e-11
C40_85 V40 V85 -5.486465133701087e-20

R40_86 V40 V86 20552.26493065805
L40_86 V40 V86 3.636575630973424e-10
C40_86 V40 V86 1.3511270007733165e-23

R40_87 V40 V87 -86658.35825810413
L40_87 V40 V87 -1.7627732543296095e-11
C40_87 V40 V87 -3.041291190672061e-20

R40_88 V40 V88 -45926.429152030156
L40_88 V40 V88 -1.2473120318021747e-11
C40_88 V40 V88 -3.4864796351378666e-20

R40_89 V40 V89 142363.29659848372
L40_89 V40 V89 1.3366414936701118e-11
C40_89 V40 V89 5.1776463239882413e-20

R40_90 V40 V90 92424.46913187046
L40_90 V40 V90 3.7372590335589816e-11
C40_90 V40 V90 5.050962802701711e-20

R40_91 V40 V91 -332756.0776907527
L40_91 V40 V91 3.8896890123123623e-10
C40_91 V40 V91 1.97748511540765e-20

R40_92 V40 V92 14985.388209254214
L40_92 V40 V92 3.601775873354107e-12
C40_92 V40 V92 1.6048800562560017e-19

R40_93 V40 V93 53088.05494678646
L40_93 V40 V93 -2.487128796907425e-11
C40_93 V40 V93 -1.4309588540585133e-20

R40_94 V40 V94 -36097.38437954896
L40_94 V40 V94 -6.777956267614217e-12
C40_94 V40 V94 -8.631123662982767e-20

R40_95 V40 V95 441331.49520851305
L40_95 V40 V95 1.058371315827806e-10
C40_95 V40 V95 2.0003078781948954e-20

R40_96 V40 V96 21209.622255587943
L40_96 V40 V96 3.2854329902268507e-12
C40_96 V40 V96 1.6627863236906438e-19

R40_97 V40 V97 190720.76973578957
L40_97 V40 V97 -1.602048466911033e-11
C40_97 V40 V97 -2.053300018180018e-20

R40_98 V40 V98 36039.95103024821
L40_98 V40 V98 7.875807989073128e-12
C40_98 V40 V98 6.145988344886247e-20

R40_99 V40 V99 -81343.86269475697
L40_99 V40 V99 -2.7210499139744374e-11
C40_99 V40 V99 -3.398909290616599e-20

R40_100 V40 V100 -23237.543267004992
L40_100 V40 V100 -1.0458403055130514e-11
C40_100 V40 V100 -7.875481883987205e-20

R40_101 V40 V101 45168.26887957184
L40_101 V40 V101 8.688490829569477e-12
C40_101 V40 V101 7.28747734073249e-20

R40_102 V40 V102 25586.6956733621
L40_102 V40 V102 2.108958409406661e-11
C40_102 V40 V102 6.208906140656974e-20

R40_103 V40 V103 113132.83994047658
L40_103 V40 V103 -8.188276389207822e-11
C40_103 V40 V103 -4.421854044992032e-20

R40_104 V40 V104 16518.4580559114
L40_104 V40 V104 3.598285154695377e-12
C40_104 V40 V104 1.9557383646488803e-19

R40_105 V40 V105 -15051.566121700751
L40_105 V40 V105 -5.642232878992031e-12
C40_105 V40 V105 -1.5196914920031994e-19

R40_106 V40 V106 26018.953524773126
L40_106 V40 V106 6.668123534860794e-12
C40_106 V40 V106 1.5236758615585922e-19

R40_107 V40 V107 67335.12806432156
L40_107 V40 V107 1.9330127593903846e-11
C40_107 V40 V107 6.564977052960934e-20

R40_108 V40 V108 -16687.79891566802
L40_108 V40 V108 -7.405700032357075e-12
C40_108 V40 V108 -1.3923189967900761e-19

R40_109 V40 V109 15887.077961593997
L40_109 V40 V109 5.643274648595242e-12
C40_109 V40 V109 1.5196739174870525e-19

R40_110 V40 V110 -75442.98751193658
L40_110 V40 V110 -7.632873845791863e-12
C40_110 V40 V110 -1.0895655067671104e-19

R40_111 V40 V111 -38615.77692781693
L40_111 V40 V111 -3.18575109425746e-11
C40_111 V40 V111 -5.334357911453346e-20

R40_112 V40 V112 30166.260014568496
L40_112 V40 V112 1.675420937453907e-11
C40_112 V40 V112 4.790020751945473e-20

R40_113 V40 V113 -22007.306167158626
L40_113 V40 V113 3.9582478631598865e-11
C40_113 V40 V113 -4.026001288226595e-21

R40_114 V40 V114 17350.401961490224
L40_114 V40 V114 9.273569872289948e-11
C40_114 V40 V114 2.6125340896670887e-20

R40_115 V40 V115 30492.367367851108
L40_115 V40 V115 4.813135846465809e-11
C40_115 V40 V115 3.7018970300417676e-20

R40_116 V40 V116 -27976.644632398016
L40_116 V40 V116 -1.0232976563501458e-11
C40_116 V40 V116 -7.002239193805384e-20

R40_117 V40 V117 41179.12721355172
L40_117 V40 V117 -1.8967278639327455e-11
C40_117 V40 V117 -3.143660832303123e-20

R40_118 V40 V118 3343563.893252558
L40_118 V40 V118 -4.226449139050691e-11
C40_118 V40 V118 -2.25053265652973e-20

R40_119 V40 V119 -13918.445429827512
L40_119 V40 V119 -1.655992351915063e-11
C40_119 V40 V119 -6.158931513804492e-20

R40_120 V40 V120 263704.21467666386
L40_120 V40 V120 -1.5560763493415652e-11
C40_120 V40 V120 -4.5758861779780814e-20

R40_121 V40 V121 -4483420.999291257
L40_121 V40 V121 5.0871258002054216e-11
C40_121 V40 V121 1.2550561267081134e-20

R40_122 V40 V122 34736.08953810531
L40_122 V40 V122 9.516892031685769e-11
C40_122 V40 V122 1.3575558895346414e-20

R40_123 V40 V123 18694.35772834318
L40_123 V40 V123 -1.9839141322044672e-10
C40_123 V40 V123 4.952513643903566e-21

R40_124 V40 V124 79969.7248901227
L40_124 V40 V124 -1.988389904712829e-11
C40_124 V40 V124 -7.936213066697972e-20

R40_125 V40 V125 27529.616911029912
L40_125 V40 V125 -1.7488453642833465e-11
C40_125 V40 V125 -7.454184095781877e-21

R40_126 V40 V126 -27294.64284506409
L40_126 V40 V126 3.8527232273489744e-11
C40_126 V40 V126 3.6352947530628103e-22

R40_127 V40 V127 69371.35422366149
L40_127 V40 V127 -1.0826912686422849e-10
C40_127 V40 V127 -1.5632545279140474e-20

R40_128 V40 V128 -56111.909608147886
L40_128 V40 V128 -1.1844045372966151e-11
C40_128 V40 V128 -5.115798837887724e-20

R40_129 V40 V129 15785.859129061653
L40_129 V40 V129 -3.46011540834794e-11
C40_129 V40 V129 -3.032092241450605e-20

R40_130 V40 V130 -13035.624217780012
L40_130 V40 V130 -1.2192032434872635e-11
C40_130 V40 V130 -7.932436707488567e-20

R40_131 V40 V131 -19960.501421615743
L40_131 V40 V131 -1.347056271567294e-10
C40_131 V40 V131 1.274290291101786e-21

R40_132 V40 V132 -46836.33126344825
L40_132 V40 V132 -1.1858365166018924e-11
C40_132 V40 V132 -4.3370388665955003e-20

R40_133 V40 V133 -1469753.9954045552
L40_133 V40 V133 1.3597005807415746e-11
C40_133 V40 V133 6.549883667600194e-20

R40_134 V40 V134 -173389.57163193653
L40_134 V40 V134 -1.0059298792605505e-10
C40_134 V40 V134 -1.4266433280423083e-21

R40_135 V40 V135 114729.48959691642
L40_135 V40 V135 -3.0223946201497355e-11
C40_135 V40 V135 -2.6836571065519346e-20

R40_136 V40 V136 -68663.24542791508
L40_136 V40 V136 1.5367169953106532e-11
C40_136 V40 V136 4.69725790823229e-20

R40_137 V40 V137 89965.2510541432
L40_137 V40 V137 -2.365297762196526e-11
C40_137 V40 V137 -5.811817768799623e-20

R40_138 V40 V138 -11955.162255767927
L40_138 V40 V138 1.6826751102207493e-11
C40_138 V40 V138 3.402432957078248e-21

R40_139 V40 V139 26578.49870375687
L40_139 V40 V139 1.0677600836047349e-10
C40_139 V40 V139 3.494446364303769e-20

R40_140 V40 V140 -32709.924995363283
L40_140 V40 V140 -8.138117177585792e-11
C40_140 V40 V140 1.2556831954293643e-20

R40_141 V40 V141 26465.991996072346
L40_141 V40 V141 1.3049056174781132e-11
C40_141 V40 V141 4.1547774757319676e-20

R40_142 V40 V142 -10196.68280868557
L40_142 V40 V142 -1.0252532999276624e-10
C40_142 V40 V142 -2.8409638861048616e-20

R40_143 V40 V143 -23802.772124716714
L40_143 V40 V143 -1.8530152472119693e-10
C40_143 V40 V143 -1.8788783649102974e-20

R40_144 V40 V144 -60614.02831224319
L40_144 V40 V144 -4.144658705584011e-11
C40_144 V40 V144 -5.60493196693307e-20

R41_41 V41 0 28.345120995990737
L41_41 V41 0 1.2005468008971494e-14
C41_41 V41 0 1.6657962186053675e-17

R41_42 V41 V42 -273.30314243537356
L41_42 V41 V42 -7.503218291662258e-14
C41_42 V41 V42 -4.491533254251016e-18

R41_43 V41 V43 -489.6892729638458
L41_43 V41 V43 -1.3777547652956036e-13
C41_43 V41 V43 -2.508997082731321e-18

R41_44 V41 V44 -2595.699759436652
L41_44 V41 V44 -7.429667011510104e-13
C41_44 V41 V44 -3.905878453775551e-19

R41_45 V41 V45 -53246.57220837672
L41_45 V41 V45 1.4741240449269106e-13
C41_45 V41 V45 4.8710487248257724e-18

R41_46 V41 V46 -1367.3779795006687
L41_46 V41 V46 6.64246699422355e-13
C41_46 V41 V46 2.2633735360592677e-18

R41_47 V41 V47 -1215.2569227962013
L41_47 V41 V47 -3.2656696222777724e-12
C41_47 V41 V47 9.277826502876348e-19

R41_48 V41 V48 4499.681718138094
L41_48 V41 V48 1.0777029181398774e-12
C41_48 V41 V48 2.918764366814437e-19

R41_49 V41 V49 -37728.772977014996
L41_49 V41 V49 -7.934053142974496e-13
C41_49 V41 V49 -1.1774580904129064e-18

R41_50 V41 V50 -1012.504581694435
L41_50 V41 V50 -2.935630160272511e-13
C41_50 V41 V50 -1.1346348869882048e-18

R41_51 V41 V51 935.3892298837897
L41_51 V41 V51 3.500896227431891e-13
C41_51 V41 V51 7.124091528603481e-19

R41_52 V41 V52 -903.8462046948455
L41_52 V41 V52 -1.6157322319602443e-13
C41_52 V41 V52 -3.2084277007226716e-18

R41_53 V41 V53 -941.6996290425668
L41_53 V41 V53 -2.333806637262889e-13
C41_53 V41 V53 -1.755690737833756e-18

R41_54 V41 V54 -888.0426593542609
L41_54 V41 V54 -4.743998192847319e-13
C41_54 V41 V54 -1.877500137866448e-19

R41_55 V41 V55 -570.7501797424079
L41_55 V41 V55 -2.4273991987368865e-13
C41_55 V41 V55 -9.520709527325893e-19

R41_56 V41 V56 -927.8478338979696
L41_56 V41 V56 -3.1094034149995714e-13
C41_56 V41 V56 -9.840684544899257e-19

R41_57 V41 V57 -95.60089768625436
L41_57 V41 V57 -5.419503240259144e-14
C41_57 V41 V57 6.416081462638085e-19

R41_58 V41 V58 -537.9976344173812
L41_58 V41 V58 -3.386581994150934e-13
C41_58 V41 V58 3.344918906429457e-19

R41_59 V41 V59 5159.507946730527
L41_59 V41 V59 1.967868487383994e-12
C41_59 V41 V59 4.419329478028761e-19

R41_60 V41 V60 -566.7198874566527
L41_60 V41 V60 -3.0797930818981686e-13
C41_60 V41 V60 1.1446294372739193e-19

R41_61 V41 V61 547.1848329952085
L41_61 V41 V61 1.4592476094146122e-12
C41_61 V41 V61 -2.2108496522845656e-18

R41_62 V41 V62 444.72661478868014
L41_62 V41 V62 5.859587060729437e-13
C41_62 V41 V62 -1.74599255633976e-18

R41_63 V41 V63 4320.432411486005
L41_63 V41 V63 -1.9808451093343636e-12
C41_63 V41 V63 -5.229564183459715e-19

R41_64 V41 V64 -4378.220999180524
L41_64 V41 V64 -1.2978843008360516e-12
C41_64 V41 V64 -3.5921866545211747e-19

R41_65 V41 V65 -215.9049548559424
L41_65 V41 V65 -1.2118451173731347e-13
C41_65 V41 V65 -6.593841340502958e-19

R41_66 V41 V66 -240.64425924938178
L41_66 V41 V66 -1.4537007003527866e-13
C41_66 V41 V66 -5.2093673797977965e-19

R41_67 V41 V67 -959.7463987538886
L41_67 V41 V67 -4.951835536412379e-13
C41_67 V41 V67 -4.0106794088292164e-19

R41_68 V41 V68 -1859.8205066225373
L41_68 V41 V68 -6.372524551800756e-13
C41_68 V41 V68 -2.316853099466668e-19

R41_69 V41 V69 2573.8960792872463
L41_69 V41 V69 1.020465551802528e-12
C41_69 V41 V69 1.4185465219513114e-19

R41_70 V41 V70 1185.539379902779
L41_70 V41 V70 1.0577542435127558e-11
C41_70 V41 V70 -3.3132845943606844e-19

R41_71 V41 V71 13072.199952981615
L41_71 V41 V71 -4.713262894532168e-12
C41_71 V41 V71 -1.315295443675739e-19

R41_72 V41 V72 817.6029166535548
L41_72 V41 V72 7.570103431539186e-13
C41_72 V41 V72 -6.253222581586773e-20

R41_73 V41 V73 -20872.89274282897
L41_73 V41 V73 -1.2025943489306119e-12
C41_73 V41 V73 -2.9060740537166267e-19

R41_74 V41 V74 1314.076614286867
L41_74 V41 V74 6.44761506597349e-13
C41_74 V41 V74 2.945396976373128e-19

R41_75 V41 V75 -1055.4645437658887
L41_75 V41 V75 -7.301095794504771e-13
C41_75 V41 V75 -1.8627926783387412e-19

R41_76 V41 V76 -1100.1208617937239
L41_76 V41 V76 -4.851548493848137e-13
C41_76 V41 V76 -4.1949034891108107e-19

R41_77 V41 V77 -3507.4076787629597
L41_77 V41 V77 -1.4302869595262251e-12
C41_77 V41 V77 -9.94518947738404e-20

R41_78 V41 V78 -15701.83889520307
L41_78 V41 V78 -2.1026263015686254e-12
C41_78 V41 V78 -2.0782754610391596e-19

R41_79 V41 V79 6529.474319369285
L41_79 V41 V79 -3.280836733296095e-11
C41_79 V41 V79 -1.9972201369640016e-19

R41_80 V41 V80 3265.8891346594432
L41_80 V41 V80 1.6178146828278747e-12
C41_80 V41 V80 1.6539811621829811e-19

R41_81 V41 V81 7351.966964948262
L41_81 V41 V81 5.205195262008724e-12
C41_81 V41 V81 7.39457441209294e-20

R41_82 V41 V82 7513.144042163195
L41_82 V41 V82 1.832156976514597e-12
C41_82 V41 V82 3.1025156356738143e-19

R41_83 V41 V83 13867.397884091668
L41_83 V41 V83 1.002779024015916e-11
C41_83 V41 V83 2.0451164262783066e-19

R41_84 V41 V84 31099.92842871111
L41_84 V41 V84 -3.223200252150346e-12
C41_84 V41 V84 -4.344235960675627e-20

R41_85 V41 V85 4717.033687044853
L41_85 V41 V85 -3.161607573705764e-12
C41_85 V41 V85 -1.4585626046230277e-19

R41_86 V41 V86 13829.64558951874
L41_86 V41 V86 -4.5964698867590696e-12
C41_86 V41 V86 -8.373702403531772e-20

R41_87 V41 V87 -6454.409813926607
L41_87 V41 V87 -3.347062786680568e-12
C41_87 V41 V87 -2.0715954168530973e-19

R41_88 V41 V88 -90101.70675387283
L41_88 V41 V88 1.4051071704664684e-11
C41_88 V41 V88 -5.555414294516384e-20

R41_89 V41 V89 -7204.110983914789
L41_89 V41 V89 3.421872577095624e-12
C41_89 V41 V89 5.921389225474582e-20

R41_90 V41 V90 21348.88706904845
L41_90 V41 V90 4.41324968829081e-12
C41_90 V41 V90 1.3494252673606259e-19

R41_91 V41 V91 6523.050617378451
L41_91 V41 V91 3.0206908489376366e-12
C41_91 V41 V91 2.750315543713388e-19

R41_92 V41 V92 258133.5026676215
L41_92 V41 V92 1.988007503503811e-11
C41_92 V41 V92 8.575407635171716e-20

R41_93 V41 V93 1781.8038330100494
L41_93 V41 V93 1.6570024306366417e-11
C41_93 V41 V93 -2.847505212503878e-20

R41_94 V41 V94 4843.997361853806
L41_94 V41 V94 -2.952525969549802e-11
C41_94 V41 V94 -4.7760027289888185e-20

R41_95 V41 V95 15113.204930060805
L41_95 V41 V95 5.610087681934494e-12
C41_95 V41 V95 1.8797730758263724e-19

R41_96 V41 V96 -10706.624959109215
L41_96 V41 V96 -4.9179794842421444e-11
C41_96 V41 V96 8.91463605103581e-20

R41_97 V41 V97 3377.5785410293133
L41_97 V41 V97 1.3888786174168961e-11
C41_97 V41 V97 9.640536734773467e-21

R41_98 V41 V98 2531.5754385886567
L41_98 V41 V98 6.656036144847023e-12
C41_98 V41 V98 1.1248885565155871e-19

R41_99 V41 V99 6321.743327731739
L41_99 V41 V99 -1.1409715603208402e-11
C41_99 V41 V99 -2.872083698613011e-20

R41_100 V41 V100 -14609.735992549367
L41_100 V41 V100 1.9605536823163286e-11
C41_100 V41 V100 1.5042888852899567e-20

R41_101 V41 V101 4170.634359200671
L41_101 V41 V101 7.117777214138386e-12
C41_101 V41 V101 4.5316037379827206e-20

R41_102 V41 V102 3976.321190508458
L41_102 V41 V102 2.306338577319566e-12
C41_102 V41 V102 2.454493300790846e-19

R41_103 V41 V103 36972.67142916854
L41_103 V41 V103 -8.93317896213848e-12
C41_103 V41 V103 -2.3192246585136417e-19

R41_104 V41 V104 -22328.22594955606
L41_104 V41 V104 -9.860478167215645e-12
C41_104 V41 V104 4.11452718506889e-21

R41_105 V41 V105 -3199.120112638822
L41_105 V41 V105 -5.214041370152883e-12
C41_105 V41 V105 -1.1830708817338357e-19

R41_106 V41 V106 -6980.852376522548
L41_106 V41 V106 2.713708131204878e-12
C41_106 V41 V106 3.886514545581972e-19

R41_107 V41 V107 4699.681416887644
L41_107 V41 V107 2.9761165823754664e-12
C41_107 V41 V107 3.0874208588223057e-19

R41_108 V41 V108 -29888.65435629369
L41_108 V41 V108 -3.96670526230345e-12
C41_108 V41 V108 -8.65732583884494e-20

R41_109 V41 V109 38319.71560534915
L41_109 V41 V109 -4.4606799131765355e-12
C41_109 V41 V109 -7.010113876841504e-20

R41_110 V41 V110 -5877.676348663597
L41_110 V41 V110 -2.902274695894464e-12
C41_110 V41 V110 -2.9251676332144335e-19

R41_111 V41 V111 -5860.093796566463
L41_111 V41 V111 -4.608256361622461e-12
C41_111 V41 V111 -1.9098932072720259e-19

R41_112 V41 V112 -75477.16586822018
L41_112 V41 V112 5.213225104742305e-12
C41_112 V41 V112 1.7203785661331325e-19

R41_113 V41 V113 -10259.647527165782
L41_113 V41 V113 5.959731986588489e-12
C41_113 V41 V113 1.2330844324883006e-19

R41_114 V41 V114 7716.798998663634
L41_114 V41 V114 5.3475360135977246e-12
C41_114 V41 V114 2.0108929648530737e-19

R41_115 V41 V115 4836.555880486176
L41_115 V41 V115 5.6197957432712136e-12
C41_115 V41 V115 2.185323209524955e-19

R41_116 V41 V116 16929.185575085434
L41_116 V41 V116 -6.75203230405292e-12
C41_116 V41 V116 -5.0497321090750295e-20

R41_117 V41 V117 4861.224676684947
L41_117 V41 V117 -9.228333064241088e-12
C41_117 V41 V117 -8.386996965800338e-20

R41_118 V41 V118 -3562.9375971924237
L41_118 V41 V118 -4.3074749266628e-12
C41_118 V41 V118 -1.739759495777685e-19

R41_119 V41 V119 -3196.9035801976197
L41_119 V41 V119 -4.323098131042938e-12
C41_119 V41 V119 -2.0213037464184896e-19

R41_120 V41 V120 4588.427689039053
L41_120 V41 V120 6.6982698091222e-12
C41_120 V41 V120 -8.996141483875943e-20

R41_121 V41 V121 -6702.702435647665
L41_121 V41 V121 2.857592368310736e-11
C41_121 V41 V121 3.0009502289936276e-20

R41_122 V41 V122 -4532.832123826647
L41_122 V41 V122 5.926816214434682e-12
C41_122 V41 V122 5.857908006368e-20

R41_123 V41 V123 16949.72313035497
L41_123 V41 V123 -4.0559125784260484e-11
C41_123 V41 V123 -5.832468199668378e-20

R41_124 V41 V124 -33159.66712676171
L41_124 V41 V124 -1.1362728403256471e-11
C41_124 V41 V124 -1.0590956072987943e-19

R41_125 V41 V125 2942.32409180698
L41_125 V41 V125 7.598495114013422e-11
C41_125 V41 V125 3.232914965704277e-21

R41_126 V41 V126 4475.28791997728
L41_126 V41 V126 -3.801519140818534e-12
C41_126 V41 V126 8.400816211916411e-21

R41_127 V41 V127 19185.048235484406
L41_127 V41 V127 4.534059235633161e-12
C41_127 V41 V127 -3.097970996408902e-20

R41_128 V41 V128 8533.278360920101
L41_128 V41 V128 1.5249311556400713e-10
C41_128 V41 V128 -5.2154420245381154e-20

R41_129 V41 V129 8256.55570780457
L41_129 V41 V129 2.017901327928579e-11
C41_129 V41 V129 -5.395373575721802e-20

R41_130 V41 V130 27338.31654161387
L41_130 V41 V130 -6.182566859719274e-12
C41_130 V41 V130 -9.917948933607443e-20

R41_131 V41 V131 7378.339104437448
L41_131 V41 V131 -1.6391604550437945e-10
C41_131 V41 V131 5.335453181936808e-20

R41_132 V41 V132 -73057.34096758788
L41_132 V41 V132 -3.650316031065581e-11
C41_132 V41 V132 1.720348810549783e-20

R41_133 V41 V133 -31653.269320908916
L41_133 V41 V133 7.126287492517475e-12
C41_133 V41 V133 1.067813443758376e-19

R41_134 V41 V134 -2839.7308378803905
L41_134 V41 V134 -1.2033268580820203e-11
C41_134 V41 V134 -5.913710093488732e-20

R41_135 V41 V135 -11625.416380021574
L41_135 V41 V135 7.649083985466655e-12
C41_135 V41 V135 -4.5094150165424505e-20

R41_136 V41 V136 15013.756094020546
L41_136 V41 V136 1.1432496300591934e-10
C41_136 V41 V136 -2.0308513467107154e-20

R41_137 V41 V137 3478.0918850806847
L41_137 V41 V137 -4.7313632689572906e-11
C41_137 V41 V137 -1.148653638227658e-19

R41_138 V41 V138 15103.787395248102
L41_138 V41 V138 -4.325416969617007e-12
C41_138 V41 V138 -1.4725887381427716e-19

R41_139 V41 V139 3455.9472368533566
L41_139 V41 V139 3.307714044370077e-12
C41_139 V41 V139 1.2327483978913677e-19

R41_140 V41 V140 -4914.550369941359
L41_140 V41 V140 -1.575959048083575e-11
C41_140 V41 V140 6.978508589871891e-20

R41_141 V41 V141 7485.496174446418
L41_141 V41 V141 -1.39815365600504e-11
C41_141 V41 V141 -4.6654801772223404e-20

R41_142 V41 V142 -4163.813751004959
L41_142 V41 V142 -1.3143048741831743e-11
C41_142 V41 V142 5.1046894310107577e-20

R41_143 V41 V143 -33479.103505950705
L41_143 V41 V143 -7.0792642272521445e-12
C41_143 V41 V143 -2.989251567001868e-20

R41_144 V41 V144 -4296.59991134321
L41_144 V41 V144 9.292345284918476e-12
C41_144 V41 V144 -3.146931847853705e-20

R42_42 V42 0 47.812386984238174
L42_42 V42 0 1.71156850879221e-14
C42_42 V42 0 1.1185320529278961e-17

R42_43 V42 V43 -1461.7002250331268
L42_43 V42 V43 -3.7649101591987785e-13
C42_43 V42 V43 -1.0308543969325767e-18

R42_44 V42 V44 -63904.66300520263
L42_44 V42 V44 7.333670896178598e-12
C42_44 V42 V44 1.175397842273417e-19

R42_45 V42 V45 2351.993686134684
L42_45 V42 V45 1.7728166225344717e-13
C42_45 V42 V45 3.895635427149329e-18

R42_46 V42 V46 -3088.7288402214563
L42_46 V42 V46 6.405474169437698e-13
C42_46 V42 V46 2.2800565640701664e-18

R42_47 V42 V47 1620.5924368222218
L42_47 V42 V47 -1.807147063412666e-11
C42_47 V42 V47 -1.5752856850173381e-19

R42_48 V42 V48 1741.4442493879505
L42_48 V42 V48 7.710021096265638e-13
C42_48 V42 V48 1.0183259395603327e-20

R42_49 V42 V49 -3678.630671734295
L42_49 V42 V49 -9.306663967091601e-13
C42_49 V42 V49 -1.022663171695625e-18

R42_50 V42 V50 -1640.8175136633638
L42_50 V42 V50 -3.276507286714825e-13
C42_50 V42 V50 -8.71813810745859e-19

R42_51 V42 V51 952.5485302257024
L42_51 V42 V51 2.422859154434149e-13
C42_51 V42 V51 1.5436276305183438e-18

R42_52 V42 V52 -909.6522047620828
L42_52 V42 V52 -1.9135856478218526e-13
C42_52 V42 V52 -2.4967496348230295e-18

R42_53 V42 V53 31852.019422162954
L42_53 V42 V53 -5.749379122149012e-13
C42_53 V42 V53 -1.0306207278962095e-18

R42_54 V42 V54 -1487.8145605236298
L42_54 V42 V54 -4.3118352291267405e-13
C42_54 V42 V54 -6.011234832878871e-19

R42_55 V42 V55 -846.1374265199146
L42_55 V42 V55 -3.0516859796753217e-13
C42_55 V42 V55 -7.752797307452578e-19

R42_56 V42 V56 -5685.3146092501165
L42_56 V42 V56 -7.487947353408493e-13
C42_56 V42 V56 -4.372159356486724e-19

R42_57 V42 V57 -170.01828380292045
L42_57 V42 V57 -7.45415214125882e-14
C42_57 V42 V57 4.2582057433374876e-19

R42_58 V42 V58 -269.73512874278373
L42_58 V42 V58 -1.3404098693583972e-13
C42_58 V42 V58 3.741873384278801e-19

R42_59 V42 V59 2188.0160645894134
L42_59 V42 V59 5.334261304983421e-11
C42_59 V42 V59 4.074615901333624e-19

R42_60 V42 V60 -1947.8890141062168
L42_60 V42 V60 -6.114402444337584e-13
C42_60 V42 V60 1.5637277884520971e-19

R42_61 V42 V61 906.1153719878703
L42_61 V42 V61 8.831929449251876e-13
C42_61 V42 V61 -1.5078074847525031e-18

R42_62 V42 V62 831.5919360349844
L42_62 V42 V62 1.0090282163958817e-12
C42_62 V42 V62 -1.5560602366387405e-18

R42_63 V42 V63 -4009.1149959695563
L42_63 V42 V63 -9.081858476024374e-13
C42_63 V42 V63 7.03370141483133e-21

R42_64 V42 V64 6130.457881863278
L42_64 V42 V64 -3.21790055842335e-11
C42_64 V42 V64 5.0848043764692154e-20

R42_65 V42 V65 -391.42677612465184
L42_65 V42 V65 -1.603137566142631e-13
C42_65 V42 V65 -5.384837634505755e-19

R42_66 V42 V66 -390.61952438032336
L42_66 V42 V66 -1.7470734491625726e-13
C42_66 V42 V66 -3.5449676356227403e-19

R42_67 V42 V67 14022.68280725037
L42_67 V42 V67 6.643471893038891e-12
C42_67 V42 V67 -1.3516272129548385e-19

R42_68 V42 V68 -3792.8414971268935
L42_68 V42 V68 -1.1323645273452842e-12
C42_68 V42 V68 -1.488165890595751e-19

R42_69 V42 V69 9393.731577940584
L42_69 V42 V69 8.258571395723408e-13
C42_69 V42 V69 2.2118475263260425e-19

R42_70 V42 V70 1512.3614745051966
L42_70 V42 V70 2.5050888476267933e-12
C42_70 V42 V70 3.591087817220903e-20

R42_71 V42 V71 5365.117747437514
L42_71 V42 V71 1.161359639548342e-11
C42_71 V42 V71 3.7674934986846726e-20

R42_72 V42 V72 1703.7176108566687
L42_72 V42 V72 9.695042974822265e-13
C42_72 V42 V72 2.243987761421788e-20

R42_73 V42 V73 -4138.958506861063
L42_73 V42 V73 -1.6253305886877886e-12
C42_73 V42 V73 -2.1147345275209251e-19

R42_74 V42 V74 4423.346868151771
L42_74 V42 V74 9.017532403779546e-13
C42_74 V42 V74 2.0720918368412778e-19

R42_75 V42 V75 -2206.878442183398
L42_75 V42 V75 -1.0311189346850635e-12
C42_75 V42 V75 -2.9086736313247806e-19

R42_76 V42 V76 -1646.4268083700629
L42_76 V42 V76 -6.889958121096973e-13
C42_76 V42 V76 -1.6029686939720106e-19

R42_77 V42 V77 -3273.6582164810175
L42_77 V42 V77 -1.3442121115700412e-12
C42_77 V42 V77 -1.339670756901836e-19

R42_78 V42 V78 -15668.298050571788
L42_78 V42 V78 -5.889614025627719e-12
C42_78 V42 V78 -1.1137494179077295e-20

R42_79 V42 V79 119725.64211324898
L42_79 V42 V79 5.668196256488056e-12
C42_79 V42 V79 1.3772538202668637e-19

R42_80 V42 V80 11380.226447072399
L42_80 V42 V80 1.5234781969144163e-11
C42_80 V42 V80 -2.1361271593133182e-19

R42_81 V42 V81 8173.4182014319285
L42_81 V42 V81 2.5565897587963594e-12
C42_81 V42 V81 1.309785510209373e-19

R42_82 V42 V82 -21199.675907297813
L42_82 V42 V82 -2.965123023293371e-12
C42_82 V42 V82 -2.1316669184703912e-19

R42_83 V42 V83 -310283.7634510225
L42_83 V42 V83 -2.2688206433715105e-12
C42_83 V42 V83 -2.4229124043878674e-19

R42_84 V42 V84 -10302.88520828004
L42_84 V42 V84 -8.230149999513506e-12
C42_84 V42 V84 8.92740506507054e-20

R42_85 V42 V85 7802.837983242259
L42_85 V42 V85 5.5466285518570796e-12
C42_85 V42 V85 2.1525509090402317e-19

R42_86 V42 V86 215957.3666366634
L42_86 V42 V86 4.23862946314344e-11
C42_86 V42 V86 1.1198914789563944e-19

R42_87 V42 V87 222138.7518657337
L42_87 V42 V87 2.764505950001617e-12
C42_87 V42 V87 1.586906912231691e-19

R42_88 V42 V88 19223.24745197811
L42_88 V42 V88 4.876791177295453e-12
C42_88 V42 V88 2.733945721814806e-22

R42_89 V42 V89 -7276.216701439742
L42_89 V42 V89 -5.132425603249352e-12
C42_89 V42 V89 -1.6173952408013041e-19

R42_90 V42 V90 -110342.81494094095
L42_90 V42 V90 -4.698590670357993e-12
C42_90 V42 V90 -2.0842750948163644e-19

R42_91 V42 V91 1011714.2433027704
L42_91 V42 V91 -2.511918603612735e-12
C42_91 V42 V91 -1.4868250642479304e-19

R42_92 V42 V92 -9820.205130676366
L42_92 V42 V92 -2.1185963899966785e-12
C42_92 V42 V92 -2.0450899435473363e-19

R42_93 V42 V93 3462.4642939981823
L42_93 V42 V93 4.817115265147414e-12
C42_93 V42 V93 3.9991110391807135e-20

R42_94 V42 V94 6471.880635520518
L42_94 V42 V94 3.182208139436475e-12
C42_94 V42 V94 2.951522728974193e-20

R42_95 V42 V95 -18399.70742279077
L42_95 V42 V95 -4.678595436354677e-12
C42_95 V42 V95 -8.952353380433839e-20

R42_96 V42 V96 -9867.359914027853
L42_96 V42 V96 -2.8912010968966084e-12
C42_96 V42 V96 -9.8413668508209e-20

R42_97 V42 V97 6480.148185363045
L42_97 V42 V97 -1.8040955602767904e-11
C42_97 V42 V97 -2.1421610172659126e-20

R42_98 V42 V98 10785.0787579494
L42_98 V42 V98 -1.9544234135348648e-12
C42_98 V42 V98 -2.090142696317407e-19

R42_99 V42 V99 12906.624267562513
L42_99 V42 V99 7.0253808765872e-12
C42_99 V42 V99 3.409135997505959e-20

R42_100 V42 V100 -36562.63532832884
L42_100 V42 V100 6.985729427776589e-12
C42_100 V42 V100 2.3001478152494053e-20

R42_101 V42 V101 23029.705878996603
L42_101 V42 V101 -2.3199216355767754e-12
C42_101 V42 V101 -2.3656447153782425e-19

R42_102 V42 V102 -6327.359673173187
L42_102 V42 V102 -1.3545273185465182e-12
C42_102 V42 V102 -6.27496264264685e-19

R42_103 V42 V103 6554.916910897023
L42_103 V42 V103 3.3265601363829774e-12
C42_103 V42 V103 2.1341113518686111e-19

R42_104 V42 V104 -18285.541135156724
L42_104 V42 V104 -7.421518913074837e-12
C42_104 V42 V104 -2.99445320610473e-20

R42_105 V42 V105 -12838.519020990027
L42_105 V42 V105 1.830917099908335e-12
C42_105 V42 V105 2.826068771934306e-19

R42_106 V42 V106 -3477.896140099144
L42_106 V42 V106 -1.3699826485185198e-12
C42_106 V42 V106 -4.0642034700483157e-19

R42_107 V42 V107 -10405.908033974507
L42_107 V42 V107 -1.7608692479999444e-12
C42_107 V42 V107 -3.9792153726412277e-19

R42_108 V42 V108 7222.167296517753
L42_108 V42 V108 1.600054774866403e-12
C42_108 V42 V108 4.911285413722502e-19

R42_109 V42 V109 10266.159342818604
L42_109 V42 V109 2.491710976842484e-11
C42_109 V42 V109 2.020756929874996e-19

R42_110 V42 V110 18504.16526462546
L42_110 V42 V110 1.7256076028335037e-12
C42_110 V42 V110 3.1567732986013086e-19

R42_111 V42 V111 28879.389763818
L42_111 V42 V111 3.0916595846447163e-12
C42_111 V42 V111 2.064123641636831e-19

R42_112 V42 V112 -4404.614827280308
L42_112 V42 V112 -1.256834858823463e-12
C42_112 V42 V112 -3.815334378075544e-19

R42_113 V42 V113 -6421.691834071572
L42_113 V42 V113 -3.3843978853145565e-12
C42_113 V42 V113 -1.5228199755787437e-19

R42_114 V42 V114 -41437.99659285987
L42_114 V42 V114 -2.532054668736929e-12
C42_114 V42 V114 -1.4800681573572572e-19

R42_115 V42 V115 -14019.575774563398
L42_115 V42 V115 -3.1983965448380632e-12
C42_115 V42 V115 -1.954321470023047e-19

R42_116 V42 V116 6276.217127271738
L42_116 V42 V116 1.9781584546539666e-12
C42_116 V42 V116 3.22566600828722e-19

R42_117 V42 V117 4022.648915553596
L42_117 V42 V117 3.6309294458867e-12
C42_117 V42 V117 2.500898304321644e-19

R42_118 V42 V118 -15256.140744448709
L42_118 V42 V118 2.7271352679328432e-12
C42_118 V42 V118 1.5344976910447388e-19

R42_119 V42 V119 -15952.861016571802
L42_119 V42 V119 2.2797571270674195e-12
C42_119 V42 V119 1.9746611270321236e-19

R42_120 V42 V120 5109.759225804835
L42_120 V42 V120 1.795490112833616e-11
C42_120 V42 V120 4.383569465043651e-20

R42_121 V42 V121 -8682.974953164963
L42_121 V42 V121 -3.2322297140029634e-12
C42_121 V42 V121 -5.408964463678725e-20

R42_122 V42 V122 -7059.812139509173
L42_122 V42 V122 -1.945802525470848e-12
C42_122 V42 V122 3.936767354635216e-20

R42_123 V42 V123 17183.06743492806
L42_123 V42 V123 -2.0512365825428376e-11
C42_123 V42 V123 2.454029118586976e-20

R42_124 V42 V124 -45536.65640665418
L42_124 V42 V124 7.98087689815248e-12
C42_124 V42 V124 -2.0091122222528958e-20

R42_125 V42 V125 4521.552942127839
L42_125 V42 V125 3.2129613228652795e-12
C42_125 V42 V125 8.638934445892361e-20

R42_126 V42 V126 15414.297317175924
L42_126 V42 V126 2.498450987197372e-12
C42_126 V42 V126 -5.940067205136291e-20

R42_127 V42 V127 28074.52162642285
L42_127 V42 V127 -3.2068877969455627e-12
C42_127 V42 V127 -5.428570897308858e-20

R42_128 V42 V128 12672.580297990942
L42_128 V42 V128 -2.296876438125809e-11
C42_128 V42 V128 -2.253084373300748e-20

R42_129 V42 V129 14868.848253135531
L42_129 V42 V129 -2.1885775706116673e-11
C42_129 V42 V129 -1.8559389560232908e-20

R42_130 V42 V130 13676.29582427361
L42_130 V42 V130 4.215752631751985e-12
C42_130 V42 V130 9.356921229175345e-20

R42_131 V42 V131 87405.4578344392
L42_131 V42 V131 -2.5447710621731266e-11
C42_131 V42 V131 -1.2055857698145606e-19

R42_132 V42 V132 10933003.490921997
L42_132 V42 V132 6.734584369567697e-12
C42_132 V42 V132 4.0787823287904536e-20

R42_133 V42 V133 -14973.015687131427
L42_133 V42 V133 -8.755759379248136e-12
C42_133 V42 V133 -1.0564428826640401e-19

R42_134 V42 V134 -4991.1598558399955
L42_134 V42 V134 1.3930926538145483e-11
C42_134 V42 V134 -7.222817540667502e-20

R42_135 V42 V135 55391.124621779614
L42_135 V42 V135 -5.8456588685075096e-12
C42_135 V42 V135 3.1380480208868375e-20

R42_136 V42 V136 24469.25305700685
L42_136 V42 V136 -6.037085538960451e-10
C42_136 V42 V136 -2.2553668485320437e-20

R42_137 V42 V137 5898.956518974596
L42_137 V42 V137 4.012141506482585e-12
C42_137 V42 V137 -2.9572732314295464e-20

R42_138 V42 V138 15108.104771667768
L42_138 V42 V138 2.0755432967305643e-12
C42_138 V42 V138 -5.602329541293371e-20

R42_139 V42 V139 7782.309853277378
L42_139 V42 V139 -2.0740838508296224e-12
C42_139 V42 V139 -1.3326938674921058e-21

R42_140 V42 V140 -8889.192944592634
L42_140 V42 V140 4.28792934336906e-12
C42_140 V42 V140 1.02255481439866e-19

R42_141 V42 V141 13386.855834246893
L42_141 V42 V141 7.037820907298975e-12
C42_141 V42 V141 -1.0462945048421074e-20

R42_142 V42 V142 -8630.544420298653
L42_142 V42 V142 4.255028280312402e-12
C42_142 V42 V142 1.2191123319430478e-19

R42_143 V42 V143 -29865.56009131582
L42_143 V42 V143 8.998674392648843e-12
C42_143 V42 V143 -8.11344966347436e-21

R42_144 V42 V144 -9637.703626518762
L42_144 V42 V144 -6.463336506665466e-12
C42_144 V42 V144 -7.064980799038666e-20

R43_43 V43 0 104.59129971657819
L43_43 V43 0 3.69380716280854e-14
C43_43 V43 0 5.627627785318977e-18

R43_44 V43 V44 19411.251636939352
L43_44 V43 V44 4.2662796671176284e-12
C43_44 V43 V44 5.90218161259857e-20

R43_45 V43 V45 2158.1698318474023
L43_45 V43 V45 3.070381398549739e-13
C43_45 V43 V45 2.1806583809102772e-18

R43_46 V43 V46 -3166.788049999525
L43_46 V43 V46 -1.3094007624459773e-12
C43_46 V43 V46 -2.9193640232608366e-20

R43_47 V43 V47 -1769.1868519273899
L43_47 V43 V47 -1.205347584272044e-12
C43_47 V43 V47 6.17593526515475e-19

R43_48 V43 V48 -253367.4075269333
L43_48 V43 V48 3.2998667192389523e-12
C43_48 V43 V48 1.5005457436828823e-19

R43_49 V43 V49 50902.443702462224
L43_49 V43 V49 -4.723488675087949e-12
C43_49 V43 V49 -5.605996458708375e-19

R43_50 V43 V50 -4711.840016029359
L43_50 V43 V50 -8.551293258633004e-13
C43_50 V43 V50 -1.6906513609471807e-19

R43_51 V43 V51 -121737.6907908612
L43_51 V43 V51 2.3025878328147417e-12
C43_51 V43 V51 2.896353981745732e-21

R43_52 V43 V52 -2958.8528780646716
L43_52 V43 V52 -5.196856883352898e-13
C43_52 V43 V52 -1.092675246338353e-18

R43_53 V43 V53 -2293.796660176585
L43_53 V43 V53 -5.502378772730864e-13
C43_53 V43 V53 -5.525449359102424e-19

R43_54 V43 V54 -4420.981093862938
L43_54 V43 V54 -2.0249627367668044e-12
C43_54 V43 V54 9.926059292736096e-20

R43_55 V43 V55 -2344.296801899205
L43_55 V43 V55 -6.731465434591622e-13
C43_55 V43 V55 -5.202128270552504e-19

R43_56 V43 V56 -2138.7603142901353
L43_56 V43 V56 -7.734005947507004e-13
C43_56 V43 V56 -2.237144100935082e-19

R43_57 V43 V57 -381.9895884324515
L43_57 V43 V57 -1.614676341901721e-13
C43_57 V43 V57 1.911111717128055e-19

R43_58 V43 V58 2861.2545668589296
L43_58 V43 V58 1.0057925321784106e-12
C43_58 V43 V58 1.656433652938122e-19

R43_59 V43 V59 -5708.907807877614
L43_59 V43 V59 -1.4368543258495583e-12
C43_59 V43 V59 2.4230971160074773e-19

R43_60 V43 V60 -2786.2068370666284
L43_60 V43 V60 -1.0920515909742812e-12
C43_60 V43 V60 3.6239875638369493e-20

R43_61 V43 V61 2766.469522884354
L43_61 V43 V61 3.360591321007428e-12
C43_61 V43 V61 -6.567897821730181e-19

R43_62 V43 V62 2556.4004846149205
L43_62 V43 V62 3.4222822891570297e-12
C43_62 V43 V62 -6.614757309081346e-19

R43_63 V43 V63 19289.488686017383
L43_63 V43 V63 8.076374290960537e-12
C43_63 V43 V63 -7.990831539528518e-20

R43_64 V43 V64 -13173.498266637058
L43_64 V43 V64 -4.6262668618425e-12
C43_64 V43 V64 6.24565925238154e-20

R43_65 V43 V65 -928.3638523300955
L43_65 V43 V65 -3.61526363784129e-13
C43_65 V43 V65 -2.173373354128059e-19

R43_66 V43 V66 -1985.4708944199738
L43_66 V43 V66 -5.575400105027954e-13
C43_66 V43 V66 -1.9556619149605603e-19

R43_67 V43 V67 -1145.0201542981647
L43_67 V43 V67 -7.58872448003274e-13
C43_67 V43 V67 -1.9162661506374667e-19

R43_68 V43 V68 -5865.37641680861
L43_68 V43 V68 -4.371227740091444e-12
C43_68 V43 V68 -4.538457319918478e-20

R43_69 V43 V69 -53891.88102914934
L43_69 V43 V69 1.2652426800382165e-12
C43_69 V43 V69 1.4594111843860405e-19

R43_70 V43 V70 4083.2751963490678
L43_70 V43 V70 -1.875124996329796e-11
C43_70 V43 V70 5.390910698457801e-21

R43_71 V43 V71 1908.7405283788707
L43_71 V43 V71 -4.9324051928282856e-11
C43_71 V43 V71 1.0945307660641251e-20

R43_72 V43 V72 -313856.7987256888
L43_72 V43 V72 2.721527495281001e-12
C43_72 V43 V72 6.960681817984008e-21

R43_73 V43 V73 -4333.263851786982
L43_73 V43 V73 -8.181818069637068e-12
C43_73 V43 V73 -7.126190391168196e-20

R43_74 V43 V74 9576.013238448168
L43_74 V43 V74 1.3050324790459302e-12
C43_74 V43 V74 9.936795388655438e-20

R43_75 V43 V75 -3872.2040434426085
L43_75 V43 V75 -1.447400805598708e-12
C43_75 V43 V75 -1.8943966542398103e-19

R43_76 V43 V76 -14500.012976418515
L43_76 V43 V76 -3.778592975034233e-12
C43_76 V43 V76 -4.197344739166951e-20

R43_77 V43 V77 -3547613.27411637
L43_77 V43 V77 -1.0723799253386439e-11
C43_77 V43 V77 -3.167657859107982e-20

R43_78 V43 V78 86292.92983712682
L43_78 V43 V78 -3.328888565407134e-11
C43_78 V43 V78 -7.441255270384925e-21

R43_79 V43 V79 11299.848574959007
L43_79 V43 V79 1.7223204479542104e-12
C43_79 V43 V79 1.8265368524793166e-19

R43_80 V43 V80 -87962.70186765096
L43_80 V43 V80 -3.340232206056379e-12
C43_80 V43 V80 -1.8362731040358439e-19

R43_81 V43 V81 74047.27950384907
L43_81 V43 V81 -1.061608741231731e-11
C43_81 V43 V81 -2.76987743930385e-20

R43_82 V43 V82 -22509.72804917308
L43_82 V43 V82 1.992920202260421e-10
C43_82 V43 V82 -8.928551460693487e-20

R43_83 V43 V83 23794.43076479688
L43_83 V43 V83 -2.9012875390265233e-12
C43_83 V43 V83 -1.7336157893241924e-19

R43_84 V43 V84 -29071.44401983396
L43_84 V43 V84 3.740532812278847e-12
C43_84 V43 V84 1.1740249338251302e-19

R43_85 V43 V85 15247.392509956982
L43_85 V43 V85 3.3725194140751974e-12
C43_85 V43 V85 1.6006255970660976e-19

R43_86 V43 V86 -23209.90940501934
L43_86 V43 V86 9.828074696672071e-12
C43_86 V43 V86 6.922755784914849e-20

R43_87 V43 V87 19408.603518924796
L43_87 V43 V87 5.1127728570048226e-12
C43_87 V43 V87 1.1893681894252478e-19

R43_88 V43 V88 66520.44443225078
L43_88 V43 V88 -2.456509968165096e-11
C43_88 V43 V88 -2.8596093190209844e-20

R43_89 V43 V89 -13352.632332592724
L43_89 V43 V89 -1.2987568478578249e-11
C43_89 V43 V89 -9.712745017829435e-20

R43_90 V43 V90 -26404.069924045965
L43_90 V43 V90 -1.5935906905263857e-12
C43_90 V43 V90 -2.4451580885343877e-19

R43_91 V43 V91 -36605.13627448568
L43_91 V43 V91 -6.206879882611782e-12
C43_91 V43 V91 -1.4457919299763045e-19

R43_92 V43 V92 -27730.58097540405
L43_92 V43 V92 -7.938795503062773e-12
C43_92 V43 V92 -9.358791487425089e-20

R43_93 V43 V93 6170.0294276333425
L43_93 V43 V93 7.341874155648837e-12
C43_93 V43 V93 2.6056940154850517e-20

R43_94 V43 V94 22656.377962498646
L43_94 V43 V94 2.917299172183756e-11
C43_94 V43 V94 1.559247746272075e-20

R43_95 V43 V95 133675.21839968787
L43_95 V43 V95 -1.5620122962811856e-11
C43_95 V43 V95 -6.297881649091512e-20

R43_96 V43 V96 -20993.891821412963
L43_96 V43 V96 -1.811964580772772e-11
C43_96 V43 V96 -4.133503199185685e-20

R43_97 V43 V97 288125.1377815
L43_97 V43 V97 -2.8269406589224084e-12
C43_97 V43 V97 -1.0625919515796944e-19

R43_98 V43 V98 21312.090332969707
L43_98 V43 V98 -3.2402121036757293e-12
C43_98 V43 V98 -1.2006275733270603e-19

R43_99 V43 V99 13464.379440955401
L43_99 V43 V99 5.1510091639520794e-12
C43_99 V43 V99 4.490414490886437e-20

R43_100 V43 V100 -30526.32195385869
L43_100 V43 V100 -1.3372153922067081e-11
C43_100 V43 V100 -4.605748326505961e-20

R43_101 V43 V101 -290576.09879972535
L43_101 V43 V101 -8.489032790825687e-12
C43_101 V43 V101 -1.1371860444448615e-19

R43_102 V43 V102 -9323.016375777905
L43_102 V43 V102 -9.780142636356938e-13
C43_102 V43 V102 -4.633953143825353e-19

R43_103 V43 V103 13036.103748622794
L43_103 V43 V103 1.833279426364542e-12
C43_103 V43 V103 2.4015960657216968e-19

R43_104 V43 V104 -127620.95244586784
L43_104 V43 V104 1.2354074810835848e-10
C43_104 V43 V104 1.6821120449199714e-22

R43_105 V43 V105 36773.85056880619
L43_105 V43 V105 3.1887246056740846e-12
C43_105 V43 V105 1.626610629883194e-19

R43_106 V43 V106 -5273.141180907391
L43_106 V43 V106 -2.3239299007630666e-12
C43_106 V43 V106 -3.066028925554202e-19

R43_107 V43 V107 -8362.412471444635
L43_107 V43 V107 -1.260621727651461e-12
C43_107 V43 V107 -3.8506985758200326e-19

R43_108 V43 V108 5753.655051003822
L43_108 V43 V108 1.6015947739546676e-12
C43_108 V43 V108 3.594703026462002e-19

R43_109 V43 V109 11406.152245362433
L43_109 V43 V109 3.146270999183768e-12
C43_109 V43 V109 1.926240358644528e-19

R43_110 V43 V110 9919.209566498053
L43_110 V43 V110 4.738381783328663e-12
C43_110 V43 V110 2.5913363207134124e-19

R43_111 V43 V111 66600.0711780292
L43_111 V43 V111 2.896006422904196e-12
C43_111 V43 V111 1.329348139340117e-19

R43_112 V43 V112 -9202.323118479675
L43_112 V43 V112 -1.501064832415491e-12
C43_112 V43 V112 -2.30823756147107e-19

R43_113 V43 V113 -14210.669443153942
L43_113 V43 V113 -3.066287102511642e-12
C43_113 V43 V113 -1.2531860360104983e-19

R43_114 V43 V114 -18992.377021563403
L43_114 V43 V114 -5.255259504911291e-12
C43_114 V43 V114 -9.568354244219905e-20

R43_115 V43 V115 320569.2842076984
L43_115 V43 V115 -2.093746258406632e-12
C43_115 V43 V115 -2.043055458472024e-19

R43_116 V43 V116 10468.074222799612
L43_116 V43 V116 1.9912225191356795e-12
C43_116 V43 V116 2.4189572231295163e-19

R43_117 V43 V117 8162.723245740001
L43_117 V43 V117 3.5466344738403885e-12
C43_117 V43 V117 1.959028947381748e-19

R43_118 V43 V118 64636.20316749424
L43_118 V43 V118 3.3916578543262815e-12
C43_118 V43 V118 1.5995466891232899e-19

R43_119 V43 V119 -223848.4825834619
L43_119 V43 V119 3.5888324964794325e-12
C43_119 V43 V119 1.412886114656871e-19

R43_120 V43 V120 13430.195770405795
L43_120 V43 V120 -4.171027395534117e-12
C43_120 V43 V120 4.833586883997557e-20

R43_121 V43 V121 -19237.841033517798
L43_121 V43 V121 -5.224111667963447e-12
C43_121 V43 V121 -2.1062517445152328e-20

R43_122 V43 V122 -24459.34306234073
L43_122 V43 V122 -1.5313354133085262e-12
C43_122 V43 V122 2.1631707141191628e-20

R43_123 V43 V123 162368.0744409186
L43_123 V43 V123 -7.581300171794886e-12
C43_123 V43 V123 1.216538764314562e-20

R43_124 V43 V124 144021.50136698567
L43_124 V43 V124 1.8258224065004572e-11
C43_124 V43 V124 1.7148037598618932e-20

R43_125 V43 V125 8285.573188141576
L43_125 V43 V125 8.020598323413828e-12
C43_125 V43 V125 6.336135785581217e-20

R43_126 V43 V126 35848.8042729767
L43_126 V43 V126 1.3996465563174573e-12
C43_126 V43 V126 -5.4167886865971954e-20

R43_127 V43 V127 54326.16344997309
L43_127 V43 V127 -1.7236445219660171e-12
C43_127 V43 V127 -1.674412264137942e-20

R43_128 V43 V128 29120.573479666105
L43_128 V43 V128 -2.3546556584858338e-11
C43_128 V43 V128 5.084548076098907e-22

R43_129 V43 V129 27218.681831551185
L43_129 V43 V129 -4.480441369397664e-12
C43_129 V43 V129 1.2189472902039946e-21

R43_130 V43 V130 10892.57597867174
L43_130 V43 V130 2.821314806999305e-12
C43_130 V43 V130 9.50649700330179e-20

R43_131 V43 V131 282482.53023573314
L43_131 V43 V131 1.2256914685513081e-11
C43_131 V43 V131 -6.975804859644898e-20

R43_132 V43 V132 -127281.04242927062
L43_132 V43 V132 5.423968912707122e-12
C43_132 V43 V132 1.4096781965534986e-20

R43_133 V43 V133 -20417.178889553106
L43_133 V43 V133 -1.1815077411506953e-10
C43_133 V43 V133 -7.411184082782928e-20

R43_134 V43 V134 -12353.460856905702
L43_134 V43 V134 1.0897100098121089e-11
C43_134 V43 V134 -2.022365595096233e-20

R43_135 V43 V135 -43057.948626255245
L43_135 V43 V135 -3.0200982088326263e-12
C43_135 V43 V135 2.615516281216212e-20

R43_136 V43 V136 51152.1074740807
L43_136 V43 V136 -3.5091427353968397e-10
C43_136 V43 V136 -3.478986021644856e-22

R43_137 V43 V137 9606.11643669409
L43_137 V43 V137 1.5244940424291373e-11
C43_137 V43 V137 -1.126816327178231e-22

R43_138 V43 V138 67656.5165089432
L43_138 V43 V138 1.4405526736529379e-12
C43_138 V43 V138 -2.1962920453730323e-20

R43_139 V43 V139 13543.844366273961
L43_139 V43 V139 -1.3424260283811802e-12
C43_139 V43 V139 9.723683580827882e-22

R43_140 V43 V140 -168335.50813398763
L43_140 V43 V140 3.530831884338491e-12
C43_140 V43 V140 4.031739016317549e-20

R43_141 V43 V141 23930.12441397139
L43_141 V43 V141 6.487665699979647e-12
C43_141 V43 V141 -9.368208898600032e-22

R43_142 V43 V142 -36363.83896628378
L43_142 V43 V142 3.32711470065176e-12
C43_142 V43 V142 2.763111240538977e-20

R43_143 V43 V143 577682.8540722929
L43_143 V43 V143 3.0807907160342066e-12
C43_143 V43 V143 5.602672335598164e-20

R43_144 V43 V144 -8766.165506374578
L43_144 V43 V144 -4.156379968338506e-12
C43_144 V43 V144 -9.439737869804996e-20

R44_44 V44 0 221.5155243002925
L44_44 V44 0 8.633756731360533e-14
C44_44 V44 0 1.9510336642066873e-18

R44_45 V44 V45 9787.860208918826
L44_45 V44 V45 3.750506018639371e-12
C44_45 V44 V45 2.465818817322986e-19

R44_46 V44 V46 4820.699483691091
L44_46 V44 V46 1.8883005091645907e-12
C44_46 V44 V46 1.0328579235546068e-19

R44_47 V44 V47 8822.719984078756
L44_47 V44 V47 2.02586312717267e-12
C44_47 V44 V47 3.0047337945873713e-19

R44_48 V44 V48 -1575.14799079356
L44_48 V44 V48 -1.4467126878792576e-12
C44_48 V44 V48 5.93530638096295e-19

R44_49 V44 V49 -3221.383080194561
L44_49 V44 V49 -2.7219388715101474e-12
C44_49 V44 V49 1.0755096828393208e-19

R44_50 V44 V50 2887.6878953580467
L44_50 V44 V50 8.151834649717855e-12
C44_50 V44 V50 -2.7879579800817285e-19

R44_51 V44 V51 -4112.337202895947
L44_51 V44 V51 -3.1501725220370568e-12
C44_51 V44 V51 -5.429116257208637e-20

R44_52 V44 V52 4567.798387922815
L44_52 V44 V52 -3.468589475705256e-12
C44_52 V44 V52 -3.4899231163986864e-19

R44_53 V44 V53 17366.54225789076
L44_53 V44 V53 2.5659360775951843e-12
C44_53 V44 V53 4.501101134924161e-19

R44_54 V44 V54 22569.818495879463
L44_54 V44 V54 4.677216690742987e-12
C44_54 V44 V54 2.3904475268101664e-19

R44_55 V44 V55 -15941.385578184394
L44_55 V44 V55 1.475554320560685e-11
C44_55 V44 V55 2.1685675940044817e-19

R44_56 V44 V56 6753.627770456132
L44_56 V44 V56 -8.06287138329062e-13
C44_56 V44 V56 -1.025888340486205e-18

R44_57 V44 V57 -6092.441330230169
L44_57 V44 V57 -2.1031877524680945e-12
C44_57 V44 V57 -3.769366021056664e-20

R44_58 V44 V58 5538.340811857355
L44_58 V44 V58 1.4551554196251355e-12
C44_58 V44 V58 1.0147177110461736e-19

R44_59 V44 V59 1466.085472123109
L44_59 V44 V59 7.261681134902023e-13
C44_59 V44 V59 1.5971875114586925e-20

R44_60 V44 V60 -431.94464960686173
L44_60 V44 V60 -2.1893516072013536e-13
C44_60 V44 V60 8.278056322887371e-20

R44_61 V44 V61 9654.554917151936
L44_61 V44 V61 7.396534969541475e-12
C44_61 V44 V61 -9.110966905441324e-21

R44_62 V44 V62 -5835.322350584058
L44_62 V44 V62 -3.1238356979465214e-12
C44_62 V44 V62 -9.153001024693683e-20

R44_63 V44 V63 -8936.748584509549
L44_63 V44 V63 -5.260203403867868e-12
C44_63 V44 V63 -1.461199063723936e-20

R44_64 V44 V64 -11803.895719288746
L44_64 V44 V64 -1.6054817982283958e-12
C44_64 V44 V64 -5.887981764284814e-19

R44_65 V44 V65 101355.01078693708
L44_65 V44 V65 -3.388921661791083e-12
C44_65 V44 V65 -2.1821569246869893e-20

R44_66 V44 V66 10623.898142900105
L44_66 V44 V66 -3.494887516530287e-12
C44_66 V44 V66 -7.099420345535822e-20

R44_67 V44 V67 -8397.568422058323
L44_67 V44 V67 -1.2789725376841447e-11
C44_67 V44 V67 -4.8368372103136104e-20

R44_68 V44 V68 -1134.888900541574
L44_68 V44 V68 -4.3425191625813465e-13
C44_68 V44 V68 -1.375522737227052e-19

R44_69 V44 V69 20900.382886337586
L44_69 V44 V69 2.5971434126454072e-12
C44_69 V44 V69 2.1944911957121428e-20

R44_70 V44 V70 -33189.43939459222
L44_70 V44 V70 9.969993540089497e-12
C44_70 V44 V70 7.942987433224793e-20

R44_71 V44 V71 7970.639617814562
L44_71 V44 V71 3.255622319873711e-10
C44_71 V44 V71 1.6184989824693186e-20

R44_72 V44 V72 -62691.72744028713
L44_72 V44 V72 2.568477993228909e-12
C44_72 V44 V72 1.0270550702158726e-20

R44_73 V44 V73 -3526.73710330618
L44_73 V44 V73 -2.470676861127664e-12
C44_73 V44 V73 9.6453386932548e-21

R44_74 V44 V74 -12906.31029018969
L44_74 V44 V74 1.7248927774500148e-11
C44_74 V44 V74 3.006511581747698e-20

R44_75 V44 V75 31062.585883478725
L44_75 V44 V75 -1.1544730978970641e-11
C44_75 V44 V75 -8.229009973884107e-20

R44_76 V44 V76 18273.323425911218
L44_76 V44 V76 -4.383130101904746e-11
C44_76 V44 V76 2.0665710072140733e-20

R44_77 V44 V77 8816.497841267033
L44_77 V44 V77 3.356433721787042e-12
C44_77 V44 V77 3.7198062292159216e-20

R44_78 V44 V78 24870.87200837508
L44_78 V44 V78 9.921763309260363e-12
C44_78 V44 V78 5.590158577322023e-20

R44_79 V44 V79 -250226.7276013521
L44_79 V44 V79 5.1437207945279235e-12
C44_79 V44 V79 1.10538060251236e-19

R44_80 V44 V80 -18144.104307393318
L44_80 V44 V80 -6.641008064104702e-12
C44_80 V44 V80 -1.9462787007906986e-19

R44_81 V44 V81 -55116.330028371616
L44_81 V44 V81 -1.305184876361018e-11
C44_81 V44 V81 1.1372207686052307e-19

R44_82 V44 V82 -23870.858300387234
L44_82 V44 V82 -4.650875663822285e-12
C44_82 V44 V82 -1.0575541016709208e-19

R44_83 V44 V83 -53469.914860712444
L44_83 V44 V83 -5.214977866877439e-12
C44_83 V44 V83 -1.5525200458743228e-19

R44_84 V44 V84 161771.58437992286
L44_84 V44 V84 6.2295817412580136e-12
C44_84 V44 V84 6.136268176104269e-20

R44_85 V44 V85 -45085.78489192709
L44_85 V44 V85 6.204483518681681e-12
C44_85 V44 V85 8.878990436839955e-20

R44_86 V44 V86 -9185.150499643198
L44_86 V44 V86 1.5737576003021777e-11
C44_86 V44 V86 -3.2156851534772926e-20

R44_87 V44 V87 22184.783082900067
L44_87 V44 V87 5.468629488167084e-12
C44_87 V44 V87 1.1761242799459633e-19

R44_88 V44 V88 19617.56517218194
L44_88 V44 V88 4.597479899227456e-11
C44_88 V44 V88 5.511149903073951e-20

R44_89 V44 V89 -105588.21733293822
L44_89 V44 V89 -7.818968311375713e-12
C44_89 V44 V89 -8.829249052543747e-20

R44_90 V44 V90 -22516.967513182906
L44_90 V44 V90 -4.3081410720992485e-12
C44_90 V44 V90 -1.292507551835077e-19

R44_91 V44 V91 -108143.81725718273
L44_91 V44 V91 -4.675108553064989e-12
C44_91 V44 V91 -4.6033069031240114e-20

R44_92 V44 V92 -10693.803276173267
L44_92 V44 V92 -8.326225204247756e-12
C44_92 V44 V92 -2.3489531365675303e-19

R44_93 V44 V93 90428.05374296362
L44_93 V44 V93 1.7867516526383494e-11
C44_93 V44 V93 1.1531496224738145e-20

R44_94 V44 V94 26583.053426329367
L44_94 V44 V94 1.4355685527153948e-11
C44_94 V44 V94 8.701418578326309e-20

R44_95 V44 V95 339459.017494736
L44_95 V44 V95 -9.864228408612907e-12
C44_95 V44 V95 -4.8938322137614514e-20

R44_96 V44 V96 -90158.1150401418
L44_96 V44 V96 -2.98515082555285e-11
C44_96 V44 V96 -1.924913704525738e-19

R44_97 V44 V97 -52898.21752931703
L44_97 V44 V97 -1.0745399782222511e-11
C44_97 V44 V97 8.678389985664455e-21

R44_98 V44 V98 -21785.543362069464
L44_98 V44 V98 -4.939297829426422e-12
C44_98 V44 V98 -1.020703034981938e-19

R44_99 V44 V99 54287.091251537364
L44_99 V44 V99 1.2633999326846027e-11
C44_99 V44 V99 4.6330428014188256e-20

R44_100 V44 V100 11258.536073660034
L44_100 V44 V100 -3.67327122972078e-09
C44_100 V44 V100 1.2385487966410688e-19

R44_101 V44 V101 -22259.8864468283
L44_101 V44 V101 -6.528191760262885e-12
C44_101 V44 V101 -1.241184787210878e-19

R44_102 V44 V102 -12497.091669634188
L44_102 V44 V102 -2.2635765246970753e-12
C44_102 V44 V102 -2.0907269274923767e-19

R44_103 V44 V103 49690.9963518335
L44_103 V44 V103 5.5550706292566884e-12
C44_103 V44 V103 1.3224978210936643e-19

R44_104 V44 V104 -12494.054805040287
L44_104 V44 V104 5.850142621087368e-11
C44_104 V44 V104 -1.7932591783354797e-19

R44_105 V44 V105 7774.9872272695475
L44_105 V44 V105 4.76609488208775e-12
C44_105 V44 V105 1.9281553707812312e-19

R44_106 V44 V106 -13949.491327104817
L44_106 V44 V106 -3.169721125728528e-12
C44_106 V44 V106 -2.4515077646508277e-19

R44_107 V44 V107 -16924.865909141587
L44_107 V44 V107 -3.001485010334773e-12
C44_107 V44 V107 -1.8797712819889203e-19

R44_108 V44 V108 6344.450695508334
L44_108 V44 V108 3.3709775876168187e-12
C44_108 V44 V108 2.9320294156669325e-19

R44_109 V44 V109 -8019.129180893989
L44_109 V44 V109 8.208349654109815e-12
C44_109 V44 V109 -1.3535694069820162e-19

R44_110 V44 V110 23303.373468351
L44_110 V44 V110 4.439513727597788e-12
C44_110 V44 V110 1.7105297041856688e-19

R44_111 V44 V111 31176.984894943194
L44_111 V44 V111 6.285957282971166e-12
C44_111 V44 V111 1.2208888515626604e-19

R44_112 V44 V112 -9627.815307486368
L44_112 V44 V112 -2.95223790097297e-12
C44_112 V44 V112 -1.8872107735131246e-19

R44_113 V44 V113 14405.331524235537
L44_113 V44 V113 -5.648270993151774e-12
C44_113 V44 V113 3.9480318072498616e-20

R44_114 V44 V114 -79314.5652683174
L44_114 V44 V114 -6.938212413701836e-12
C44_114 V44 V114 -9.796613103983916e-20

R44_115 V44 V115 -21043.622915930668
L44_115 V44 V115 -5.204061751126508e-12
C44_115 V44 V115 -1.3731163488287823e-19

R44_116 V44 V116 11836.294581522508
L44_116 V44 V116 4.5639285163686e-12
C44_116 V44 V116 1.609271350313609e-19

R44_117 V44 V117 -94421.88632858044
L44_117 V44 V117 7.045857616476053e-12
C44_117 V44 V117 3.148793126791381e-20

R44_118 V44 V118 -140208.72009107776
L44_118 V44 V118 5.426154025080677e-12
C44_118 V44 V118 2.746800418443298e-20

R44_119 V44 V119 16970.269164875757
L44_119 V44 V119 5.35169665355098e-12
C44_119 V44 V119 1.7243339132164867e-19

R44_120 V44 V120 17607.029959757965
L44_120 V44 V120 -2.244555062983596e-11
C44_120 V44 V120 1.1718414978182035e-19

R44_121 V44 V121 -17030.255423665432
L44_121 V44 V121 -8.692593261105939e-12
C44_121 V44 V121 -2.5411551218099563e-20

R44_122 V44 V122 -25961.8270872046
L44_122 V44 V122 -3.5736422653706534e-12
C44_122 V44 V122 -1.2764331034013806e-20

R44_123 V44 V123 -111385.68109297438
L44_123 V44 V123 -4.051289889185055e-11
C44_123 V44 V123 1.2436658322905758e-20

R44_124 V44 V124 17873.327741185996
L44_124 V44 V124 1.5769827521953633e-11
C44_124 V44 V124 1.224689998327684e-19

R44_125 V44 V125 40122.26953111863
L44_125 V44 V125 1.11150198606653e-11
C44_125 V44 V125 -2.227375802075602e-21

R44_126 V44 V126 31709.42873287272
L44_126 V44 V126 3.69963355578174e-12
C44_126 V44 V126 -9.835957736631987e-21

R44_127 V44 V127 120781.15173936405
L44_127 V44 V127 -4.6291619122229106e-12
C44_127 V44 V127 3.99705592418004e-20

R44_128 V44 V128 2906537.4605114837
L44_128 V44 V128 -8.974890205990952e-11
C44_128 V44 V128 4.238234538540724e-21

R44_129 V44 V129 159699.09809199383
L44_129 V44 V129 -1.8191840497249854e-11
C44_129 V44 V129 4.1983704555369576e-20

R44_130 V44 V130 74292.09703609663
L44_130 V44 V130 6.7487315860030714e-12
C44_130 V44 V130 4.4621537678948345e-20

R44_131 V44 V131 -37742.073619741896
L44_131 V44 V131 6.915281089991059e-11
C44_131 V44 V131 -6.262520041565818e-20

R44_132 V44 V132 -1836041.0993428535
L44_132 V44 V132 1.5454406638411285e-11
C44_132 V44 V132 1.2464231045357781e-20

R44_133 V44 V133 430123.4540905294
L44_133 V44 V133 -1.5373763697063915e-11
C44_133 V44 V133 -5.0568122764580905e-20

R44_134 V44 V134 -88950.94740045538
L44_134 V44 V134 2.1010776841698717e-11
C44_134 V44 V134 -1.7248135744627136e-20

R44_135 V44 V135 63272.59083054629
L44_135 V44 V135 -8.34083351412354e-12
C44_135 V44 V135 4.3885295670021953e-20

R44_136 V44 V136 78553.97369812027
L44_136 V44 V136 1.4349691466152923e-10
C44_136 V44 V136 1.8341390354391033e-20

R44_137 V44 V137 16098.853745198476
L44_137 V44 V137 1.1058096700889484e-11
C44_137 V44 V137 8.857803459480492e-20

R44_138 V44 V138 18284.117920371653
L44_138 V44 V138 3.64992630720907e-12
C44_138 V44 V138 7.626027652520818e-20

R44_139 V44 V139 -42689.84984229875
L44_139 V44 V139 -3.338075296484179e-12
C44_139 V44 V139 -2.9872895516170517e-20

R44_140 V44 V140 38056.9685863191
L44_140 V44 V140 7.903351570783568e-12
C44_140 V44 V140 -2.0109670663157347e-21

R44_141 V44 V141 -81348.70367891248
L44_141 V44 V141 1.8320714174664818e-11
C44_141 V44 V141 -3.6609703641602344e-21

R44_142 V44 V142 10993.589941669152
L44_142 V44 V142 7.9897720795759e-12
C44_142 V44 V142 6.24688742031646e-20

R44_143 V44 V143 36247.876590399035
L44_143 V44 V143 9.353022783014625e-12
C44_143 V44 V143 4.0457619811987625e-20

R44_144 V44 V144 29316.60964948937
L44_144 V44 V144 -1.0170125068176483e-11
C44_144 V44 V144 1.8874420805962083e-20

R45_45 V45 0 88.44956372226778
L45_45 V45 0 -2.5928195029726207e-14
C45_45 V45 0 -1.3418993254047006e-17

R45_46 V45 V46 -666.5757142157087
L45_46 V45 V46 3.218458073493163e-13
C45_46 V45 V46 -4.793954084127268e-19

R45_47 V45 V47 -1992.1134693977979
L45_47 V45 V47 4.2695031514909447e-13
C45_47 V45 V47 -9.066856002739071e-20

R45_48 V45 V48 87890.9249816804
L45_48 V45 V48 -1.8331522846314954e-12
C45_48 V45 V48 -1.0580077146562461e-19

R45_49 V45 V49 1848.4858514584769
L45_49 V45 V49 4.080955592426741e-12
C45_49 V45 V49 1.4737266513232615e-18

R45_50 V45 V50 2011.1298786262619
L45_50 V45 V50 4.900082033016579e-13
C45_50 V45 V50 3.1614932428384233e-19

R45_51 V45 V51 5009.722559200599
L45_51 V45 V51 -5.873471522137242e-13
C45_51 V45 V51 -9.457902555914882e-19

R45_52 V45 V52 623.4838319376595
L45_52 V45 V52 3.3380293240796504e-13
C45_52 V45 V52 2.571696450493292e-18

R45_53 V45 V53 1509.9695798209962
L45_53 V45 V53 8.085983265025631e-13
C45_53 V45 V53 9.4870040867081e-19

R45_54 V45 V54 -1655.707227317204
L45_54 V45 V54 9.208600885335048e-13
C45_54 V45 V54 2.5705083254776703e-19

R45_55 V45 V55 -1179.3662912593447
L45_55 V45 V55 4.750515414672639e-13
C45_55 V45 V55 1.216122013895094e-18

R45_56 V45 V56 -3876.3505280262516
L45_56 V45 V56 5.648461851695908e-13
C45_56 V45 V56 1.1059652705925858e-18

R45_57 V45 V57 -120.64472549264408
L45_57 V45 V57 1.4070609888885598e-13
C45_57 V45 V57 -3.6799014170605145e-19

R45_58 V45 V58 -468.01599340915044
L45_58 V45 V58 5.887642365154734e-13
C45_58 V45 V58 -2.8508665507692666e-19

R45_59 V45 V59 1187.1712911709026
L45_59 V45 V59 3.555557682969705e-13
C45_59 V45 V59 -3.9621178146189142e-19

R45_60 V45 V60 -1915.1279352138934
L45_60 V45 V60 3.518219424253885e-13
C45_60 V45 V60 -1.236441036003232e-19

R45_61 V45 V61 346.3017271779423
L45_61 V45 V61 -1.15935123967254e-12
C45_61 V45 V61 1.455039172290973e-18

R45_62 V45 V62 277.4846109407784
L45_62 V45 V62 1.4741420300246888e-12
C45_62 V45 V62 1.3797270191917378e-18

R45_63 V45 V63 3302.5469874696146
L45_63 V45 V63 2.1418103127630256e-12
C45_63 V45 V63 3.4214942827327507e-19

R45_64 V45 V64 6257.19982923443
L45_64 V45 V64 1.5335431104752235e-12
C45_64 V45 V64 2.974969387576229e-19

R45_65 V45 V65 -382.376957804489
L45_65 V45 V65 2.933398914926946e-13
C45_65 V45 V65 4.1452581306235826e-19

R45_66 V45 V66 -389.67536750421453
L45_66 V45 V66 3.5918079414344403e-13
C45_66 V45 V66 4.548364779230632e-19

R45_67 V45 V67 -5998.909390435958
L45_67 V45 V67 8.258813928640818e-13
C45_67 V45 V67 3.8014523067422527e-19

R45_68 V45 V68 -12670.358852358613
L45_68 V45 V68 1.1882534859301618e-12
C45_68 V45 V68 2.2238455684831948e-19

R45_69 V45 V69 -3568.9409555366483
L45_69 V45 V69 -4.691378456332873e-13
C45_69 V45 V69 -2.9888654134346852e-19

R45_70 V45 V70 1322.5782679224722
L45_70 V45 V70 3.0781451349833197e-12
C45_70 V45 V70 9.023134714041277e-20

R45_71 V45 V71 -6813.23194633584
L45_71 V45 V71 -5.570782532709476e-12
C45_71 V45 V71 3.5919739712935325e-20

R45_72 V45 V72 1249.3240182984782
L45_72 V45 V72 -2.0329806869449013e-12
C45_72 V45 V72 1.9619297474235822e-20

R45_73 V45 V73 6667.763116392364
L45_73 V45 V73 2.3404670809803207e-12
C45_73 V45 V73 2.1576189893941657e-19

R45_74 V45 V74 4622.67407585531
L45_74 V45 V74 -1.1511447565462658e-12
C45_74 V45 V74 -1.742376888917954e-19

R45_75 V45 V75 -2249.8694394661366
L45_75 V45 V75 1.9213433803558425e-12
C45_75 V45 V75 3.0847053678913406e-19

R45_76 V45 V76 -3384.401263241196
L45_76 V45 V76 1.466439185548649e-12
C45_76 V45 V76 1.8239076375497758e-19

R45_77 V45 V77 -8020.35716731651
L45_77 V45 V77 5.247296392362691e-12
C45_77 V45 V77 4.5483651114761994e-20

R45_78 V45 V78 8119.9837699850295
L45_78 V45 V78 4.116543494342469e-12
C45_78 V45 V78 -2.572920174459658e-20

R45_79 V45 V79 8492.562567138331
L45_79 V45 V79 -7.0778808065130644e-12
C45_79 V45 V79 -3.642438155777885e-20

R45_80 V45 V80 6713.066793874306
L45_80 V45 V80 -1.6180443860952358e-11
C45_80 V45 V80 9.402651647066888e-20

R45_81 V45 V81 63003.996075380295
L45_81 V45 V81 -6.450860592996811e-11
C45_81 V45 V81 -4.6260856611731124e-20

R45_82 V45 V82 5074.385507749035
L45_82 V45 V82 2.0458935013343977e-12
C45_82 V45 V82 3.95694719271046e-19

R45_83 V45 V83 31148.20050391531
L45_83 V45 V83 2.221194457289018e-12
C45_83 V45 V83 4.2173238913976076e-19

R45_84 V45 V84 -22414.623192819916
L45_84 V45 V84 1.0832348028616193e-11
C45_84 V45 V84 3.5994517326416217e-20

R45_85 V45 V85 11293.421439132038
L45_85 V45 V85 -9.16485620117939e-12
C45_85 V45 V85 -1.0760117770867889e-19

R45_86 V45 V86 34329.20775868423
L45_86 V45 V86 -6.951701278178057e-12
C45_86 V45 V86 -1.537873439881134e-19

R45_87 V45 V87 -6975.058787364953
L45_87 V45 V87 -3.803607467246263e-12
C45_87 V45 V87 -2.0005387487027517e-19

R45_88 V45 V88 25636.760546259426
L45_88 V45 V88 -1.2621615167206258e-11
C45_88 V45 V88 -4.6189790425520543e-20

R45_89 V45 V89 -102744.96073619416
L45_89 V45 V89 7.878743016944726e-12
C45_89 V45 V89 1.2337601645366585e-19

R45_90 V45 V90 42495.053506863
L45_90 V45 V90 7.375261550471195e-12
C45_90 V45 V90 8.105033036672101e-20

R45_91 V45 V91 5301.63512088274
L45_91 V45 V91 1.6519824882889657e-12
C45_91 V45 V91 4.47583911300063e-19

R45_92 V45 V92 21493.6339116128
L45_92 V45 V92 3.8684007936532585e-12
C45_92 V45 V92 2.3829045457352396e-19

R45_93 V45 V93 2258.6289138075886
L45_93 V45 V93 -8.281021441373769e-12
C45_93 V45 V93 -5.945014535254816e-20

R45_94 V45 V94 8299.500179601531
L45_94 V45 V94 -4.644438301386502e-12
C45_94 V45 V94 -1.5557461243392452e-19

R45_95 V45 V95 17563.320733515568
L45_95 V45 V95 3.4228678073104085e-12
C45_95 V45 V95 2.1342557557107615e-19

R45_96 V45 V96 -16807.89647745897
L45_96 V45 V96 1.5914911900241674e-11
C45_96 V45 V96 1.0221428058926696e-19

R45_97 V45 V97 4848.8200669937105
L45_97 V45 V97 -1.569174690037336e-11
C45_97 V45 V97 -8.750890784947789e-20

R45_98 V45 V98 3451.289371969474
L45_98 V45 V98 3.468219595787165e-12
C45_98 V45 V98 2.188423364310042e-19

R45_99 V45 V99 11192.781945658397
L45_99 V45 V99 -1.3556784203739554e-11
C45_99 V45 V99 -4.9469635255516004e-20

R45_100 V45 V100 -16662.5205074794
L45_100 V45 V100 -2.2912135082802272e-11
C45_100 V45 V100 -4.080679910233618e-20

R45_101 V45 V101 3579.407507911137
L45_101 V45 V101 4.677755361691859e-12
C45_101 V45 V101 2.107420185774541e-19

R45_102 V45 V102 4602.300221152566
L45_102 V45 V102 2.2070131053053855e-12
C45_102 V45 V102 3.2774250916590597e-19

R45_103 V45 V103 9478.790568304212
L45_103 V45 V103 -1.4040890561005245e-11
C45_103 V45 V103 -2.127110277053935e-20

R45_104 V45 V104 -22801.157281997635
L45_104 V45 V104 -1.3033606420952849e-11
C45_104 V45 V104 -3.434544116769459e-20

R45_105 V45 V105 -3116.0329374843295
L45_105 V45 V105 -2.4698288610658243e-12
C45_105 V45 V105 -3.3998369751284525e-19

R45_106 V45 V106 -163872.22416710365
L45_106 V45 V106 1.5602846266293492e-12
C45_106 V45 V106 5.217768614277037e-19

R45_107 V45 V107 6846.835111104121
L45_107 V45 V107 2.8803230622373412e-12
C45_107 V45 V107 2.5733877592554587e-19

R45_108 V45 V108 -5671.834365653518
L45_108 V45 V108 -3.6736187380874e-12
C45_108 V45 V108 -2.783304212135235e-19

R45_109 V45 V109 -28654.030106587987
L45_109 V45 V109 -6.986482423517462e-12
C45_109 V45 V109 -1.1266471300403953e-19

R45_110 V45 V110 -4206.9537310949545
L45_110 V45 V110 -1.8310085158161907e-12
C45_110 V45 V110 -4.92083100239449e-19

R45_111 V45 V111 -7499.038317399949
L45_111 V45 V111 -4.417254246355857e-12
C45_111 V45 V111 -1.5962903417998527e-19

R45_112 V45 V112 -22739.48634127844
L45_112 V45 V112 2.70614085593349e-12
C45_112 V45 V112 2.2639703116837375e-19

R45_113 V45 V113 -10017.307185014926
L45_113 V45 V113 4.400795633856655e-12
C45_113 V45 V113 1.1587131446700501e-19

R45_114 V45 V114 6634.227698165426
L45_114 V45 V114 3.372327315585018e-12
C45_114 V45 V114 2.532608406276814e-19

R45_115 V45 V115 11457.90116952748
L45_115 V45 V115 5.061633088834013e-12
C45_115 V45 V115 9.321018256544679e-20

R45_116 V45 V116 -87384.76694808256
L45_116 V45 V116 -4.304803286817498e-12
C45_116 V45 V116 -1.7784085348227189e-19

R45_117 V45 V117 7480.560896151716
L45_117 V45 V117 -5.153043838366933e-12
C45_117 V45 V117 -1.4289532769885034e-19

R45_118 V45 V118 -4013.6048466453867
L45_118 V45 V118 -2.9582671879073877e-12
C45_118 V45 V118 -2.530836267617288e-19

R45_119 V45 V119 -3166.290750735177
L45_119 V45 V119 -2.6802551847735252e-12
C45_119 V45 V119 -2.9532134627102984e-19

R45_120 V45 V120 4467.410630735627
L45_120 V45 V120 4.230108876144003e-11
C45_120 V45 V120 -4.736614113810552e-20

R45_121 V45 V121 -5262.274886051405
L45_121 V45 V121 6.258904037657242e-12
C45_121 V45 V121 7.22120280907224e-20

R45_122 V45 V122 -3265.4075666385475
L45_122 V45 V122 5.160401686117127e-12
C45_122 V45 V122 -4.542633240133042e-20

R45_123 V45 V123 19406.751499889484
L45_123 V45 V123 -1.049940302752202e-11
C45_123 V45 V123 -6.923263644399339e-20

R45_124 V45 V124 -68199.93825958602
L45_124 V45 V124 -8.554022832527334e-12
C45_124 V45 V124 -4.7627485832729256e-20

R45_125 V45 V125 3078.432493999154
L45_125 V45 V125 -1.2789905756022817e-11
C45_125 V45 V125 -6.327219370229238e-20

R45_126 V45 V126 4394.366477733735
L45_126 V45 V126 -5.358476057629323e-12
C45_126 V45 V126 5.903548325878146e-20

R45_127 V45 V127 26537.0292456593
L45_127 V45 V127 5.569625964729813e-12
C45_127 V45 V127 1.4143125149159962e-20

R45_128 V45 V128 9954.988370125622
L45_128 V45 V128 -2.482383453402751e-10
C45_128 V45 V128 -9.714188583277769e-21

R45_129 V45 V129 9474.220730586663
L45_129 V45 V129 -7.985423613299462e-11
C45_129 V45 V129 -1.75012701241266e-20

R45_130 V45 V130 -215246.4350454083
L45_130 V45 V130 -9.399922413419666e-12
C45_130 V45 V130 -7.134285687410018e-20

R45_131 V45 V131 10009.515347564235
L45_131 V45 V131 2.030007406674658e-11
C45_131 V45 V131 6.567816554183505e-20

R45_132 V45 V132 -732773.0403936993
L45_132 V45 V132 -2.3813474434492335e-11
C45_132 V45 V132 -3.9771812125050416e-21

R45_133 V45 V133 25378.107986134753
L45_133 V45 V133 4.890961380131156e-12
C45_133 V45 V133 1.792458024472954e-19

R45_134 V45 V134 -4624.113133197513
L45_134 V45 V134 -8.413524796058062e-11
C45_134 V45 V134 1.6768795177618972e-20

R45_135 V45 V135 -20879.58513315043
L45_135 V45 V135 1.1360660238016316e-11
C45_135 V45 V135 -1.1409860427768017e-20

R45_136 V45 V136 16109.034695067528
L45_136 V45 V136 4.777493202826904e-11
C45_136 V45 V136 6.406619161202838e-21

R45_137 V45 V137 3508.2095475639394
L45_137 V45 V137 -8.420722366685262e-12
C45_137 V45 V137 -4.123277564588659e-20

R45_138 V45 V138 5971.3565274602515
L45_138 V45 V138 -4.58738330508238e-12
C45_138 V45 V138 4.032880056103956e-20

R45_139 V45 V139 7000.079697111921
L45_139 V45 V139 4.132879750690874e-12
C45_139 V45 V139 -1.8586910143762567e-20

R45_140 V45 V140 -5045.983510364862
L45_140 V45 V140 -1.1245741791447217e-11
C45_140 V45 V140 -6.768009827067688e-20

R45_141 V45 V141 7300.1806249819765
L45_141 V45 V141 -1.399486993228018e-11
C45_141 V45 V141 3.44051869120625e-21

R45_142 V45 V142 -3994.749904242611
L45_142 V45 V142 -5.5955410370717535e-12
C45_142 V45 V142 -1.0778736007346173e-19

R45_143 V45 V143 -25643.965239147663
L45_143 V45 V143 -1.3990329634246296e-11
C45_143 V45 V143 -5.111490798086521e-21

R45_144 V45 V144 -8205.006089995775
L45_144 V45 V144 1.0578359586533157e-11
C45_144 V45 V144 9.127844376188982e-20

R46_46 V46 0 53.68863392472322
L46_46 V46 0 9.012648958080489e-12
C46_46 V46 0 -4.239582939171132e-18

R46_47 V46 V47 -2183.7329652502835
L46_47 V46 V47 -5.130159258347011e-13
C46_47 V46 V47 -3.1404824768166117e-19

R46_48 V46 V48 1278.818393669409
L46_48 V46 V48 4.264538447837492e-11
C46_48 V46 V48 -8.001318166207294e-20

R46_49 V46 V49 969.3309533162278
L46_49 V46 V49 2.4282857047854655e-12
C46_49 V46 V49 -6.567131720617283e-20

R46_50 V46 V50 -1555.6435540911436
L46_50 V46 V50 -2.651291408886586e-12
C46_50 V46 V50 8.380006630772637e-19

R46_51 V46 V51 5462.610086003539
L46_51 V46 V51 -1.2210935068872412e-11
C46_51 V46 V51 -4.923659140188194e-19

R46_52 V46 V52 1791.6703275014868
L46_52 V46 V52 9.89624050218225e-11
C46_52 V46 V52 9.74215619782428e-19

R46_53 V46 V53 1839.3068785197008
L46_53 V46 V53 7.751271264365236e-12
C46_53 V46 V53 6.353857326252116e-19

R46_54 V46 V54 -1970.7968311445604
L46_54 V46 V54 2.438706819716106e-10
C46_54 V46 V54 2.0835339273163541e-19

R46_55 V46 V55 -1585.6390678972539
L46_55 V46 V55 -3.073613563524476e-12
C46_55 V46 V55 -2.724992311575676e-19

R46_56 V46 V56 -4177.167906731161
L46_56 V46 V56 -1.864979613387886e-12
C46_56 V46 V56 -1.1686739975520383e-19

R46_57 V46 V57 -127.32922719871638
L46_57 V46 V57 1.2600787607496108e-12
C46_57 V46 V57 -1.860323319533004e-19

R46_58 V46 V58 -268.51034579313466
L46_58 V46 V58 9.623059744986658e-13
C46_58 V46 V58 -1.2897790774315752e-19

R46_59 V46 V59 -797.7514125278714
L46_59 V46 V59 -3.8525590420652535e-13
C46_59 V46 V59 -7.036903933106633e-20

R46_60 V46 V60 -1015.6887809418174
L46_60 V46 V60 -9.35188974415767e-13
C46_60 V46 V60 -8.202621302372946e-20

R46_61 V46 V61 356.87496163347674
L46_61 V46 V61 3.1661395803201715e-12
C46_61 V46 V61 6.983675007332022e-19

R46_62 V46 V62 422.6832285141205
L46_62 V46 V62 -9.188190650639723e-13
C46_62 V46 V62 6.075008451517292e-19

R46_63 V46 V63 -4278.970836801852
L46_63 V46 V63 -4.5105923786278204e-11
C46_63 V46 V63 1.8505970463690616e-20

R46_64 V46 V64 -9581.233646866092
L46_64 V46 V64 -3.54456523039568e-12
C46_64 V46 V64 -1.6003670223025386e-20

R46_65 V46 V65 -350.6757954796324
L46_65 V46 V65 2.0166687893085515e-12
C46_65 V46 V65 3.739078589285411e-19

R46_66 V46 V66 -359.6172950242289
L46_66 V46 V66 1.9328763427337988e-12
C46_66 V46 V66 -8.596746111105893e-20

R46_67 V46 V67 -3861.0165033041026
L46_67 V46 V67 -1.3805695019025818e-12
C46_67 V46 V67 -1.309718697382661e-19

R46_68 V46 V68 -13150.293262438381
L46_68 V46 V68 8.502643715915287e-11
C46_68 V46 V68 6.292424838386694e-20

R46_69 V46 V69 1977.2816241679157
L46_69 V46 V69 7.740966099995122e-13
C46_69 V46 V69 9.698445258913258e-20

R46_70 V46 V70 1759.372531947505
L46_70 V46 V70 -1.6691132803068346e-12
C46_70 V46 V70 2.9125067301609813e-20

R46_71 V46 V71 7045.7869095763235
L46_71 V46 V71 -2.2979363162086217e-11
C46_71 V46 V71 -1.5208167652070542e-20

R46_72 V46 V72 1527.0195925752846
L46_72 V46 V72 -3.279789756185009e-12
C46_72 V46 V72 7.735701235108815e-21

R46_73 V46 V73 55240.75544795044
L46_73 V46 V73 2.9153556851526666e-11
C46_73 V46 V73 1.533225852482724e-19

R46_74 V46 V74 2952.1625893844957
L46_74 V46 V74 4.732844563714841e-12
C46_74 V46 V74 -4.2214908779051624e-20

R46_75 V46 V75 -2608.4028722214825
L46_75 V46 V75 3.972368618700134e-12
C46_75 V46 V75 5.3485117998900246e-20

R46_76 V46 V76 -2206.8090656647128
L46_76 V46 V76 3.485097258298165e-12
C46_76 V46 V76 1.3506309228594534e-19

R46_77 V46 V77 -5307.628263283821
L46_77 V46 V77 5.48305077459202e-11
C46_77 V46 V77 1.9210063789623206e-20

R46_78 V46 V78 -17222.58803679997
L46_78 V46 V78 -4.788407113363975e-12
C46_78 V46 V78 -1.7880246786448426e-20

R46_79 V46 V79 16754.033999519204
L46_79 V46 V79 -1.8854183556295065e-11
C46_79 V46 V79 -6.708958925887737e-21

R46_80 V46 V80 5730.450562536759
L46_80 V46 V80 -9.192809825589854e-12
C46_80 V46 V80 2.1387266962709207e-20

R46_81 V46 V81 12615.966308845533
L46_81 V46 V81 3.3518687333567174e-12
C46_81 V46 V81 5.956832849896642e-20

R46_82 V46 V82 14075.776091815796
L46_82 V46 V82 5.792042534335672e-12
C46_82 V46 V82 8.166678962009447e-21

R46_83 V46 V83 20309.801202024384
L46_83 V46 V83 2.5971466113539833e-11
C46_83 V46 V83 1.7293630134183768e-20

R46_84 V46 V84 -7747.494019434174
L46_84 V46 V84 -3.77255811806965e-11
C46_84 V46 V84 1.0920047627833718e-20

R46_85 V46 V85 14185.027707820358
L46_85 V46 V85 4.4809556920684004e-11
C46_85 V46 V85 3.893624957372223e-20

R46_86 V46 V86 -76582.82982059388
L46_86 V46 V86 -2.7901028389140225e-11
C46_86 V46 V86 -1.0158329344312541e-20

R46_87 V46 V87 -67089.39288960204
L46_87 V46 V87 2.7217711591528816e-11
C46_87 V46 V87 4.0807602829992326e-20

R46_88 V46 V88 11898.32288396677
L46_88 V46 V88 1.1539458622591376e-11
C46_88 V46 V88 4.521610611971888e-20

R46_89 V46 V89 -16971.030373907466
L46_89 V46 V89 2.2262626790159753e-11
C46_89 V46 V89 1.6224595852817278e-20

R46_90 V46 V90 16816.126306905742
L46_90 V46 V90 1.3756995955418164e-11
C46_90 V46 V90 3.779699305198158e-20

R46_91 V46 V91 21610.00340582502
L46_91 V46 V91 3.8718974634079065e-12
C46_91 V46 V91 3.4122036586964276e-20

R46_92 V46 V92 -53408.43246726883
L46_92 V46 V92 -7.473616695937627e-12
C46_92 V46 V92 5.2623748268973815e-21

R46_93 V46 V93 2654.2684198523584
L46_93 V46 V93 9.431419200324227e-11
C46_93 V46 V93 4.527940892147848e-21

R46_94 V46 V94 4873.203380330225
L46_94 V46 V94 -5.458257387327025e-10
C46_94 V46 V94 1.0563690077288873e-20

R46_95 V46 V95 -31116.49668120447
L46_95 V46 V95 1.1554699065922839e-11
C46_95 V46 V95 -1.2492714404489045e-20

R46_96 V46 V96 -5423.0316439269745
L46_96 V46 V96 -3.527503768681309e-12
C46_96 V46 V96 -1.0274643330961452e-19

R46_97 V46 V97 6059.288009541803
L46_97 V46 V97 1.8030910124825273e-11
C46_97 V46 V97 7.346442920971402e-23

R46_98 V46 V98 5093.920771944323
L46_98 V46 V98 -5.5379430729774526e-11
C46_98 V46 V98 -3.0991114744592256e-21

R46_99 V46 V99 6597.321422949368
L46_99 V46 V99 2.121041788436649e-10
C46_99 V46 V99 1.8271122428980318e-20

R46_100 V46 V100 -20547.604442382108
L46_100 V46 V100 9.037632094658237e-12
C46_100 V46 V100 1.8963299919675144e-20

R46_101 V46 V101 5308.099041866806
L46_101 V46 V101 -1.8192427912055043e-11
C46_101 V46 V101 -1.1992715514060598e-20

R46_102 V46 V102 4714.751183391303
L46_102 V46 V102 1.6793222357232494e-11
C46_102 V46 V102 8.135316126948716e-20

R46_103 V46 V103 8700.440134000837
L46_103 V46 V103 1.469980705952606e-11
C46_103 V46 V103 6.989904533405963e-20

R46_104 V46 V104 -13332.313475796547
L46_104 V46 V104 -4.602006721218854e-12
C46_104 V46 V104 -5.800566740902628e-20

R46_105 V46 V105 -4604.313261462441
L46_105 V46 V105 3.107540930337244e-11
C46_105 V46 V105 6.79441539893655e-22

R46_106 V46 V106 -5301.497814318316
L46_106 V46 V106 2.1224271666130214e-11
C46_106 V46 V106 -5.579883740602692e-20

R46_107 V46 V107 17352.938767568136
L46_107 V46 V107 1.857686468444823e-11
C46_107 V46 V107 4.920444332742326e-21

R46_108 V46 V108 -7063.082286659454
L46_108 V46 V108 1.3649139768319553e-11
C46_108 V46 V108 -4.7429201481150793e-20

R46_109 V46 V109 -28752.232410142376
L46_109 V46 V109 -5.80752041966149e-12
C46_109 V46 V109 -6.400746693370124e-20

R46_110 V46 V110 -18766.18325174671
L46_110 V46 V110 -2.490962699654008e-11
C46_110 V46 V110 3.6199472728367003e-20

R46_111 V46 V111 -54012.41369547911
L46_111 V46 V111 1.8408705060088206e-11
C46_111 V46 V111 4.384714275619236e-20

R46_112 V46 V112 -12451.42779081455
L46_112 V46 V112 -1.2907515900147612e-10
C46_112 V46 V112 1.0246765869127762e-20

R46_113 V46 V113 -6995.053730901558
L46_113 V46 V113 1.2933340052009669e-11
C46_113 V46 V113 -3.1999574663955754e-21

R46_114 V46 V114 -23095.866538296887
L46_114 V46 V114 4.0928230380701116e-10
C46_114 V46 V114 -6.701020357351988e-20

R46_115 V46 V115 24325.85778297363
L46_115 V46 V115 1.2895736431232632e-11
C46_115 V46 V115 3.1455254771014454e-20

R46_116 V46 V116 -60648.05155150271
L46_116 V46 V116 2.4234399042581765e-11
C46_116 V46 V116 -5.921111885324399e-20

R46_117 V46 V117 10588.44210456076
L46_117 V46 V117 -1.7460164838273894e-11
C46_117 V46 V117 -4.5521739898636805e-20

R46_118 V46 V118 -9089.626671357304
L46_118 V46 V118 -8.614719773624148e-12
C46_118 V46 V118 -5.124672004840455e-21

R46_119 V46 V119 -7839.769644436443
L46_119 V46 V119 -9.427324816547145e-11
C46_119 V46 V119 1.0466398344151057e-20

R46_120 V46 V120 7954.306018530766
L46_120 V46 V120 2.2422131034371003e-11
C46_120 V46 V120 2.5709986056910097e-20

R46_121 V46 V121 -7106.872840103944
L46_121 V46 V121 3.96241001389227e-11
C46_121 V46 V121 1.080244471077721e-20

R46_122 V46 V122 -2511.929194898338
L46_122 V46 V122 1.2649158740231737e-11
C46_122 V46 V122 -2.109281474314527e-20

R46_123 V46 V123 58575.291780198415
L46_123 V46 V123 -3.5127759648286104e-11
C46_123 V46 V123 -1.7882576340176382e-20

R46_124 V46 V124 14928.617272077438
L46_124 V46 V124 2.197159578388396e-10
C46_124 V46 V124 3.667563806529883e-20

R46_125 V46 V125 4466.545111611077
L46_125 V46 V125 4.3578684773730744e-11
C46_125 V46 V125 -7.576245674291192e-21

R46_126 V46 V126 2865.1121681559353
L46_126 V46 V126 -1.0771360800312055e-11
C46_126 V46 V126 -1.2618517972766381e-20

R46_127 V46 V127 -16631.766496242286
L46_127 V46 V127 1.4231870591552768e-11
C46_127 V46 V127 3.8889982438278366e-20

R46_128 V46 V128 8925.370789334303
L46_128 V46 V128 -9.072360396122445e-11
C46_128 V46 V128 2.996326392220112e-20

R46_129 V46 V129 12006.940468774463
L46_129 V46 V129 4.937083263087079e-11
C46_129 V46 V129 3.347913826181115e-20

R46_130 V46 V130 7991.518546408562
L46_130 V46 V130 -5.887746783081493e-11
C46_130 V46 V130 4.494659516692877e-20

R46_131 V46 V131 7231.826094944314
L46_131 V46 V131 -1.70775163310625e-11
C46_131 V46 V131 -4.210474925930876e-21

R46_132 V46 V132 40405.742548563576
L46_132 V46 V132 2.3797889698743604e-11
C46_132 V46 V132 -1.5329599119383289e-21

R46_133 V46 V133 -31980.862812886964
L46_133 V46 V133 2.1094111957512773e-11
C46_133 V46 V133 -3.927234524066008e-22

R46_134 V46 V134 -8715.657026597204
L46_134 V46 V134 1.1003051343662025e-10
C46_134 V46 V134 5.1666098242434477e-20

R46_135 V46 V135 -7429.8402861618715
L46_135 V46 V135 4.104574962505117e-11
C46_135 V46 V135 -4.20410462159113e-21

R46_136 V46 V136 18067.31077634035
L46_136 V46 V136 -2.992350782266549e-11
C46_136 V46 V136 -7.322145558864947e-21

R46_137 V46 V137 3232.990311321537
L46_137 V46 V137 -2.3310986515947624e-11
C46_137 V46 V137 5.126590837965206e-20

R46_138 V46 V138 2792.4861709857937
L46_138 V46 V138 -1.511533018648774e-11
C46_138 V46 V138 5.82892560308116e-20

R46_139 V46 V139 -11277.905105107933
L46_139 V46 V139 1.869393252795057e-11
C46_139 V46 V139 -5.1832547551393745e-20

R46_140 V46 V140 -6305.5558050943
L46_140 V46 V140 9.156941438014341e-10
C46_140 V46 V140 -3.7331747804259966e-20

R46_141 V46 V141 5748.4470244663735
L46_141 V46 V141 6.336461600172296e-10
C46_141 V46 V141 2.5040124173141344e-20

R46_142 V46 V142 -4678.389233391981
L46_142 V46 V142 -3.5869672754524925e-11
C46_142 V46 V142 -5.029444150091227e-20

R46_143 V46 V143 24763.752495300854
L46_143 V46 V143 -2.070934462290761e-11
C46_143 V46 V143 -1.358770166339697e-20

R46_144 V46 V144 -7220.187064478743
L46_144 V46 V144 1.2332944934131858e-11
C46_144 V46 V144 7.072028304936343e-20

R47_47 V47 0 102.57229814789527
L47_47 V47 0 1.6980056209549814e-13
C47_47 V47 0 -7.147427552622363e-19

R47_48 V47 V48 -1868.9529800656064
L47_48 V47 V48 1.4207137385143032e-11
C47_48 V47 V48 -2.4716758357420522e-19

R47_49 V47 V49 837.3538158160825
L47_49 V47 V49 5.8922320807947785e-12
C47_49 V47 V49 -1.276848700693052e-19

R47_50 V47 V50 -1105.0700578026212
L47_50 V47 V50 -2.6438296846023866e-12
C47_50 V47 V50 2.925158566389758e-19

R47_51 V47 V51 1989.2493295654403
L47_51 V47 V51 1.298325507503704e-11
C47_51 V47 V51 2.369448175562672e-19

R47_52 V47 V52 1636.988579966059
L47_52 V47 V52 -2.7867622058370874e-12
C47_52 V47 V52 2.4584640619188005e-19

R47_53 V47 V53 -1152.6163568011161
L47_53 V47 V53 -6.6153460115027144e-12
C47_53 V47 V53 1.6613965790304216e-19

R47_54 V47 V54 -1319.4280210206311
L47_54 V47 V54 -6.263112986204172e-12
C47_54 V47 V54 -2.213136259324448e-19

R47_55 V47 V55 5735.158805424207
L47_55 V47 V55 -2.6580182719003966e-12
C47_55 V47 V55 -1.2542007521932065e-19

R47_56 V47 V56 -1666.8580806162918
L47_56 V47 V56 -2.3370840267323968e-12
C47_56 V47 V56 -8.592373340229158e-20

R47_57 V47 V57 -225.02009495973698
L47_57 V47 V57 -1.4550979051224696e-12
C47_57 V47 V57 -2.920768305268922e-20

R47_58 V47 V58 275.6454691182696
L47_58 V47 V58 5.93521132774262e-12
C47_58 V47 V58 -1.3003053984613341e-19

R47_59 V47 V59 -552.8994290066695
L47_59 V47 V59 -6.096396578138363e-13
C47_59 V47 V59 -8.445326738219105e-20

R47_60 V47 V60 -618.4040462279734
L47_60 V47 V60 -1.6318938581082635e-12
C47_60 V47 V60 -1.0728178652946131e-20

R47_61 V47 V61 799.6994248145097
L47_61 V47 V61 4.428612144570495e-12
C47_61 V47 V61 1.1913284121778842e-19

R47_62 V47 V62 2506.1316891250412
L47_62 V47 V62 -1.9056015856453467e-12
C47_62 V47 V62 1.9547506242448973e-19

R47_63 V47 V63 797.6636285762481
L47_63 V47 V63 -9.194960522586212e-12
C47_63 V47 V63 -1.5056136657655194e-19

R47_64 V47 V64 -3856.551202198208
L47_64 V47 V64 -3.3257636306204344e-12
C47_64 V47 V64 -8.258512710138977e-20

R47_65 V47 V65 -596.2040513690995
L47_65 V47 V65 -5.384122042942186e-12
C47_65 V47 V65 1.095890646675333e-19

R47_66 V47 V66 -1709.5993100626224
L47_66 V47 V66 -7.1341600494775066e-12
C47_66 V47 V66 -6.386681214399322e-20

R47_67 V47 V67 -646.3126130788926
L47_67 V47 V67 -1.6096919059253513e-12
C47_67 V47 V67 -1.4631304855880388e-20

R47_68 V47 V68 -4820.816264009468
L47_68 V47 V68 7.294773432595927e-11
C47_68 V47 V68 8.538345726202155e-21

R47_69 V47 V69 1880.6971445172032
L47_69 V47 V69 1.4219609832550738e-12
C47_69 V47 V69 3.037776091322421e-20

R47_70 V47 V70 -87128.16765503431
L47_70 V47 V70 -2.525181491172157e-12
C47_70 V47 V70 -6.757406166476876e-20

R47_71 V47 V71 4818.4446114118655
L47_71 V47 V71 6.115377562266666e-12
C47_71 V47 V71 5.487832809543847e-20

R47_72 V47 V72 4811.059459600367
L47_72 V47 V72 -4.190839135391675e-12
C47_72 V47 V72 -4.5357428322660275e-20

R47_73 V47 V73 15764.092474982026
L47_73 V47 V73 -5.777387688128781e-12
C47_73 V47 V73 -1.9820112509939154e-20

R47_74 V47 V74 2451.0663180315105
L47_74 V47 V74 9.709144743259772e-12
C47_74 V47 V74 -4.2620177191099694e-20

R47_75 V47 V75 -3501.888922648421
L47_75 V47 V75 7.511610655865967e-12
C47_75 V47 V75 6.29258596829299e-20

R47_76 V47 V76 -21903.182154707578
L47_76 V47 V76 -8.852921687040807e-12
C47_76 V47 V76 -4.5035211152992585e-20

R47_77 V47 V77 10448.564024193898
L47_77 V47 V77 2.077907406315367e-11
C47_77 V47 V77 3.0650545269071216e-20

R47_78 V47 V78 28224.68540330349
L47_78 V47 V78 -4.748798645268292e-12
C47_78 V47 V78 -1.022048382759497e-20

R47_79 V47 V79 5594.840891922161
L47_79 V47 V79 -8.974002433862189e-12
C47_79 V47 V79 -8.567987973329439e-20

R47_80 V47 V80 11684.36203633366
L47_80 V47 V80 1.1188018742006887e-11
C47_80 V47 V80 7.84081124097394e-20

R47_81 V47 V81 -64436.33496544469
L47_81 V47 V81 -1.3723523518197875e-11
C47_81 V47 V81 -4.207908951768794e-22

R47_82 V47 V82 14243.23024848169
L47_82 V47 V82 7.225309590355301e-12
C47_82 V47 V82 -2.2194928049366403e-20

R47_83 V47 V83 -44653.556747132825
L47_83 V47 V83 5.815305377132741e-12
C47_83 V47 V83 6.509034378145347e-20

R47_84 V47 V84 14561.011498055821
L47_84 V47 V84 -6.2143774803470415e-12
C47_84 V47 V84 -9.15371051377235e-20

R47_85 V47 V85 11231.980718979234
L47_85 V47 V85 -5.328851223986678e-12
C47_85 V47 V85 -1.0427621251166494e-19

R47_86 V47 V86 16309.59200525712
L47_86 V47 V86 -9.18969427174923e-12
C47_86 V47 V86 -1.6768816046952254e-20

R47_87 V47 V87 -85613.65456081521
L47_87 V47 V87 -8.165247612783736e-12
C47_87 V47 V87 -5.426781184630807e-20

R47_88 V47 V88 -30828.974066702096
L47_88 V47 V88 -5.133694473937011e-11
C47_88 V47 V88 1.354346828322948e-20

R47_89 V47 V89 -25212.840832700756
L47_89 V47 V89 1.2312481222737924e-11
C47_89 V47 V89 1.4508232755682102e-20

R47_90 V47 V90 45754.448584118276
L47_90 V47 V90 8.219443594248286e-12
C47_90 V47 V90 1.326328663699279e-19

R47_91 V47 V91 134758.47227074558
L47_91 V47 V91 7.260652034121945e-12
C47_91 V47 V91 1.1560770054568723e-20

R47_92 V47 V92 25984.849173673585
L47_92 V47 V92 1.1139850104486631e-11
C47_92 V47 V92 2.2335816770801375e-20

R47_93 V47 V93 3904.979329297779
L47_93 V47 V93 -3.0492786374714054e-11
C47_93 V47 V93 -9.8866571130637e-21

R47_94 V47 V94 32720.468593999743
L47_94 V47 V94 -3.0404311368451636e-10
C47_94 V47 V94 5.511727566467855e-20

R47_95 V47 V95 13673.360670146543
L47_95 V47 V95 1.3591685730393686e-11
C47_95 V47 V95 9.60061933910789e-21

R47_96 V47 V96 -16551.615453991042
L47_96 V47 V96 1.4813537601205372e-11
C47_96 V47 V96 1.460509943100921e-20

R47_97 V47 V97 10807.469717485736
L47_97 V47 V97 3.6192141518238575e-11
C47_97 V47 V97 7.4500717213726e-20

R47_98 V47 V98 4611.907966986902
L47_98 V47 V98 7.935411794005512e-12
C47_98 V47 V98 4.3776970619726884e-20

R47_99 V47 V99 16849.53781782712
L47_99 V47 V99 -3.330455613338753e-11
C47_99 V47 V99 -1.4239262445168457e-20

R47_100 V47 V100 -17645.2403781556
L47_100 V47 V100 -3.336275596044429e-11
C47_100 V47 V100 2.174253574811814e-21

R47_101 V47 V101 13447.559519866025
L47_101 V47 V101 8.008539706837438e-12
C47_101 V47 V101 4.1817638596978957e-20

R47_102 V47 V102 3938.574521374944
L47_102 V47 V102 3.1435895002958375e-12
C47_102 V47 V102 3.2291973136656035e-19

R47_103 V47 V103 -22873.87192583665
L47_103 V47 V103 -5.8700080986449615e-12
C47_103 V47 V103 -1.9732921847215108e-19

R47_104 V47 V104 -405225.1646437965
L47_104 V47 V104 2.4326981299300856e-10
C47_104 V47 V104 1.0757549328462057e-20

R47_105 V47 V105 -11440.164312291701
L47_105 V47 V105 -6.140900941723377e-12
C47_105 V47 V105 -9.351258549137866e-20

R47_106 V47 V106 -10689.98263698839
L47_106 V47 V106 3.989463853221691e-12
C47_106 V47 V106 1.556310402747845e-19

R47_107 V47 V107 10708.98969107395
L47_107 V47 V107 5.474091695337619e-12
C47_107 V47 V107 2.27149676079933e-19

R47_108 V47 V108 33816.00429987641
L47_108 V47 V108 -5.504299363404656e-12
C47_108 V47 V108 -2.0648750603973716e-19

R47_109 V47 V109 214965.53481708674
L47_109 V47 V109 -1.719107966079049e-11
C47_109 V47 V109 -9.321206890789635e-20

R47_110 V47 V110 10204.533914612186
L47_110 V47 V110 -8.191904990913837e-12
C47_110 V47 V110 -4.7862803840553693e-20

R47_111 V47 V111 -5571.315537037231
L47_111 V47 V111 -7.950283151461846e-12
C47_111 V47 V111 -1.0247284563261009e-19

R47_112 V47 V112 6054.173036829147
L47_112 V47 V112 3.920969714492078e-12
C47_112 V47 V112 1.800203432723438e-19

R47_113 V47 V113 24307.197409675675
L47_113 V47 V113 9.13166581445895e-12
C47_113 V47 V113 6.922409160286565e-20

R47_114 V47 V114 38930.01571100259
L47_114 V47 V114 8.905168830244232e-12
C47_114 V47 V114 3.535156467968431e-20

R47_115 V47 V115 3872.601411124421
L47_115 V47 V115 9.904033843112771e-12
C47_115 V47 V115 1.1453765419133634e-19

R47_116 V47 V116 -15197.719993081144
L47_116 V47 V116 -9.115875147047214e-12
C47_116 V47 V116 -9.577262159293495e-20

R47_117 V47 V117 17801.977567473394
L47_117 V47 V117 -1.505243803652117e-11
C47_117 V47 V117 -9.259413626438923e-20

R47_118 V47 V118 -11201.60229689388
L47_118 V47 V118 -9.168546515899827e-12
C47_118 V47 V118 -4.454838206196146e-20

R47_119 V47 V119 -6375.768331982408
L47_119 V47 V119 -8.288506390060063e-12
C47_119 V47 V119 -4.234934571970173e-20

R47_120 V47 V120 3628.21769050007
L47_120 V47 V120 2.0773412180838395e-11
C47_120 V47 V120 -2.5849065824566638e-20

R47_121 V47 V121 -53691.80701331464
L47_121 V47 V121 1.584355566247003e-11
C47_121 V47 V121 1.8229724140286862e-20

R47_122 V47 V122 3879.5647749909253
L47_122 V47 V122 6.305247516847179e-12
C47_122 V47 V122 -4.776128294743938e-21

R47_123 V47 V123 17000.12474146946
L47_123 V47 V123 5.655697856101907e-11
C47_123 V47 V123 -3.2546275589275632e-21

R47_124 V47 V124 103318.67987228368
L47_124 V47 V124 -1.0085875641776654e-10
C47_124 V47 V124 6.090893846895599e-21

R47_125 V47 V125 5206.397473435353
L47_125 V47 V125 -3.9839046806046426e-11
C47_125 V47 V125 -1.0162632941277142e-20

R47_126 V47 V126 -3312.159380690534
L47_126 V47 V126 -8.811171217440989e-12
C47_126 V47 V126 4.9218961978778564e-20

R47_127 V47 V127 2953.869024221602
L47_127 V47 V127 7.834797208104732e-12
C47_127 V47 V127 2.0280065967782784e-21

R47_128 V47 V128 13762.458386584325
L47_128 V47 V128 6.615308562912755e-11
C47_128 V47 V128 1.7637480411363497e-21

R47_129 V47 V129 5576.991050473409
L47_129 V47 V129 4.7383329057564434e-11
C47_129 V47 V129 -5.9066834151660705e-21

R47_130 V47 V130 -41486.11424824292
L47_130 V47 V130 -9.645375870873221e-12
C47_130 V47 V130 -7.522761128898325e-20

R47_131 V47 V131 -89699.14156951263
L47_131 V47 V131 2.3002104887663288e-11
C47_131 V47 V131 8.423092539058648e-20

R47_132 V47 V132 -10853.04355511566
L47_132 V47 V132 -3.2903322306599e-11
C47_132 V47 V132 1.5167880146156996e-21

R47_133 V47 V133 -18852.710933920556
L47_133 V47 V133 1.0178422486906866e-11
C47_133 V47 V133 5.86498705283833e-20

R47_134 V47 V134 -6520.085951232236
L47_134 V47 V134 -3.545122182332567e-11
C47_134 V47 V134 1.5273329429369974e-20

R47_135 V47 V135 8822.481384373245
L47_135 V47 V135 1.092155936680142e-11
C47_135 V47 V135 -1.494240107655256e-20

R47_136 V47 V136 37272.68569516157
L47_136 V47 V136 1.3894627860506393e-10
C47_136 V47 V136 9.799770404303575e-21

R47_137 V47 V137 6005.439806055199
L47_137 V47 V137 -1.4026436656626166e-11
C47_137 V47 V137 -2.312805173077228e-20

R47_138 V47 V138 -2953.608608825475
L47_138 V47 V138 -5.40697349569959e-12
C47_138 V47 V138 -1.963540997341471e-20

R47_139 V47 V139 1890.7475062763417
L47_139 V47 V139 4.72999049069209e-12
C47_139 V47 V139 3.0095100543518924e-20

R47_140 V47 V140 -7026.725422130074
L47_140 V47 V140 -1.0906423453115444e-11
C47_140 V47 V140 -3.752675617783662e-20

R47_141 V47 V141 -80243.55557589539
L47_141 V47 V141 -2.5125264452974738e-11
C47_141 V47 V141 -2.2806808949209826e-21

R47_142 V47 V142 -5298.8031166518185
L47_142 V47 V142 -1.6296386985829174e-11
C47_142 V47 V142 -3.7886183215368073e-20

R47_143 V47 V143 -8498.259504843469
L47_143 V47 V143 -2.7152795742535873e-10
C47_143 V47 V143 2.564229156192956e-20

R47_144 V47 V144 -8375.067632728886
L47_144 V47 V144 2.6715339503603687e-11
C47_144 V47 V144 -1.6401157977067573e-21

R48_48 V48 0 -886.4552497120453
L48_48 V48 0 -3.291481489612017e-13
C48_48 V48 0 -5.049662099220848e-19

R48_49 V48 V49 -1472.0901888295487
L48_49 V48 V49 -4.496148331213668e-11
C48_49 V48 V49 -3.425900890302995e-20

R48_50 V48 V50 1182.339503297865
L48_50 V48 V50 2.739802859579149e-12
C48_50 V48 V50 1.210029632939311e-19

R48_51 V48 V51 -5043.655888588929
L48_51 V48 V51 -2.2134988263616374e-12
C48_51 V48 V51 2.5955240418118747e-20

R48_52 V48 V52 1841.27580257757
L48_52 V48 V52 2.6534854716531675e-12
C48_52 V48 V52 1.5331787282270632e-19

R48_53 V48 V53 -1998.0076305357786
L48_53 V48 V53 4.928546250609127e-12
C48_53 V48 V53 -8.854777495642165e-20

R48_54 V48 V54 -18926.80603655127
L48_54 V48 V54 4.644406862910109e-12
C48_54 V48 V54 -1.1208735840322457e-19

R48_55 V48 V55 -19981.730377202828
L48_55 V48 V55 3.877921361423725e-12
C48_55 V48 V55 -1.0166847975234398e-19

R48_56 V48 V56 1578.4050491773762
L48_56 V48 V56 -4.451882441147287e-12
C48_56 V48 V56 2.1038652179799582e-19

R48_57 V48 V57 732.6383950643249
L48_57 V48 V57 9.053405859068912e-13
C48_57 V48 V57 9.824225928234877e-21

R48_58 V48 V58 466.1767159627823
L48_58 V48 V58 1.443822624600319e-12
C48_58 V48 V58 -7.187959718142041e-20

R48_59 V48 V59 901.2395578752353
L48_59 V48 V59 3.6488477875146284e-12
C48_59 V48 V59 -1.5512453002646266e-20

R48_60 V48 V60 -385.61368951860624
L48_60 V48 V60 -2.3062129354672337e-12
C48_60 V48 V60 -2.5469815739313102e-20

R48_61 V48 V61 -2209.5599464910674
L48_61 V48 V61 -7.0785818141198714e-12
C48_61 V48 V61 1.5505792452493558e-20

R48_62 V48 V62 -1745.1454960720152
L48_62 V48 V62 -1.581788059484451e-11
C48_62 V48 V62 1.0547589863482134e-19

R48_63 V48 V63 3105.399589322937
L48_63 V48 V63 5.3806241651714745e-11
C48_63 V48 V63 -7.638168744290232e-20

R48_64 V48 V64 2956.228093277658
L48_64 V48 V64 1.0669312761250698e-11
C48_64 V48 V64 1.5987915036024115e-19

R48_65 V48 V65 1840.8402393554622
L48_65 V48 V65 1.940102726130009e-12
C48_65 V48 V65 5.344449040778053e-20

R48_66 V48 V66 1695.8460983843158
L48_66 V48 V66 2.1314951408470603e-12
C48_66 V48 V66 -2.270179242790436e-20

R48_67 V48 V67 -4355.151181050757
L48_67 V48 V67 -9.426493483240878e-12
C48_67 V48 V67 -2.2069319962159582e-20

R48_68 V48 V68 -1046.2710568834696
L48_68 V48 V68 -2.923397893583777e-12
C48_68 V48 V68 3.379117053239459e-20

R48_69 V48 V69 -16755.93520425296
L48_69 V48 V69 -9.347455285969223e-12
C48_69 V48 V69 1.9196131408446067e-20

R48_70 V48 V70 -6076.5809178379595
L48_70 V48 V70 -2.973016495481699e-11
C48_70 V48 V70 -8.340699378148953e-20

R48_71 V48 V71 -26934.169009579586
L48_71 V48 V71 1.0568966886420153e-11
C48_71 V48 V71 1.0708556794609885e-20

R48_72 V48 V72 17317.495847727547
L48_72 V48 V72 -1.3689611345886158e-11
C48_72 V48 V72 -4.732698276238752e-20

R48_73 V48 V73 -4840.207575071459
L48_73 V48 V73 -1.423698618314759e-11
C48_73 V48 V73 1.400093694089645e-20

R48_74 V48 V74 -8486.965526713895
L48_74 V48 V74 -6.87196368418678e-12
C48_74 V48 V74 -4.350422859407915e-21

R48_75 V48 V75 16294.39660884987
L48_75 V48 V75 9.678337193524674e-12
C48_75 V48 V75 4.3812984045867416e-20

R48_76 V48 V76 5799.1371223128335
L48_76 V48 V76 6.1456109720580545e-12
C48_76 V48 V76 9.789799069719346e-21

R48_77 V48 V77 8474.050815492155
L48_77 V48 V77 -1.5354562749926435e-11
C48_77 V48 V77 -6.735365662551461e-20

R48_78 V48 V78 74806.0565419197
L48_78 V48 V78 -2.3726547544445958e-11
C48_78 V48 V78 -8.027360433133425e-20

R48_79 V48 V79 169956.45323345342
L48_79 V48 V79 -3.2672555912376116e-11
C48_79 V48 V79 -4.190564172134546e-20

R48_80 V48 V80 -66388.47312932735
L48_80 V48 V80 -8.525713281639005e-12
C48_80 V48 V80 2.368805575328021e-21

R48_81 V48 V81 -72296.72974039415
L48_81 V48 V81 3.4431427958710094e-12
C48_81 V48 V81 1.0512748440504057e-19

R48_82 V48 V82 31829.01257478297
L48_82 V48 V82 7.1562869923964515e-12
C48_82 V48 V82 1.7057328357212708e-19

R48_83 V48 V83 150086.53350051545
L48_83 V48 V83 1.6184465318812018e-11
C48_83 V48 V83 1.153498692925609e-19

R48_84 V48 V84 8949.629027577637
L48_84 V48 V84 -1.4540067229796492e-11
C48_84 V48 V84 -5.802300305884437e-20

R48_85 V48 V85 -52739.327420035406
L48_85 V48 V85 -1.8257168776390877e-11
C48_85 V48 V85 -7.088119316273676e-20

R48_86 V48 V86 -11780.235758841112
L48_86 V48 V86 -1.0445591890465089e-11
C48_86 V48 V86 -4.607178180733709e-20

R48_87 V48 V87 -21406.42722866266
L48_87 V48 V87 -1.5586240389736177e-11
C48_87 V48 V87 -1.014205463500734e-19

R48_88 V48 V88 -62942.65487912244
L48_88 V48 V88 2.611717348820172e-11
C48_88 V48 V88 -9.36006862410698e-21

R48_89 V48 V89 28491.571054195232
L48_89 V48 V89 1.1890770623206944e-10
C48_89 V48 V89 3.587887338850893e-20

R48_90 V48 V90 -60293.680722574725
L48_90 V48 V90 1.0672833608674467e-11
C48_90 V48 V90 6.866735385090385e-20

R48_91 V48 V91 15041.899324369995
L48_91 V48 V91 4.784787928359098e-12
C48_91 V48 V91 1.5365961846881793e-19

R48_92 V48 V92 -86505.10974920625
L48_92 V48 V92 -6.8284461576477156e-12
C48_92 V48 V92 1.4266612277908006e-20

R48_93 V48 V93 -19954.646026878472
L48_93 V48 V93 -9.292677844576722e-11
C48_93 V48 V93 -1.388517349995206e-20

R48_94 V48 V94 -19169.190922936497
L48_94 V48 V94 2.154007103090478e-11
C48_94 V48 V94 -7.4527436597987565e-22

R48_95 V48 V95 14030.368307293884
L48_95 V48 V95 1.0189187635855281e-11
C48_95 V48 V95 9.161823964129807e-20

R48_96 V48 V96 15776.152335585986
L48_96 V48 V96 -3.828937250658807e-12
C48_96 V48 V96 -6.220562890721815e-20

R48_97 V48 V97 -36702.656885334334
L48_97 V48 V97 1.0690223071697358e-11
C48_97 V48 V97 1.0277555171028555e-20

R48_98 V48 V98 325481.3678789775
L48_98 V48 V98 2.0797636601988233e-11
C48_98 V48 V98 6.234579407530671e-20

R48_99 V48 V99 -24383.40600544851
L48_99 V48 V99 -8.344792558655977e-11
C48_99 V48 V99 -8.900145883036296e-21

R48_100 V48 V100 19026.365177467746
L48_100 V48 V100 9.127688517317364e-12
C48_100 V48 V100 1.62472753304612e-20

R48_101 V48 V101 -61468.71083110287
L48_101 V48 V101 -4.847966517965744e-09
C48_101 V48 V101 5.1688317419403815e-20

R48_102 V48 V102 49084.293268976384
L48_102 V48 V102 4.064499349721755e-12
C48_102 V48 V102 2.0182682768342274e-19

R48_103 V48 V103 -12467.300542381663
L48_103 V48 V103 -1.2457417741434035e-11
C48_103 V48 V103 -9.247835861330868e-20

R48_104 V48 V104 -38923.164115448126
L48_104 V48 V104 -3.904041903327669e-12
C48_104 V48 V104 -9.869806283345733e-20

R48_105 V48 V105 15505.621915872343
L48_105 V48 V105 -3.698994469837345e-11
C48_105 V48 V105 -8.34146803956067e-20

R48_106 V48 V106 8831.64593979092
L48_106 V48 V106 7.53267204173077e-12
C48_106 V48 V106 1.9484140732014473e-19

R48_107 V48 V107 18413.079153497412
L48_107 V48 V107 6.571430160902586e-12
C48_107 V48 V107 1.5377510275877994e-19

R48_108 V48 V108 14908.516729208832
L48_108 V48 V108 -4.1446894297724016e-11
C48_108 V48 V108 -1.0985851357954913e-19

R48_109 V48 V109 -11059.847403836598
L48_109 V48 V109 -4.3066561840838386e-12
C48_109 V48 V109 -1.085765357860687e-19

R48_110 V48 V110 -26899.36898343192
L48_110 V48 V110 -1.0232605727954803e-11
C48_110 V48 V110 -1.617140592449417e-19

R48_111 V48 V111 -15214.129505628278
L48_111 V48 V111 -1.1097104530459627e-11
C48_111 V48 V111 -1.0123668113451509e-19

R48_112 V48 V112 15144.344289212231
L48_112 V48 V112 6.820919591134918e-12
C48_112 V48 V112 1.3311109086335227e-19

R48_113 V48 V113 7625.972598898026
L48_113 V48 V113 9.198752546603617e-12
C48_113 V48 V113 4.0182763800723995e-20

R48_114 V48 V114 15413.112557329534
L48_114 V48 V114 8.818930712355033e-12
C48_114 V48 V114 1.181824875720392e-19

R48_115 V48 V115 18125.771892289762
L48_115 V48 V115 1.3251496064972829e-11
C48_115 V48 V115 8.084459975155885e-20

R48_116 V48 V116 135525.069654537
L48_116 V48 V116 -1.8490049230758855e-11
C48_116 V48 V116 -7.557218173688277e-20

R48_117 V48 V117 -17702.730534575272
L48_117 V48 V117 -1.4884371955506822e-11
C48_117 V48 V117 -5.1619961898057214e-20

R48_118 V48 V118 -21737.331505226375
L48_118 V48 V118 -7.842379005313247e-12
C48_118 V48 V118 -8.317991926065448e-20

R48_119 V48 V119 -55993.416391916755
L48_119 V48 V119 -1.2770403464640034e-11
C48_119 V48 V119 -1.2000954897504648e-19

R48_120 V48 V120 20472.16491703786
L48_120 V48 V120 1.1408621351247653e-11
C48_120 V48 V120 -3.854793635821289e-20

R48_121 V48 V121 159871.9294153288
L48_121 V48 V121 1.4851685762654556e-11
C48_121 V48 V121 2.968696065458338e-20

R48_122 V48 V122 5899.927472944346
L48_122 V48 V122 6.768851790886687e-12
C48_122 V48 V122 -8.59241952573064e-21

R48_123 V48 V123 -75877.86017965192
L48_123 V48 V123 4.631310783871031e-10
C48_123 V48 V123 -3.266282180967515e-20

R48_124 V48 V124 -34225.907799879176
L48_124 V48 V124 2.0026108582647346e-10
C48_124 V48 V124 -2.2618984921630453e-20

R48_125 V48 V125 -69002.48469100532
L48_125 V48 V125 -3.143926358080176e-11
C48_125 V48 V125 -1.6983878565281563e-20

R48_126 V48 V126 -6309.652948914025
L48_126 V48 V126 -6.270366417959342e-12
C48_126 V48 V126 2.3459240645286182e-20

R48_127 V48 V127 9375.395504894526
L48_127 V48 V127 7.729390008227368e-12
C48_127 V48 V127 -8.533278563230732e-21

R48_128 V48 V128 -63292.24697782435
L48_128 V48 V128 2.3141606387466863e-11
C48_128 V48 V128 1.6431178220431347e-20

R48_129 V48 V129 -116147.8652957491
L48_129 V48 V129 2.1997164778597228e-11
C48_129 V48 V129 -1.4008763754393926e-20

R48_130 V48 V130 -16366.057457107776
L48_130 V48 V130 -2.137641599420365e-11
C48_130 V48 V130 -4.226017606440734e-21

R48_131 V48 V131 -33049.783478068384
L48_131 V48 V131 5.97097317478814e-11
C48_131 V48 V131 6.953237509362229e-20

R48_132 V48 V132 -46471.66499792223
L48_132 V48 V132 5.525924815555613e-11
C48_132 V48 V132 2.4105234257283748e-20

R48_133 V48 V133 28918.8316238842
L48_133 V48 V133 -6.441100117319443e-11
C48_133 V48 V133 2.5537489567348824e-20

R48_134 V48 V134 -47602.734553882314
L48_134 V48 V134 -2.4491232696585484e-11
C48_134 V48 V134 4.672286066919429e-22

R48_135 V48 V135 12764.351028423163
L48_135 V48 V135 1.0338221044937515e-11
C48_135 V48 V135 -8.272882637204967e-21

R48_136 V48 V136 -387696.897371919
L48_136 V48 V136 -2.2636436461117813e-11
C48_136 V48 V136 -3.7505479853862555e-20

R48_137 V48 V137 -16770.48621813654
L48_137 V48 V137 1.2589726214481165e-09
C48_137 V48 V137 -1.560136332732423e-20

R48_138 V48 V138 -5743.401826878692
L48_138 V48 V138 -4.371409514222054e-12
C48_138 V48 V138 -5.9402039739826e-20

R48_139 V48 V139 5663.55728350173
L48_139 V48 V139 5.889514442442079e-12
C48_139 V48 V139 6.362592567695064e-21

R48_140 V48 V140 28312.988669403054
L48_140 V48 V140 -1.7189656704674766e-11
C48_140 V48 V140 -1.3853374621542016e-20

R48_141 V48 V141 -11417.780660438595
L48_141 V48 V141 -1.101235762129747e-11
C48_141 V48 V141 -3.171028926399457e-20

R48_142 V48 V142 12803.806281633857
L48_142 V48 V142 -9.86144748166205e-12
C48_142 V48 V142 -4.298414447464283e-20

R48_143 V48 V143 -35848.16764383133
L48_143 V48 V143 -1.6790785875184025e-11
C48_143 V48 V143 -8.055176230525335e-21

R48_144 V48 V144 24256.97590749989
L48_144 V48 V144 6.740805725538533e-11
C48_144 V48 V144 -1.6069027154909061e-21

R49_49 V49 0 -135.255951030648
L49_49 V49 0 1.6091449618941675e-13
C49_49 V49 0 3.7115172741404205e-18

R49_50 V49 V50 740.8106801403608
L49_50 V49 V50 -4.376602372356534e-12
C49_50 V49 V50 -8.492943044020479e-21

R49_51 V49 V51 -12508.404285327708
L49_51 V49 V51 3.7603925755981725e-12
C49_51 V49 V51 2.6858093046875297e-19

R49_52 V49 V52 -4430.364486807394
L49_52 V49 V52 -1.4281723437981814e-12
C49_52 V49 V52 -6.55784823506873e-19

R49_53 V49 V53 45410.48705325697
L49_53 V49 V53 -1.84140363869981e-12
C49_53 V49 V53 -2.7524138184162766e-19

R49_54 V49 V54 3614.9548904025582
L49_54 V49 V54 -4.7872361598119295e-12
C49_54 V49 V54 -1.3110033799192396e-19

R49_55 V49 V55 -1925.8410626588548
L49_55 V49 V55 -3.4555381768450064e-12
C49_55 V49 V55 -4.862556270382082e-19

R49_56 V49 V56 9913.83031759671
L49_56 V49 V56 -8.321615440816396e-12
C49_56 V49 V56 -3.1361566798592387e-19

R49_57 V49 V57 329.62779430586806
L49_57 V49 V57 -1.0570000991944482e-12
C49_57 V49 V57 1.29723045083667e-19

R49_58 V49 V58 2564.9189768916794
L49_58 V49 V58 -2.645825078547105e-12
C49_58 V49 V58 4.479352614470791e-20

R49_59 V49 V59 428.080637503594
L49_59 V49 V59 2.4360596932786646e-12
C49_59 V49 V59 1.354814326120116e-19

R49_60 V49 V60 2768.4697432092803
L49_60 V49 V60 -3.658688256632994e-12
C49_60 V49 V60 1.0975077694330064e-20

R49_61 V49 V61 -840.4418646994309
L49_61 V49 V61 -5.277189795772428e-12
C49_61 V49 V61 -4.367451953062685e-19

R49_62 V49 V62 -4322.176978176267
L49_62 V49 V62 9.956560898643906e-12
C49_62 V49 V62 -3.493780294263289e-19

R49_63 V49 V63 -4472.741435097381
L49_63 V49 V63 1.0508364597703308e-11
C49_63 V49 V63 -1.3241324948560585e-19

R49_64 V49 V64 4713.414144822979
L49_64 V49 V64 -6.7024159628844145e-12
C49_64 V49 V64 -7.434652279509314e-20

R49_65 V49 V65 785.9920374357553
L49_65 V49 V65 -1.105546131845833e-12
C49_65 V49 V65 -2.333115212451193e-20

R49_66 V49 V66 1949.538842224134
L49_66 V49 V66 -7.553925230028275e-13
C49_66 V49 V66 -2.850682840266509e-19

R49_67 V49 V67 2007.0478332038178
L49_67 V49 V67 -5.383449623190699e-12
C49_67 V49 V67 -1.9922053890607062e-19

R49_68 V49 V68 -4933.183174202226
L49_68 V49 V68 -6.0364528383454075e-12
C49_68 V49 V68 -2.5815204985432414e-20

R49_69 V49 V69 -1593.34778812706
L49_69 V49 V69 -3.707027149720045e-11
C49_69 V49 V69 9.956804027273324e-20

R49_70 V49 V70 -364003.6638395544
L49_70 V49 V70 2.745388696092977e-12
C49_70 V49 V70 -1.1196850730973338e-19

R49_71 V49 V71 -3396.0843160668087
L49_71 V49 V71 4.534019096787028e-12
C49_71 V49 V71 -1.6493835930098946e-20

R49_72 V49 V72 -81371.61439544654
L49_72 V49 V72 1.870885789337876e-12
C49_72 V49 V72 -4.258896862191358e-20

R49_73 V49 V73 -1457259.6596615624
L49_73 V49 V73 1.217782404436968e-11
C49_73 V49 V73 -6.828985590124704e-20

R49_74 V49 V74 -3615.4500067229606
L49_74 V49 V74 4.5986427803253765e-12
C49_74 V49 V74 1.071847735680177e-19

R49_75 V49 V75 22711.039363639116
L49_75 V49 V75 -3.677954142340214e-12
C49_75 V49 V75 -1.0954357029203105e-20

R49_76 V49 V76 8078.084309539196
L49_76 V49 V76 -2.266884031226643e-12
C49_76 V49 V76 -8.16602761801994e-20

R49_77 V49 V77 25078.487181955647
L49_77 V49 V77 -1.1092840279567885e-11
C49_77 V49 V77 -5.194048553360782e-21

R49_78 V49 V78 -663340.429837889
L49_78 V49 V78 -3.255195025184428e-12
C49_78 V49 V78 -1.9542406194375126e-19

R49_79 V49 V79 -21803.62676821086
L49_79 V49 V79 1.1664211491555544e-11
C49_79 V49 V79 -3.679061171852636e-21

R49_80 V49 V80 -16979.090115987576
L49_80 V49 V80 5.343590294632824e-12
C49_80 V49 V80 -6.84507787572219e-21

R49_81 V49 V81 -75697.00886488952
L49_81 V49 V81 -3.1591589825303323e-11
C49_81 V49 V81 2.079008500225357e-20

R49_82 V49 V82 27724.287041078966
L49_82 V49 V82 7.127238727505984e-12
C49_82 V49 V82 2.25771282671513e-19

R49_83 V49 V83 -40903.45793682082
L49_83 V49 V83 2.987919597030081e-12
C49_83 V49 V83 1.3955639757316629e-19

R49_84 V49 V84 12171.070617108777
L49_84 V49 V84 6.003400028524153e-12
C49_84 V49 V84 4.022061900770832e-21

R49_85 V49 V85 -58521.255031795365
L49_85 V49 V85 1.9574912751727722e-11
C49_85 V49 V85 -6.412688475314245e-20

R49_86 V49 V86 -42479.84446921611
L49_86 V49 V86 -1.523735662450084e-11
C49_86 V49 V86 -7.25445609128308e-20

R49_87 V49 V87 -10746.349742632849
L49_87 V49 V87 -6.267143212720956e-12
C49_87 V49 V87 -8.375318130699883e-20

R49_88 V49 V88 -46186.611472207005
L49_88 V49 V88 -8.526963438286203e-12
C49_88 V49 V88 -3.177603736251925e-20

R49_89 V49 V89 23367.3013493949
L49_89 V49 V89 2.3001044858242408e-09
C49_89 V49 V89 4.1154441248655906e-20

R49_90 V49 V90 -22503.97915917657
L49_90 V49 V90 1.1252522548047658e-10
C49_90 V49 V90 8.126125041382517e-21

R49_91 V49 V91 13206.120670746002
L49_91 V49 V91 5.6000487772812545e-12
C49_91 V49 V91 1.7603556546660794e-19

R49_92 V49 V92 208758.43909422483
L49_92 V49 V92 5.680600731624142e-12
C49_92 V49 V92 3.8214302734694945e-20

R49_93 V49 V93 -10772.54540467793
L49_93 V49 V93 -5.930536964698665e-11
C49_93 V49 V93 -1.3499765800585772e-20

R49_94 V49 V94 -16589.192368789405
L49_94 V49 V94 -7.318872328061235e-12
C49_94 V49 V94 -7.372170570464918e-20

R49_95 V49 V95 23482.72947832185
L49_95 V49 V95 8.519228986685745e-12
C49_95 V49 V95 1.0902511166705065e-19

R49_96 V49 V96 9866.523130604628
L49_96 V49 V96 6.2089293252923755e-12
C49_96 V49 V96 -4.950205817999491e-21

R49_97 V49 V97 -17323.9019058713
L49_97 V49 V97 -1.301075217161008e-11
C49_97 V49 V97 -5.0275501878743305e-20

R49_98 V49 V98 -9334.723194129128
L49_98 V49 V98 6.21136487093818e-12
C49_98 V49 V98 6.67281371440673e-20

R49_99 V49 V99 -13856.682448615848
L49_99 V49 V99 -2.8612723088344117e-11
C49_99 V49 V99 -1.0489304856105648e-20

R49_100 V49 V100 25931.43369796119
L49_100 V49 V100 -1.3353156773175343e-11
C49_100 V49 V100 -1.535476254220336e-20

R49_101 V49 V101 -44260.22806520364
L49_101 V49 V101 8.439535590402954e-12
C49_101 V49 V101 6.078840748679873e-20

R49_102 V49 V102 -8389.405845589792
L49_102 V49 V102 1.040287084049134e-11
C49_102 V49 V102 6.53550226156138e-20

R49_103 V49 V103 -35075.16002294798
L49_103 V49 V103 -6.203207116483334e-11
C49_103 V49 V103 -1.0075536032474393e-20

R49_104 V49 V104 55423.32319070893
L49_104 V49 V104 1.2968660701455729e-11
C49_104 V49 V104 -1.8945429493456285e-20

R49_105 V49 V105 22946.747868734616
L49_105 V49 V105 -5.014464136747895e-12
C49_105 V49 V105 -1.0608645412620527e-19

R49_106 V49 V106 5484.113662353245
L49_106 V49 V106 3.914242235120251e-12
C49_106 V49 V106 1.97285793311581e-19

R49_107 V49 V107 -691025.9206056959
L49_107 V49 V107 9.600027638829487e-12
C49_107 V49 V107 5.359410783513773e-20

R49_108 V49 V108 -91650.95230036575
L49_108 V49 V108 -1.0127529147481408e-11
C49_108 V49 V108 -1.8823729859272965e-20

R49_109 V49 V109 -24455.016866259033
L49_109 V49 V109 2.123606323712366e-11
C49_109 V49 V109 -2.1363251112250817e-20

R49_110 V49 V110 -9863.783622336527
L49_110 V49 V110 -3.5127225387816173e-12
C49_110 V49 V110 -1.935662334510967e-19

R49_111 V49 V111 -50794.35366828147
L49_111 V49 V111 -1.0461183346252534e-11
C49_111 V49 V111 -6.307565334081154e-20

R49_112 V49 V112 -16104.247636633125
L49_112 V49 V112 8.882514795934286e-12
C49_112 V49 V112 4.7762194906360057e-20

R49_113 V49 V113 29066.273304586102
L49_113 V49 V113 2.329085319053479e-11
C49_113 V49 V113 4.9979847661730977e-20

R49_114 V49 V114 10606.458553642173
L49_114 V49 V114 6.680209202423926e-12
C49_114 V49 V114 1.0339598412410122e-19

R49_115 V49 V115 -17212.65779435968
L49_115 V49 V115 3.6057128439073795e-11
C49_115 V49 V115 2.829977373789121e-20

R49_116 V49 V116 31549.267247296288
L49_116 V49 V116 -1.1829759684461386e-11
C49_116 V49 V116 -2.224116059302667e-20

R49_117 V49 V117 -35528.26164349062
L49_117 V49 V117 -2.4609344341497447e-11
C49_117 V49 V117 -4.454673442432385e-20

R49_118 V49 V118 -129525.60134680365
L49_118 V49 V118 -9.791633798187079e-12
C49_118 V49 V118 -8.862109130753055e-20

R49_119 V49 V119 -29394.35365550544
L49_119 V49 V119 -7.2450373412194395e-12
C49_119 V49 V119 -8.404012116441899e-20

R49_120 V49 V120 -60940.887197217184
L49_120 V49 V120 -2.7536267237279563e-11
C49_120 V49 V120 -8.15501323873271e-21

R49_121 V49 V121 -14344.972209014064
L49_121 V49 V121 1.4869766863354384e-11
C49_121 V49 V121 3.5726259098462665e-20

R49_122 V49 V122 -29841.551058443933
L49_122 V49 V122 4.551340043143809e-11
C49_122 V49 V122 9.873730225077085e-21

R49_123 V49 V123 -85366.39743369975
L49_123 V49 V123 -3.8149014331388876e-11
C49_123 V49 V123 -2.960605037878787e-20

R49_124 V49 V124 -17166.51416026286
L49_124 V49 V124 -2.1931717826625207e-11
C49_124 V49 V124 -1.8251494056984492e-20

R49_125 V49 V125 30337.83213087805
L49_125 V49 V125 -1.7771181456201663e-11
C49_125 V49 V125 -1.2536484448616807e-20

R49_126 V49 V126 8912424.463221997
L49_126 V49 V126 8.589052868387576e-09
C49_126 V49 V126 -9.58529879412292e-22

R49_127 V49 V127 -19409.86494397678
L49_127 V49 V127 3.7909096876785705e-10
C49_127 V49 V127 1.866678548229176e-21

R49_128 V49 V128 -21460.750308502462
L49_128 V49 V128 -4.916044473923862e-11
C49_128 V49 V128 -3.428774183946762e-20

R49_129 V49 V129 -15646.864250320403
L49_129 V49 V129 -2.851919425120435e-11
C49_129 V49 V129 -1.899519050576611e-20

R49_130 V49 V130 -11387.693866007072
L49_130 V49 V130 -3.3003923163026925e-11
C49_130 V49 V130 -2.1920862101523033e-20

R49_131 V49 V131 -30010.680474164692
L49_131 V49 V131 2.7766802690717816e-11
C49_131 V49 V131 1.5009400336164948e-20

R49_132 V49 V132 42910.119208374315
L49_132 V49 V132 -2.2038361167776917e-11
C49_132 V49 V132 -4.1052883019918145e-21

R49_133 V49 V133 12836.46282822927
L49_133 V49 V133 2.8311439260130774e-11
C49_133 V49 V133 3.905611182487028e-20

R49_134 V49 V134 22841.064931880195
L49_134 V49 V134 -6.689314402896984e-11
C49_134 V49 V134 -4.877712973820946e-22

R49_135 V49 V135 35841.8232338387
L49_135 V49 V135 -9.74517438831441e-11
C49_135 V49 V135 -1.2354292472842462e-20

R49_136 V49 V136 -75651.70037917697
L49_136 V49 V136 2.689995930217967e-11
C49_136 V49 V136 1.8273880752814452e-20

R49_137 V49 V137 -13067.834619497582
L49_137 V49 V137 -3.5760998686280924e-11
C49_137 V49 V137 -1.9472275843806162e-20

R49_138 V49 V138 -50793.79583278598
L49_138 V49 V138 -7.107410315480303e-11
C49_138 V49 V138 -1.8625822483942512e-20

R49_139 V49 V139 -28288.31040301415
L49_139 V49 V139 2.935446276867357e-11
C49_139 V49 V139 2.825037376084568e-20

R49_140 V49 V140 11875.14262515825
L49_140 V49 V140 -1.5247714944798903e-10
C49_140 V49 V140 2.143005603185617e-20

R49_141 V49 V141 -22296.359721336266
L49_141 V49 V141 -4.880711221026371e-11
C49_141 V49 V141 -3.576472395152569e-21

R49_142 V49 V142 11073.599652485229
L49_142 V49 V142 -2.0456882431599104e-11
C49_142 V49 V142 -2.3949429986774734e-20

R49_143 V49 V143 -70012.28871563653
L49_143 V49 V143 -6.905157963897631e-11
C49_143 V49 V143 -1.2734380894618415e-20

R49_144 V49 V144 18971.49834266083
L49_144 V49 V144 1.1314762595717057e-08
C49_144 V49 V144 -3.1659848960763546e-20

R50_50 V50 0 100.28606617963277
L50_50 V50 0 6.477599451618449e-14
C50_50 V50 0 1.8672862815816075e-18

R50_51 V50 V51 3126.1659995798364
L50_51 V50 V51 9.46124860861197e-13
C50_51 V50 V51 1.944700356002574e-19

R50_52 V50 V52 -2135.462142293455
L50_52 V50 V52 -6.369010645711284e-13
C50_52 V50 V52 -5.035167082822346e-19

R50_53 V50 V53 -3338.0787704108657
L50_53 V50 V53 -1.2271892459161416e-12
C50_53 V50 V53 -2.5578230761375933e-19

R50_54 V50 V54 -2835.0047128275596
L50_54 V50 V54 -1.7130552215889934e-12
C50_54 V50 V54 -1.4873993027789806e-20

R50_55 V50 V55 2715.212790515406
L50_55 V50 V55 -1.037549032340698e-12
C50_55 V50 V55 1.0256210649900245e-19

R50_56 V50 V56 -3805.427514435849
L50_56 V50 V56 -1.7634083353493206e-12
C50_56 V50 V56 -5.798200756824404e-20

R50_57 V50 V57 -360.2344690187314
L50_57 V50 V57 -3.033955486003932e-13
C50_57 V50 V57 9.686318240012701e-20

R50_58 V50 V58 -1122.500402165471
L50_58 V50 V58 -8.829943242807259e-13
C50_58 V50 V58 1.1698469078413777e-19

R50_59 V50 V59 -409.66381835486425
L50_59 V50 V59 -1.5143429251997058e-12
C50_59 V50 V59 3.358304137291205e-20

R50_60 V50 V60 -4152.923053890629
L50_60 V50 V60 -1.4379827877702523e-12
C50_60 V50 V60 4.086403941040711e-20

R50_61 V50 V61 1122.099881327017
L50_61 V50 V61 5.61451280942801e-12
C50_61 V50 V61 -3.3650703186655925e-19

R50_62 V50 V62 -48431.49975305771
L50_62 V50 V62 -1.4594267325979448e-11
C50_62 V50 V62 -3.3482669676554363e-19

R50_63 V50 V63 -264376.43184726173
L50_63 V50 V63 4.0718814770079724e-11
C50_63 V50 V63 8.224479478558026e-20

R50_64 V50 V64 -2990.618056740266
L50_64 V50 V64 -6.513861281144726e-12
C50_64 V50 V64 -4.894845115512216e-20

R50_65 V50 V65 -701.0776007107977
L50_65 V50 V65 -5.006670064608729e-13
C50_65 V50 V65 -2.0460004236212104e-19

R50_66 V50 V66 -1215.4725713812554
L50_66 V50 V66 -5.501184868004733e-13
C50_66 V50 V66 3.563681952931397e-20

R50_67 V50 V67 -3242.2580480955016
L50_67 V50 V67 -2.2680066773362767e-11
C50_67 V50 V67 8.624381731512515e-20

R50_68 V50 V68 4131.361007209418
L50_68 V50 V68 -5.6979967040208295e-12
C50_68 V50 V68 -5.553964943607597e-20

R50_69 V50 V69 1206.985478284506
L50_69 V50 V69 1.1921556134598219e-12
C50_69 V50 V69 -3.013797127379395e-20

R50_70 V50 V70 -12883.971115125185
L50_70 V50 V70 8.96678739194082e-12
C50_70 V50 V70 2.6911547408630225e-20

R50_71 V50 V71 9467.995364791335
L50_71 V50 V71 -4.3508558428342486e-12
C50_71 V50 V71 -4.44889533587754e-20

R50_72 V50 V72 8739.457282484369
L50_72 V50 V72 1.4740401605146974e-12
C50_72 V50 V72 5.415408161314382e-20

R50_73 V50 V73 14946.731954345092
L50_73 V50 V73 6.482471944731746e-12
C50_73 V50 V73 -3.048333100428631e-20

R50_74 V50 V74 2453.0674628208726
L50_74 V50 V74 1.7665529989724118e-12
C50_74 V50 V74 5.412202774685193e-21

R50_75 V50 V75 -13936.198288013185
L50_75 V50 V75 -2.586733721563855e-12
C50_75 V50 V75 -5.533083993156e-20

R50_76 V50 V76 -4780.342824505421
L50_76 V50 V76 -2.0875080132338905e-12
C50_76 V50 V76 -9.018261009466984e-20

R50_77 V50 V77 -15651.620555789708
L50_77 V50 V77 -3.349566112576793e-12
C50_77 V50 V77 -4.888396349309064e-20

R50_78 V50 V78 -28508.71178035867
L50_78 V50 V78 2.51198497010595e-11
C50_78 V50 V78 1.090606676419104e-19

R50_79 V50 V79 15414.717299545542
L50_79 V50 V79 8.227544771364243e-12
C50_79 V50 V79 -4.848273240552503e-20

R50_80 V50 V80 11581.538517404135
L50_80 V50 V80 6.272597047900132e-12
C50_80 V50 V80 1.0180550651737133e-19

R50_81 V50 V81 65026.11247333953
L50_81 V50 V81 4.101302915823037e-12
C50_81 V50 V81 -1.2769312653461563e-21

R50_82 V50 V82 289799.44779951096
L50_82 V50 V82 -2.8198696135039072e-12
C50_82 V50 V82 -1.2025910040290578e-19

R50_83 V50 V83 167729.93100001448
L50_83 V50 V83 -3.1170946085419955e-12
C50_83 V50 V83 -7.460532517250707e-20

R50_84 V50 V84 -14866.203972251627
L50_84 V50 V84 1.4503837841052444e-11
C50_84 V50 V84 -1.73196818336297e-20

R50_85 V50 V85 66200.92127449602
L50_85 V50 V85 4.392058523766568e-12
C50_85 V50 V85 3.0766828743454784e-20

R50_86 V50 V86 16545.89650705657
L50_86 V50 V86 4.783422119285105e-12
C50_86 V50 V86 5.2296182285038287e-20

R50_87 V50 V87 14574.621848984336
L50_87 V50 V87 5.070272406784745e-12
C50_87 V50 V87 2.835159560860967e-20

R50_88 V50 V88 40358.35422333217
L50_88 V50 V88 1.1468062400148081e-11
C50_88 V50 V88 2.4070361847626496e-20

R50_89 V50 V89 -80650.68780566314
L50_89 V50 V89 -3.5358804879386036e-10
C50_89 V50 V89 3.2493317481511057e-20

R50_90 V50 V90 38258.18015496512
L50_90 V50 V90 1.441850122513754e-09
C50_90 V50 V90 3.530474688605205e-20

R50_91 V50 V91 -16711.065385968894
L50_91 V50 V91 -3.724192970020229e-12
C50_91 V50 V91 -9.202881228557302e-20

R50_92 V50 V92 73499.8321900236
L50_92 V50 V92 -5.500557561582657e-12
C50_92 V50 V92 8.845589829172424e-21

R50_93 V50 V93 7438.544902311317
L50_93 V50 V93 1.1889564919750732e-11
C50_93 V50 V93 3.811113158571104e-20

R50_94 V50 V94 13183.40970108479
L50_94 V50 V94 8.091641587024036e-12
C50_94 V50 V94 2.87739124352283e-20

R50_95 V50 V95 -37819.45186672112
L50_95 V50 V95 -5.6414501008982095e-12
C50_95 V50 V95 -5.0500152800197547e-20

R50_96 V50 V96 -11654.311883887787
L50_96 V50 V96 -6.06134615962184e-12
C50_96 V50 V96 4.296749957439076e-20

R50_97 V50 V97 25141.04145097014
L50_97 V50 V97 5.620476257733258e-12
C50_97 V50 V97 5.750286551951029e-20

R50_98 V50 V98 15002.084308663629
L50_98 V50 V98 -9.306173525084951e-12
C50_98 V50 V98 -1.8431862460929868e-20

R50_99 V50 V99 11932.412570221215
L50_99 V50 V99 3.109423414254236e-11
C50_99 V50 V99 -5.942576881012892e-21

R50_100 V50 V100 -25907.293762633042
L50_100 V50 V100 9.589462625491775e-12
C50_100 V50 V100 1.9297406819912714e-20

R50_101 V50 V101 17254.545834565604
L50_101 V50 V101 -6.601165481665544e-12
C50_101 V50 V101 -1.131117060228913e-20

R50_102 V50 V102 8095.885314518114
L50_102 V50 V102 -8.059651913469775e-12
C50_102 V50 V102 -6.981959084806708e-21

R50_103 V50 V103 45317.052122912566
L50_103 V50 V103 9.57812258612238e-12
C50_103 V50 V103 -1.2051144006250926e-20

R50_104 V50 V104 119623.98899645515
L50_104 V50 V104 -5.540925594520823e-11
C50_104 V50 V104 4.914794900002586e-20

R50_105 V50 V105 -18103.409037382542
L50_105 V50 V105 3.954949391015043e-12
C50_105 V50 V105 7.391761241842765e-20

R50_106 V50 V106 -9750.848381931084
L50_106 V50 V106 -2.2674398100265027e-12
C50_106 V50 V106 -9.167105477111118e-20

R50_107 V50 V107 72633.77862607746
L50_107 V50 V107 -9.316430040576882e-12
C50_107 V50 V107 1.1233556285650267e-20

R50_108 V50 V108 -13430.971411645123
L50_108 V50 V108 7.346433137207075e-12
C50_108 V50 V108 -2.5129807485348525e-20

R50_109 V50 V109 60241.90694348716
L50_109 V50 V109 7.274258557388087e-11
C50_109 V50 V109 2.2534900321375087e-20

R50_110 V50 V110 32274.243588375335
L50_110 V50 V110 3.055127835091826e-12
C50_110 V50 V110 8.592677571108465e-20

R50_111 V50 V111 150824.09804415426
L50_111 V50 V111 4.772817058164219e-12
C50_111 V50 V111 3.144960758015697e-20

R50_112 V50 V112 57553.69206298006
L50_112 V50 V112 -1.1008826484689899e-11
C50_112 V50 V112 7.359726406526463e-21

R50_113 V50 V113 -14096.649576646665
L50_113 V50 V113 -1.8148719546021903e-11
C50_113 V50 V113 -2.2042810586100378e-20

R50_114 V50 V114 -16178.985969764813
L50_114 V50 V114 -5.324234117208215e-12
C50_114 V50 V114 -3.6588180775289624e-20

R50_115 V50 V115 19121.37787716353
L50_115 V50 V115 -3.5086606012684676e-11
C50_115 V50 V115 2.909426471600112e-20

R50_116 V50 V116 -24027.89825223603
L50_116 V50 V116 1.0318533903779771e-11
C50_116 V50 V116 2.8730116952509825e-21

R50_117 V50 V117 617073.8923419992
L50_117 V50 V117 2.470403327361805e-11
C50_117 V50 V117 1.4679691484376124e-20

R50_118 V50 V118 96481.91901967414
L50_118 V50 V118 8.046843229951844e-12
C50_118 V50 V118 4.06729777424592e-20

R50_119 V50 V119 -110351.03348391059
L50_119 V50 V119 4.582492729088922e-12
C50_119 V50 V119 1.602223807634202e-20

R50_120 V50 V120 -33223.46406636245
L50_120 V50 V120 -2.4658293187866096e-11
C50_120 V50 V120 -3.135866964454651e-20

R50_121 V50 V121 -41048.167538997266
L50_121 V50 V121 6.911495433366624e-11
C50_121 V50 V121 -3.8271888843999265e-20

R50_122 V50 V122 -5970.271216972396
L50_122 V50 V122 1.148473135674395e-11
C50_122 V50 V122 1.444305480190857e-20

R50_123 V50 V123 -92288.94431347263
L50_123 V50 V123 1.896791822699674e-11
C50_123 V50 V123 6.896561186910798e-21

R50_124 V50 V124 18982.80270752988
L50_124 V50 V124 2.5859366829340014e-11
C50_124 V50 V124 -3.39605898763492e-20

R50_125 V50 V125 20867.446685615338
L50_125 V50 V125 -3.2361507933184334e-11
C50_125 V50 V125 2.5295468858938756e-20

R50_126 V50 V126 5330.066379186579
L50_126 V50 V126 -2.6587051723731443e-11
C50_126 V50 V126 -2.5228652939915278e-21

R50_127 V50 V127 -13267.230011559517
L50_127 V50 V127 -2.4549001401835127e-11
C50_127 V50 V127 -1.6792987975152357e-20

R50_128 V50 V128 41927.977208471675
L50_128 V50 V128 -1.5496399489811486e-10
C50_128 V50 V128 1.19536813468136e-20

R50_129 V50 V129 58122.506343785106
L50_129 V50 V129 1.8103413808463641e-10
C50_129 V50 V129 -1.9819371442019468e-20

R50_130 V50 V130 13147.707928578226
L50_130 V50 V130 -3.194565058917514e-11
C50_130 V50 V130 -1.4247107435588802e-20

R50_131 V50 V131 13393.591331057125
L50_131 V50 V131 -9.804772841498354e-12
C50_131 V50 V131 -1.43385253735788e-20

R50_132 V50 V132 65099.920615091454
L50_132 V50 V132 9.583860534778004e-11
C50_132 V50 V132 -4.424828682270379e-21

R50_133 V50 V133 -30610.916352356307
L50_133 V50 V133 -9.754826549718887e-12
C50_133 V50 V133 -1.0887603986813765e-21

R50_134 V50 V134 161955.74074412097
L50_134 V50 V134 -7.441176794232861e-11
C50_134 V50 V134 -6.934311970192766e-21

R50_135 V50 V135 -9005.708343331356
L50_135 V50 V135 -1.2133552200597302e-10
C50_135 V50 V135 -7.213338969586563e-21

R50_136 V50 V136 100706.36620156182
L50_136 V50 V136 -2.634327282368432e-11
C50_136 V50 V136 -2.0498798106462042e-20

R50_137 V50 V137 8984.114205170716
L50_137 V50 V137 -1.941823365888404e-11
C50_137 V50 V137 -3.566187512189343e-20

R50_138 V50 V138 5907.721434831797
L50_138 V50 V138 -1.3713009198232915e-11
C50_138 V50 V138 -2.8977547640397176e-20

R50_139 V50 V139 -8789.082383800322
L50_139 V50 V139 -1.5415858259330108e-11
C50_139 V50 V139 2.0602986082635966e-21

R50_140 V50 V140 -25694.796285575703
L50_140 V50 V140 6.670665459470613e-10
C50_140 V50 V140 4.695545710103945e-21

R50_141 V50 V141 11084.529952255756
L50_141 V50 V141 4.838481901198675e-11
C50_141 V50 V141 -5.5483088907444515e-21

R50_142 V50 V142 -14215.198758324714
L50_142 V50 V142 4.499905399588199e-11
C50_142 V50 V142 3.500701363589195e-20

R50_143 V50 V143 23535.042181416575
L50_143 V50 V143 -2.689816499241814e-10
C50_143 V50 V143 -2.2485709435540635e-21

R50_144 V50 V144 -11780.522931118827
L50_144 V50 V144 1.6485517217446845e-11
C50_144 V50 V144 4.046410504230598e-20

R51_51 V51 0 -123.9306803152764
L51_51 V51 0 -8.084701087600171e-14
C51_51 V51 0 -1.885142725903879e-18

R51_52 V51 V52 3932.005712073585
L51_52 V51 V52 7.252124826136894e-13
C51_52 V51 V52 5.522617879867402e-19

R51_53 V51 V53 6583.644978493298
L51_53 V51 V53 2.7624424988686616e-12
C51_53 V51 V53 1.333096691884215e-19

R51_54 V51 V54 2500.7033334927146
L51_54 V51 V54 1.313840623688141e-12
C51_54 V51 V54 2.5065665491246117e-19

R51_55 V51 V55 2489.5122431139503
L51_55 V51 V55 1.0074719964490335e-12
C51_55 V51 V55 2.374396124584255e-19

R51_56 V51 V56 2214.8198508442433
L51_56 V51 V56 5.69896712521667e-12
C51_56 V51 V56 1.1238099727887973e-19

R51_57 V51 V57 396.4512948353232
L51_57 V51 V57 3.190635517492492e-13
C51_57 V51 V57 -8.258144414161319e-20

R51_58 V51 V58 1182.5588871098598
L51_58 V51 V58 4.746163155032963e-13
C51_58 V51 V58 -1.6655781855129818e-19

R51_59 V51 V59 4393.501415328589
L51_59 V51 V59 5.148400119333971e-12
C51_59 V51 V59 -1.324917948115541e-19

R51_60 V51 V60 -6735.681692410882
L51_60 V51 V60 2.8189932177515715e-12
C51_60 V51 V60 -3.988447973870303e-20

R51_61 V51 V61 -2137.516065559868
L51_61 V51 V61 -3.6467677284648965e-12
C51_61 V51 V61 2.9281135493220853e-19

R51_62 V51 V62 -1321.9371820399922
L51_62 V51 V62 -6.187742688443074e-11
C51_62 V51 V62 4.0379592785413147e-19

R51_63 V51 V63 4967.932002846851
L51_63 V51 V63 -7.1650449736810124e-12
C51_63 V51 V63 -2.389086263796552e-19

R51_64 V51 V64 5360.817488670273
L51_64 V51 V64 -6.877163797986363e-11
C51_64 V51 V64 -4.305585940154411e-20

R51_65 V51 V65 882.9880385701492
L51_65 V51 V65 6.398112081317145e-13
C51_65 V51 V65 6.057609279915992e-20

R51_66 V51 V66 871.4534534563456
L51_66 V51 V66 4.3987532421158385e-13
C51_66 V51 V66 2.1423144386040227e-19

R51_67 V51 V67 1010912.6935151784
L51_67 V51 V67 -9.976364011450243e-13
C51_67 V51 V67 -4.948090673685324e-20

R51_68 V51 V68 -9597.338533223452
L51_68 V51 V68 -1.3014645126044336e-11
C51_68 V51 V68 2.174375565956563e-20

R51_69 V51 V69 -4592.6357271517145
L51_69 V51 V69 -1.1823959940134322e-12
C51_69 V51 V69 -8.789782842582433e-20

R51_70 V51 V70 -7315.247952274407
L51_70 V51 V70 3.556686608808139e-12
C51_70 V51 V70 4.302682305012821e-20

R51_71 V51 V71 4104.850346124707
L51_71 V51 V71 7.898701831686521e-13
C51_71 V51 V71 8.845866022447022e-20

R51_72 V51 V72 -2630.174909434555
L51_72 V51 V72 -1.328462808995269e-12
C51_72 V51 V72 -3.058666050731565e-20

R51_73 V51 V73 -6993.339332001888
L51_73 V51 V73 -2.5009054336671373e-12
C51_73 V51 V73 2.6734414597195017e-20

R51_74 V51 V74 -3330.6864262890135
L51_74 V51 V74 -1.6677768824860995e-12
C51_74 V51 V74 -1.3271496876840078e-20

R51_75 V51 V75 3789.191033596694
L51_75 V51 V75 5.164123467221721e-12
C51_75 V51 V75 -6.591112476406718e-21

R51_76 V51 V76 5569.079173271592
L51_76 V51 V76 1.6868331980825647e-12
C51_76 V51 V76 1.508183643240972e-19

R51_77 V51 V77 18144.950707123993
L51_77 V51 V77 3.235559791585191e-12
C51_77 V51 V77 8.297950423658202e-20

R51_78 V51 V78 -34866.85701592242
L51_78 V51 V78 8.295514985205984e-12
C51_78 V51 V78 6.657134356713504e-20

R51_79 V51 V79 -9960.87663377739
L51_79 V51 V79 3.043984085982049e-11
C51_79 V51 V79 1.1014477313878753e-19

R51_80 V51 V80 -21519.39836198165
L51_80 V51 V80 -4.841656534443348e-12
C51_80 V51 V80 -1.0240735790089072e-19

R51_81 V51 V81 -50333.25310056847
L51_81 V51 V81 -8.903207600473766e-12
C51_81 V51 V81 -2.747746413853235e-20

R51_82 V51 V82 -25771.804900395295
L51_82 V51 V82 -3.518620846615527e-12
C51_82 V51 V82 -9.925186079122525e-20

R51_83 V51 V83 21029.52510184127
L51_83 V51 V83 5.171794326417706e-12
C51_83 V51 V83 -6.090394379121451e-20

R51_84 V51 V84 -23379.431257785694
L51_84 V51 V84 -6.824403252033349e-12
C51_84 V51 V84 -2.969300125961012e-21

R51_85 V51 V85 -13623.850438735331
L51_85 V51 V85 -1.7679572137106297e-11
C51_85 V51 V85 1.257531942427025e-20

R51_86 V51 V86 -9999.934960616065
L51_86 V51 V86 -6.097260338789468e-12
C51_86 V51 V86 -1.0730067888545182e-20

R51_87 V51 V87 35366.037279584954
L51_87 V51 V87 9.71896993404081e-12
C51_87 V51 V87 6.387352977174448e-20

R51_88 V51 V88 -132966.97327432074
L51_88 V51 V88 3.780357168874388e-10
C51_88 V51 V88 3.2588690644784847e-23

R51_89 V51 V89 44616.842151448895
L51_89 V51 V89 -9.624195725583666e-12
C51_89 V51 V89 -3.141753276845027e-20

R51_90 V51 V90 23490.881703280364
L51_90 V51 V90 1.4387696994817002e-10
C51_90 V51 V90 -5.00573045488194e-20

R51_91 V51 V91 -80922.6831855992
L51_91 V51 V91 -1.3783261894058128e-11
C51_91 V51 V91 -4.122306278777395e-20

R51_92 V51 V92 -104459.08307978249
L51_92 V51 V92 -5.35428538722364e-11
C51_92 V51 V92 -4.867847230573344e-20

R51_93 V51 V93 -6876.980414638083
L51_93 V51 V93 1.0837869010268189e-08
C51_93 V51 V93 7.705443427824045e-21

R51_94 V51 V94 -12033.67442827881
L51_94 V51 V94 3.046694167893131e-11
C51_94 V51 V94 3.2057546304985503e-20

R51_95 V51 V95 65135.974129846574
L51_95 V51 V95 -3.6354789545073574e-11
C51_95 V51 V95 -2.914116870949947e-20

R51_96 V51 V96 33481.74940694376
L51_96 V51 V96 2.5386044795119208e-11
C51_96 V51 V96 -4.2105334186120616e-20

R51_97 V51 V97 -17806.977014234893
L51_97 V51 V97 -1.49152065333408e-11
C51_97 V51 V97 -2.254890016839284e-20

R51_98 V51 V98 -20922.430673278603
L51_98 V51 V98 -1.68070917758047e-11
C51_98 V51 V98 -4.136655039692641e-20

R51_99 V51 V99 -10537.508523211864
L51_99 V51 V99 1.578731719792429e-11
C51_99 V51 V99 3.1087732481536404e-20

R51_100 V51 V100 37193.15963749452
L51_100 V51 V100 -4.823543225774317e-11
C51_100 V51 V100 8.387019911738935e-21

R51_101 V51 V101 -11573.614434562001
L51_101 V51 V101 -4.1805996852864316e-11
C51_101 V51 V101 -1.8333592038150076e-20

R51_102 V51 V102 -32900.87955774037
L51_102 V51 V102 -9.481138590257747e-12
C51_102 V51 V102 -5.943529295370342e-20

R51_103 V51 V103 -69129.09802817763
L51_103 V51 V103 -2.214621219381799e-11
C51_103 V51 V103 2.0933343213630043e-20

R51_104 V51 V104 -66865.48685712928
L51_104 V51 V104 2.0887650970669274e-11
C51_104 V51 V104 -1.7856433892242098e-20

R51_105 V51 V105 11095.397973329773
L51_105 V51 V105 1.7063656924156357e-11
C51_105 V51 V105 4.505058384530449e-20

R51_106 V51 V106 144663.4271185957
L51_106 V51 V106 -8.629442750704701e-12
C51_106 V51 V106 -9.651170501125513e-20

R51_107 V51 V107 -12772.975622455151
L51_107 V51 V107 -5.345264276116327e-12
C51_107 V51 V107 -1.255759417019807e-19

R51_108 V51 V108 9300.365407854288
L51_108 V51 V108 6.861486784136526e-12
C51_108 V51 V108 9.803733933001072e-20

R51_109 V51 V109 -73116.75904568819
L51_109 V51 V109 1.048786177319222e-11
C51_109 V51 V109 7.525983423989565e-21

R51_110 V51 V110 6736.374037880094
L51_110 V51 V110 7.227390365634788e-12
C51_110 V51 V110 1.031105644359691e-19

R51_111 V51 V111 -32953.79411775152
L51_111 V51 V111 1.1913689058760162e-11
C51_111 V51 V111 5.661471574039348e-20

R51_112 V51 V112 12639.15067614703
L51_112 V51 V112 -9.725791727690904e-12
C51_112 V51 V112 -5.318852014909812e-20

R51_113 V51 V113 10481.495812415373
L51_113 V51 V113 -1.700024515029022e-11
C51_113 V51 V113 -1.8478887357462113e-21

R51_114 V51 V114 79223.1825222976
L51_114 V51 V114 -1.0084500414872799e-11
C51_114 V51 V114 -7.384408990599785e-20

R51_115 V51 V115 308479.76967041724
L51_115 V51 V115 -9.343525028928011e-12
C51_115 V51 V115 -6.02705341017527e-20

R51_116 V51 V116 -41396.22310879863
L51_116 V51 V116 1.165905224702186e-11
C51_116 V51 V116 3.4977437060828216e-20

R51_117 V51 V117 372053.3903429188
L51_117 V51 V117 1.9138759167722888e-11
C51_117 V51 V117 9.091463870415911e-21

R51_118 V51 V118 24456.240171147158
L51_118 V51 V118 9.070565501001248e-12
C51_118 V51 V118 4.745490395490554e-20

R51_119 V51 V119 49225.324120865735
L51_119 V51 V119 9.771231424616639e-12
C51_119 V51 V119 7.551264490044658e-20

R51_120 V51 V120 4637.370621343446
L51_120 V51 V120 -1.9381972459979735e-11
C51_120 V51 V120 4.658954837095854e-20

R51_121 V51 V121 14680.70440776958
L51_121 V51 V121 -2.962071851386588e-11
C51_121 V51 V121 -1.91960537855522e-23

R51_122 V51 V122 2214.772585908828
L51_122 V51 V122 -8.373780068546265e-12
C51_122 V51 V122 9.17390561145171e-21

R51_123 V51 V123 14638.790836091717
L51_123 V51 V123 -6.837651819933125e-09
C51_123 V51 V123 1.703196415124038e-20

R51_124 V51 V124 156699.99984908517
L51_124 V51 V124 1.4981963910130703e-11
C51_124 V51 V124 5.944217668820173e-20

R51_125 V51 V125 -51496.959633289895
L51_125 V51 V125 3.577509341966407e-11
C51_125 V51 V125 5.523244842035738e-21

R51_126 V51 V126 -1833.6257312709654
L51_126 V51 V126 4.824414347813216e-12
C51_126 V51 V126 2.6502407763464545e-20

R51_127 V51 V127 2824.3239971398357
L51_127 V51 V127 -7.948823767348073e-12
C51_127 V51 V127 1.4253924345136126e-20

R51_128 V51 V128 -110157.88599699075
L51_128 V51 V128 -3.105775547114294e-10
C51_128 V51 V128 7.106220816623013e-21

R51_129 V51 V129 8242.995036489876
L51_129 V51 V129 -2.21378305728759e-11
C51_129 V51 V129 1.0009802079272999e-20

R51_130 V51 V130 -8829.502328479553
L51_130 V51 V130 1.0376447579882887e-11
C51_130 V51 V130 2.889867164835114e-20

R51_131 V51 V131 -5556.77451837373
L51_131 V51 V131 2.9248587031790626e-11
C51_131 V51 V131 -3.3221221385319616e-21

R51_132 V51 V132 -10826.73139920494
L51_132 V51 V132 5.72072077146037e-11
C51_132 V51 V132 -1.3457729952480194e-21

R51_133 V51 V133 -38122.54546098446
L51_133 V51 V133 -4.25635701297342e-11
C51_133 V51 V133 -1.3819105141192035e-20

R51_134 V51 V134 226464.54732402114
L51_134 V51 V134 9.263537083915283e-11
C51_134 V51 V134 -2.0453935592160693e-21

R51_135 V51 V135 3655.762096607576
L51_135 V51 V135 -3.045609505263525e-11
C51_135 V51 V135 4.0187927656310725e-20

R51_136 V51 V136 -64921.88699515921
L51_136 V51 V136 4.984796817003669e-11
C51_136 V51 V136 1.6587888033271065e-20

R51_137 V51 V137 -18701.973647717572
L51_137 V51 V137 1.7982031847629126e-11
C51_137 V51 V137 4.8807925505785433e-20

R51_138 V51 V138 -2199.737483027057
L51_138 V51 V138 8.493772794750993e-12
C51_138 V51 V138 7.149049057420806e-21

R51_139 V51 V139 2425.77730982243
L51_139 V51 V139 -6.129781172901213e-12
C51_139 V51 V139 -1.7936266375965796e-20

R51_140 V51 V140 -17166.027684547847
L51_140 V51 V140 2.0898969793433753e-11
C51_140 V51 V140 -1.0537221004561934e-20

R51_141 V51 V141 -8244.296380371115
L51_141 V51 V141 2.2124619402999633e-11
C51_141 V51 V141 1.1233533644778877e-20

R51_142 V51 V142 -21496.153421812043
L51_142 V51 V142 1.8716895996077373e-11
C51_142 V51 V142 6.449483015718191e-21

R51_143 V51 V143 -6976.2794517304665
L51_143 V51 V143 1.0843305644196957e-11
C51_143 V51 V143 2.3049006412515244e-20

R51_144 V51 V144 9081.36719090431
L51_144 V51 V144 -1.1681929172997347e-11
C51_144 V51 V144 -1.839771115991777e-20

R52_52 V52 0 -3348.1812259939456
L52_52 V52 0 3.4356937901469115e-14
C52_52 V52 0 7.989481654969016e-18

R52_53 V52 V53 -4377.9885138426935
L52_53 V52 V53 -5.55832001230086e-13
C52_53 V52 V53 -6.878589916519495e-19

R52_54 V52 V54 16131.261649666129
L52_54 V52 V54 -9.901495490844814e-13
C52_54 V52 V54 -1.6636685691282908e-19

R52_55 V52 V55 -20762.20883909537
L52_55 V52 V55 -6.285758292183138e-13
C52_55 V52 V55 -5.4010417105984e-19

R52_56 V52 V56 -2576.6982805515167
L52_56 V52 V56 -1.139509478076102e-12
C52_56 V52 V56 -5.995646171690174e-19

R52_57 V52 V57 836.3602566634977
L52_57 V52 V57 -1.7833882716909153e-13
C52_57 V52 V57 2.9265355580063076e-19

R52_58 V52 V58 -2068.9787934808046
L52_58 V52 V58 -5.189190575256634e-13
C52_58 V52 V58 1.9396050307606e-19

R52_59 V52 V59 -4837.582977476773
L52_59 V52 V59 -2.500248440125803e-12
C52_59 V52 V59 2.3345508353957586e-19

R52_60 V52 V60 849.7674915003653
L52_60 V52 V60 -8.434543502001501e-13
C52_60 V52 V60 7.677473148599497e-20

R52_61 V52 V61 -1550.4598579058131
L52_61 V52 V61 1.1740601571463542e-10
C52_61 V52 V61 -1.0417833352657934e-18

R52_62 V52 V62 -1785.465361900338
L52_62 V52 V62 9.206131642459382e-12
C52_62 V52 V62 -9.083412236283186e-19

R52_63 V52 V63 -5570.5958808338355
L52_63 V52 V63 -3.102396369631515e-11
C52_63 V52 V63 -1.3925025400929826e-19

R52_64 V52 V64 -6419.734420572516
L52_64 V52 V64 -2.3107305697783857e-12
C52_64 V52 V64 -1.8699961009887396e-19

R52_65 V52 V65 6386.783147678559
L52_65 V52 V65 -2.701410702442377e-13
C52_65 V52 V65 -2.951680608569196e-19

R52_66 V52 V66 -18097.306090451195
L52_66 V52 V66 -2.6607253434139725e-13
C52_66 V52 V66 -3.284722264478924e-19

R52_67 V52 V67 5974.005529918877
L52_67 V52 V67 -1.3378826028125975e-12
C52_67 V52 V67 -1.9850907499844566e-19

R52_68 V52 V68 3302.884664639461
L52_68 V52 V68 -2.3931975445163177e-12
C52_68 V52 V68 -1.4268381279929946e-19

R52_69 V52 V69 18201.534399765387
L52_69 V52 V69 1.0769105535328191e-12
C52_69 V52 V69 1.0389854418362766e-19

R52_70 V52 V70 -28280.36489525674
L52_70 V52 V70 1.5088780220022553e-12
C52_70 V52 V70 -1.1208937820844837e-19

R52_71 V52 V71 -72460.88872282162
L52_71 V52 V71 1.8363984980185297e-12
C52_71 V52 V71 -3.5491941169290245e-20

R52_72 V52 V72 -27704.376398048455
L52_72 V52 V72 8.319698045395644e-13
C52_72 V52 V72 -1.565293975260215e-20

R52_73 V52 V73 17849.269257971737
L52_73 V52 V73 6.860161687341812e-12
C52_73 V52 V73 -1.473746815045006e-19

R52_74 V52 V74 28354.330757384145
L52_74 V52 V74 1.0506821940969423e-12
C52_74 V52 V74 1.6385754337348241e-19

R52_75 V52 V75 300375.0322547944
L52_75 V52 V75 -1.207041158092874e-12
C52_75 V52 V75 -1.2547485288611557e-19

R52_76 V52 V76 -11108.639591093845
L52_76 V52 V76 -8.782108498255595e-13
C52_76 V52 V76 -1.8596998523955826e-19

R52_77 V52 V77 -15967.093599913997
L52_77 V52 V77 -2.1611661327778314e-12
C52_77 V52 V77 -3.559752806569434e-20

R52_78 V52 V78 -11595.735572960539
L52_78 V52 V78 -2.3867364610208298e-12
C52_78 V52 V78 -1.0510962305818067e-19

R52_79 V52 V79 -212966.62973174785
L52_79 V52 V79 3.01071881567866e-12
C52_79 V52 V79 1.8134965892362856e-20

R52_80 V52 V80 46857.1339524004
L52_80 V52 V80 3.628637393505343e-12
C52_80 V52 V80 4.5972173044083604e-20

R52_81 V52 V81 57440.96201059564
L52_81 V52 V81 2.7810879601624375e-12
C52_81 V52 V81 -3.969583023737993e-20

R52_82 V52 V82 47178.25958074541
L52_82 V52 V82 -7.935034165062595e-12
C52_82 V52 V82 9.867460567684576e-20

R52_83 V52 V83 35609.942467691195
L52_83 V52 V83 5.11218111862214e-12
C52_83 V52 V83 5.104677878055533e-20

R52_84 V52 V84 -104333.41738913118
L52_84 V52 V84 5.323414039658358e-12
C52_84 V52 V84 -9.209043458563418e-21

R52_85 V52 V85 -229141.18009254293
L52_85 V52 V85 3.2741971688702842e-12
C52_85 V52 V85 -1.1956477619647893e-20

R52_86 V52 V86 94610.1300016062
L52_86 V52 V86 4.575526370466644e-11
C52_86 V52 V86 -1.3305906677765696e-20

R52_87 V52 V87 -36203.5522970941
L52_87 V52 V87 -4.232408422562362e-11
C52_87 V52 V87 -5.486653615897151e-20

R52_88 V52 V88 -107599.16860376047
L52_88 V52 V88 -1.487550199832055e-11
C52_88 V52 V88 -3.6152480711814475e-20

R52_89 V52 V89 45217.046440870705
L52_89 V52 V89 -6.951623412660032e-11
C52_89 V52 V89 7.409864601554851e-20

R52_90 V52 V90 -180560.12320639138
L52_90 V52 V90 -1.91265932177762e-11
C52_90 V52 V90 -2.4012341784152757e-20

R52_91 V52 V91 50347.95136128677
L52_91 V52 V91 9.333748878368965e-12
C52_91 V52 V91 6.493394816333486e-20

R52_92 V52 V92 32426.338623750114
L52_92 V52 V92 -1.9448559348348723e-11
C52_92 V52 V92 7.401362263387948e-20

R52_93 V52 V93 45448.74521881629
L52_93 V52 V93 1.1803661345328416e-11
C52_93 V52 V93 2.6939725434466822e-20

R52_94 V52 V94 -80427.15605330929
L52_94 V52 V94 -1.6699584527998377e-10
C52_94 V52 V94 -6.597112715421467e-20

R52_95 V52 V95 35477.14938060447
L52_95 V52 V95 2.9901749771459106e-11
C52_95 V52 V95 5.974797354393713e-20

R52_96 V52 V96 37133.34362614053
L52_96 V52 V96 -7.61947830229999e-12
C52_96 V52 V96 8.242824567216154e-20

R52_97 V52 V97 -17432.978935837546
L52_97 V52 V97 7.681641677609617e-11
C52_97 V52 V97 -4.926728273966575e-20

R52_98 V52 V98 -12398.80878613066
L52_98 V52 V98 1.626939169125578e-11
C52_98 V52 V98 3.3878157013003965e-20

R52_99 V52 V99 -47202.60616298894
L52_99 V52 V99 1.8308827110752043e-11
C52_99 V52 V99 -1.731967168162916e-21

R52_100 V52 V100 -55283.912928885
L52_100 V52 V100 2.7089117510760865e-11
C52_100 V52 V100 -2.51262005632383e-20

R52_101 V52 V101 85780.39310055997
L52_101 V52 V101 4.4045415639794136e-11
C52_101 V52 V101 6.397246545851514e-20

R52_102 V52 V102 -20848.139768494562
L52_102 V52 V102 -9.295239562862808e-12
C52_102 V52 V102 -6.41020112899359e-20

R52_103 V52 V103 142292.7080171366
L52_103 V52 V103 5.859521392923104e-12
C52_103 V52 V103 3.7491739947178535e-20

R52_104 V52 V104 22954.41123115479
L52_104 V52 V104 -1.1442586916036189e-11
C52_104 V52 V104 5.079116267803154e-20

R52_105 V52 V105 425491.13503906794
L52_105 V52 V105 2.818667940515545e-11
C52_105 V52 V105 -3.64449065225207e-21

R52_106 V52 V106 11271.374683287833
L52_106 V52 V106 -8.539677493673576e-12
C52_106 V52 V106 4.8531377025473743e-20

R52_107 V52 V107 -17896.099735053223
L52_107 V52 V107 -8.03370291966189e-12
C52_107 V52 V107 -5.70350051542143e-20

R52_108 V52 V108 -15484.243147655478
L52_108 V52 V108 5.5335744925199434e-12
C52_108 V52 V108 5.28297972765333e-20

R52_109 V52 V109 73546.93552845815
L52_109 V52 V109 4.9310281382988207e-11
C52_109 V52 V109 6.94335267068285e-20

R52_110 V52 V110 -86964.74388232027
L52_110 V52 V110 -2.2506510715735525e-11
C52_110 V52 V110 -6.916373959417556e-20

R52_111 V52 V111 -28922.858554931383
L52_111 V52 V111 6.2944715888210115e-12
C52_111 V52 V111 -1.2295272683618137e-21

R52_112 V52 V112 -16045.387252627912
L52_112 V52 V112 -3.8324645972735006e-11
C52_112 V52 V112 4.198702428152296e-21

R52_113 V52 V113 -19920.362547262448
L52_113 V52 V113 8.737194345900261e-11
C52_113 V52 V113 -2.63634412279456e-21

R52_114 V52 V114 35924.70990313574
L52_114 V52 V114 2.9778857679090664e-10
C52_114 V52 V114 6.786013389791501e-20

R52_115 V52 V115 -53264.48537502633
L52_115 V52 V115 -1.0632828353784861e-11
C52_115 V52 V115 -4.111663840982687e-21

R52_116 V52 V116 -75449.34184625388
L52_116 V52 V116 9.538121090198166e-12
C52_116 V52 V116 3.0575557687605296e-20

R52_117 V52 V117 124094.55594712796
L52_117 V52 V117 2.341534906936311e-10
C52_117 V52 V117 2.1556724782102655e-20

R52_118 V52 V118 27008.089187808702
L52_118 V52 V118 -3.907722566923681e-11
C52_118 V52 V118 -9.22092915810042e-21

R52_119 V52 V119 -16065.514995293006
L52_119 V52 V119 1.3597413419732505e-11
C52_119 V52 V119 -6.41856547476576e-20

R52_120 V52 V120 15744.845663932501
L52_120 V52 V120 -7.881158105939494e-12
C52_120 V52 V120 -3.961413853068667e-20

R52_121 V52 V121 -8085.21826974479
L52_121 V52 V121 8.773901528057066e-12
C52_121 V52 V121 -4.886212169538386e-21

R52_122 V52 V122 -10550.483541904388
L52_122 V52 V122 3.7131491202344036e-11
C52_122 V52 V122 3.6338168423290437e-20

R52_123 V52 V123 -234083.86248741808
L52_123 V52 V123 -8.336629158796863e-11
C52_123 V52 V123 -2.3899334986709115e-20

R52_124 V52 V124 -28499.623591545445
L52_124 V52 V124 3.677720002790855e-11
C52_124 V52 V124 -5.598763902814838e-20

R52_125 V52 V125 6639.551647258051
L52_125 V52 V125 -9.465467257289133e-12
C52_125 V52 V125 3.098657707171629e-20

R52_126 V52 V126 315531.70897713886
L52_126 V52 V126 9.211609809808789e-12
C52_126 V52 V126 -1.2540091089266276e-21

R52_127 V52 V127 -367049.40084566514
L52_127 V52 V127 -7.375784148415228e-12
C52_127 V52 V127 -3.0851175925631875e-20

R52_128 V52 V128 -62770.59206938765
L52_128 V52 V128 -3.179298014639753e-11
C52_128 V52 V128 -1.873792891946017e-20

R52_129 V52 V129 -79544.0176005432
L52_129 V52 V129 -1.241551866756666e-11
C52_129 V52 V129 -6.039644977672066e-20

R52_130 V52 V130 -28661.161575366288
L52_130 V52 V130 6.774999578909293e-11
C52_130 V52 V130 6.042695856634111e-22

R52_131 V52 V131 -73900.29911628606
L52_131 V52 V131 -3.3074849901559875e-11
C52_131 V52 V131 -5.859763702373326e-21

R52_132 V52 V132 66216.80318794718
L52_132 V52 V132 3.467860250263416e-11
C52_132 V52 V132 -7.997666749262694e-21

R52_133 V52 V133 21871.577589781
L52_133 V52 V133 -2.7783005567085918e-11
C52_133 V52 V133 1.3023997700992654e-20

R52_134 V52 V134 16301.864504694442
L52_134 V52 V134 -2.8508765478456945e-11
C52_134 V52 V134 -2.2230383966973686e-20

R52_135 V52 V135 77378.13677427183
L52_135 V52 V135 -1.8125033388319187e-11
C52_135 V52 V135 4.541762899774585e-21

R52_136 V52 V136 -287980.9617598492
L52_136 V52 V136 -5.630875463305383e-11
C52_136 V52 V136 -1.1503332698406714e-20

R52_137 V52 V137 23726.85610833504
L52_137 V52 V137 -1.2958188552600182e-11
C52_137 V52 V137 -4.365469991567964e-20

R52_138 V52 V138 81552.80055482521
L52_138 V52 V138 9.406900078334164e-11
C52_138 V52 V138 -8.410393331319065e-20

R52_139 V52 V139 87066.94229263905
L52_139 V52 V139 -6.746039915294451e-12
C52_139 V52 V139 2.59011696544555e-20

R52_140 V52 V140 26774.086027608195
L52_140 V52 V140 5.537108158270973e-11
C52_140 V52 V140 3.69982954510824e-20

R52_141 V52 V141 94531.6238651373
L52_141 V52 V141 4.1255014397088866e-11
C52_141 V52 V141 -1.7596306449624495e-20

R52_142 V52 V142 -60416.52843344326
L52_142 V52 V142 -5.831583235528942e-11
C52_142 V52 V142 1.4388929406681936e-20

R52_143 V52 V143 -28908.598647863015
L52_143 V52 V143 1.5161125429469866e-11
C52_143 V52 V143 7.657806401014813e-22

R52_144 V52 V144 -39214.932784091085
L52_144 V52 V144 3.0216307490194763e-10
C52_144 V52 V144 -2.9756867580189704e-21

R53_53 V53 0 284.83453722908206
L53_53 V53 0 5.664386698038628e-14
C53_53 V53 0 3.678643311036725e-18

R53_54 V53 V54 -3757.6747505780777
L53_54 V53 V54 -1.9736135693178574e-12
C53_54 V53 V54 -1.0534004542024482e-19

R53_55 V53 V55 -35495.38139031781
L53_55 V53 V55 -1.069379129610579e-12
C53_55 V53 V55 -2.4475200959449555e-19

R53_56 V53 V56 -14645.328363274348
L53_56 V53 V56 -1.18355390223792e-12
C53_56 V53 V56 -6.598340098022659e-21

R53_57 V53 V57 -2155.1429466937684
L53_57 V53 V57 -3.0919073843350275e-13
C53_57 V53 V57 2.111214451775731e-19

R53_58 V53 V58 619.9403702170495
L53_58 V53 V58 6.197258774761536e-12
C53_58 V53 V58 3.229921797400745e-20

R53_59 V53 V59 -2965.799822982732
L53_59 V53 V59 -8.012822149705497e-12
C53_59 V53 V59 7.429878593935314e-20

R53_60 V53 V60 -925.9372434191489
L53_60 V53 V60 -3.830932930543872e-12
C53_60 V53 V60 -1.461562642814021e-21

R53_61 V53 V61 -13259.503100942391
L53_61 V53 V61 -2.2704542644622965e-12
C53_61 V53 V61 -6.319197197727741e-19

R53_62 V53 V62 -3696.6764231384122
L53_62 V53 V62 4.64065341062404e-12
C53_62 V53 V62 -3.856297265341744e-19

R53_63 V53 V63 2862.9682656710906
L53_63 V53 V63 3.049307350781425e-12
C53_63 V53 V63 -1.9766779080241408e-19

R53_64 V53 V64 -12317.612325025191
L53_64 V53 V64 -3.1261507802284447e-12
C53_64 V53 V64 -1.3620063379150557e-20

R53_65 V53 V65 -2193.9108372184846
L53_65 V53 V65 -3.8732912424945964e-13
C53_65 V53 V65 -1.8331617979305134e-19

R53_66 V53 V66 -5301.302643730068
L53_66 V53 V66 -3.8134865066466195e-13
C53_66 V53 V66 -1.3587317240772035e-19

R53_67 V53 V67 -2380.6803934344603
L53_67 V53 V67 -1.189108894349351e-12
C53_67 V53 V67 -7.934693363583145e-20

R53_68 V53 V68 -3952.114348000154
L53_68 V53 V68 -1.250291043008495e-11
C53_68 V53 V68 -1.5330471336986734e-20

R53_69 V53 V69 3279.078805493514
L53_69 V53 V69 1.984866698286412e-12
C53_69 V53 V69 9.719555538870223e-21

R53_70 V53 V70 -7303.875088397944
L53_70 V53 V70 2.2735051315837968e-12
C53_70 V53 V70 -1.681857622590403e-19

R53_71 V53 V71 -9390.57163381373
L53_71 V53 V71 3.1172665690836437e-12
C53_71 V53 V71 -5.722732654893083e-20

R53_72 V53 V72 5543.273191035558
L53_72 V53 V72 9.715811615082531e-13
C53_72 V53 V72 -2.133120389820544e-20

R53_73 V53 V73 14096.07200541913
L53_73 V53 V73 4.203067349355057e-12
C53_73 V53 V73 -7.397937272603103e-20

R53_74 V53 V74 4721.713477156388
L53_74 V53 V74 1.4789259532047426e-12
C53_74 V53 V74 6.132223082640596e-20

R53_75 V53 V75 -13119.977348768847
L53_75 V53 V75 -1.7527452795409062e-12
C53_75 V53 V75 8.387602877101665e-21

R53_76 V53 V76 -23466.627752589957
L53_76 V53 V76 -1.0228223867475062e-12
C53_76 V53 V76 -1.94762550582982e-19

R53_77 V53 V77 21924.67150526924
L53_77 V53 V77 -2.356051901333248e-12
C53_77 V53 V77 -6.202083586550873e-20

R53_78 V53 V78 -59507.53130106875
L53_78 V53 V78 -2.798568677143625e-12
C53_78 V53 V78 -8.020518904585039e-20

R53_79 V53 V79 17663.45941744864
L53_79 V53 V79 4.185376524534004e-11
C53_79 V53 V79 -1.811348805665662e-19

R53_80 V53 V80 11842.205739611813
L53_80 V53 V80 2.0803343767744102e-12
C53_80 V53 V80 2.277185767685179e-19

R53_81 V53 V81 1251907.0825089298
L53_81 V53 V81 2.685205990087692e-12
C53_81 V53 V81 5.795710838859762e-20

R53_82 V53 V82 12196.887604661639
L53_82 V53 V82 6.8077824216038675e-12
C53_82 V53 V82 2.190487114484863e-19

R53_83 V53 V83 100779.0898247644
L53_83 V53 V83 2.1735155167660427e-12
C53_83 V53 V83 1.8784601635211012e-19

R53_84 V53 V84 14556.695162529928
L53_84 V53 V84 7.626302803161703e-12
C53_84 V53 V84 -9.835807576695936e-20

R53_85 V53 V85 187177.0011866843
L53_85 V53 V85 1.5297549576812776e-11
C53_85 V53 V85 -1.5938810075982085e-19

R53_86 V53 V86 33290.13669540215
L53_86 V53 V86 -1.4208786979905529e-11
C53_86 V53 V86 -7.384569111832262e-20

R53_87 V53 V87 -14935.928356459524
L53_87 V53 V87 -3.426718482193405e-12
C53_87 V53 V87 -1.8531483238404043e-19

R53_88 V53 V88 -40023.28815289072
L53_88 V53 V88 -1.3892627929322286e-11
C53_88 V53 V88 -8.603646206435577e-21

R53_89 V53 V89 24234.294239446455
L53_89 V53 V89 2.3653512951543352e-11
C53_89 V53 V89 1.4117558389482426e-19

R53_90 V53 V90 36278.546186844935
L53_90 V53 V90 3.610022288467172e-12
C53_90 V53 V90 1.9517646117340189e-19

R53_91 V53 V91 16950.26835541529
L53_91 V53 V91 2.3285793310612465e-12
C53_91 V53 V91 2.1120727102805074e-19

R53_92 V53 V92 21584.169166803542
L53_92 V53 V92 8.408824602514908e-12
C53_92 V53 V92 1.1012773266639698e-19

R53_93 V53 V93 11079.346689802842
L53_93 V53 V93 -3.4749417101851565e-11
C53_93 V53 V93 1.1019628448707855e-20

R53_94 V53 V94 -133255.75683185397
L53_94 V53 V94 -1.3271282054372737e-11
C53_94 V53 V94 -2.728394489660459e-20

R53_95 V53 V95 12549.519147642524
L53_95 V53 V95 5.0347049017879795e-12
C53_95 V53 V95 1.3269581597447028e-19

R53_96 V53 V96 35137.03418602172
L53_96 V53 V96 -4.533114724591026e-11
C53_96 V53 V96 5.684494208406524e-20

R53_97 V53 V97 46008.23614706068
L53_97 V53 V97 6.097469057535887e-12
C53_97 V53 V97 6.807427935779763e-20

R53_98 V53 V98 13729.203392811498
L53_98 V53 V98 3.262862890628836e-12
C53_98 V53 V98 1.4245179231962142e-19

R53_99 V53 V99 -2063621.9578270863
L53_99 V53 V99 -8.425211336535955e-12
C53_99 V53 V99 -3.954742203645889e-20

R53_100 V53 V100 -124773.49210434363
L53_100 V53 V100 4.375185677641661e-11
C53_100 V53 V100 5.011574044969349e-21

R53_101 V53 V101 13475.059959132264
L53_101 V53 V101 7.385213575281631e-12
C53_101 V53 V101 1.4565411662674876e-19

R53_102 V53 V102 5609.180006979854
L53_102 V53 V102 1.6030987158777346e-12
C53_102 V53 V102 4.254282815323307e-19

R53_103 V53 V103 -10040.965066228135
L53_103 V53 V103 -4.280709708118432e-12
C53_103 V53 V103 -2.2470563413588654e-19

R53_104 V53 V104 57074.915759530304
L53_104 V53 V104 -8.961562437466911e-12
C53_104 V53 V104 1.1134780548886097e-20

R53_105 V53 V105 -22532.736915493868
L53_105 V53 V105 -2.998725177707481e-12
C53_105 V53 V105 -1.716330515136867e-19

R53_106 V53 V106 7365.646004783858
L53_106 V53 V106 1.952013764511615e-12
C53_106 V53 V106 3.8292301995619097e-19

R53_107 V53 V107 7908.817974775767
L53_107 V53 V107 1.880427357385677e-12
C53_107 V53 V107 3.593365280467397e-19

R53_108 V53 V108 -9673.914929156317
L53_108 V53 V108 -2.6147846775718246e-12
C53_108 V53 V108 -3.1672830557571997e-19

R53_109 V53 V109 -14735.393672825589
L53_109 V53 V109 -4.701970995817196e-12
C53_109 V53 V109 -1.277770655281622e-19

R53_110 V53 V110 -12834.525200725066
L53_110 V53 V110 -2.554514189001293e-12
C53_110 V53 V110 -2.797553076266619e-19

R53_111 V53 V111 -7784.164414471739
L53_111 V53 V111 -4.122781848990981e-12
C53_111 V53 V111 -1.7497241047165497e-19

R53_112 V53 V112 8699.452794703895
L53_112 V53 V112 1.9487543686337755e-12
C53_112 V53 V112 2.9513253056431947e-19

R53_113 V53 V113 14726.62034613476
L53_113 V53 V113 4.113464212767007e-12
C53_113 V53 V113 1.1643857546207727e-19

R53_114 V53 V114 13614.268492850048
L53_114 V53 V114 3.538878781604974e-12
C53_114 V53 V114 1.739617170541364e-19

R53_115 V53 V115 7560.31910245618
L53_115 V53 V115 3.4161656325820274e-12
C53_115 V53 V115 2.2164462929171703e-19

R53_116 V53 V116 -13538.307077795773
L53_116 V53 V116 -3.657292061225425e-12
C53_116 V53 V116 -1.653912408252176e-19

R53_117 V53 V117 -17167.523870966703
L53_117 V53 V117 -5.715374810292746e-12
C53_117 V53 V117 -1.52862244704295e-19

R53_118 V53 V118 -14695.647806635774
L53_118 V53 V118 -2.8857716620104847e-12
C53_118 V53 V118 -1.5897614832904962e-19

R53_119 V53 V119 -8670.648592340727
L53_119 V53 V119 -3.398024498325537e-12
C53_119 V53 V119 -1.9701076621238582e-19

R53_120 V53 V120 14929.412421771573
L53_120 V53 V120 1.0294237597389984e-11
C53_120 V53 V120 -9.466629507370158e-20

R53_121 V53 V121 -16088.53971707341
L53_121 V53 V121 4.9757193531355325e-12
C53_121 V53 V121 2.2512853648839272e-20

R53_122 V53 V122 51470.514863284836
L53_122 V53 V122 2.2891270098488638e-12
C53_122 V53 V122 2.524246462213519e-20

R53_123 V53 V123 -54625.52506174309
L53_123 V53 V123 2.313811752864358e-11
C53_123 V53 V123 -3.719615852907406e-20

R53_124 V53 V124 -22956.970671429463
L53_124 V53 V124 -1.1628174477814493e-11
C53_124 V53 V124 -6.96878329387588e-20

R53_125 V53 V125 9196.265052276896
L53_125 V53 V125 -9.638961252366321e-12
C53_125 V53 V125 -1.601113541600888e-20

R53_126 V53 V126 -25678.178629465718
L53_126 V53 V126 -2.4125277857317604e-12
C53_126 V53 V126 3.4230626320531835e-20

R53_127 V53 V127 13465.01413751658
L53_127 V53 V127 3.0447043339592435e-12
C53_127 V53 V127 -9.367124774748056e-21

R53_128 V53 V128 80965.16553640208
L53_128 V53 V128 3.71642459815918e-11
C53_128 V53 V128 -1.6789114160160235e-20

R53_129 V53 V129 -137085.7441278667
L53_129 V53 V129 1.3720148247419548e-11
C53_129 V53 V129 -3.5851621611741974e-20

R53_130 V53 V130 -23375.736713879884
L53_130 V53 V130 -3.8128540035702866e-12
C53_130 V53 V130 -1.1544795423897944e-19

R53_131 V53 V131 22638.614469622902
L53_131 V53 V131 -4.04800399077628e-11
C53_131 V53 V131 7.96449967170501e-20

R53_132 V53 V132 -72496.61369454287
L53_132 V53 V132 -1.5610334769450153e-11
C53_132 V53 V132 9.901950633586598e-21

R53_133 V53 V133 20138.372372934067
L53_133 V53 V133 6.191137028633136e-12
C53_133 V53 V133 1.2216505227055414e-19

R53_134 V53 V134 -91911.99960989143
L53_134 V53 V134 -1.775558581841772e-11
C53_134 V53 V134 3.412915677156309e-21

R53_135 V53 V135 84604.01252331487
L53_135 V53 V135 5.272128045745651e-12
C53_135 V53 V135 -4.949204974425689e-20

R53_136 V53 V136 64683.1548150857
L53_136 V53 V136 -5.709777566802895e-11
C53_136 V53 V136 -1.814343957835979e-20

R53_137 V53 V137 28995.610172975983
L53_137 V53 V137 -5.097074376598161e-12
C53_137 V53 V137 -1.0475147190716399e-19

R53_138 V53 V138 -12067.844910603992
L53_138 V53 V138 -2.2626491154960766e-12
C53_138 V53 V138 -6.976838083503665e-20

R53_139 V53 V139 6194.368924659699
L53_139 V53 V139 2.0797822024219936e-12
C53_139 V53 V139 7.428514158514367e-20

R53_140 V53 V140 -173947.45378576676
L53_140 V53 V140 -5.12434381076119e-12
C53_140 V53 V140 -3.2584501131124046e-21

R53_141 V53 V141 -37907.5770266999
L53_141 V53 V141 -8.479107062202711e-12
C53_141 V53 V141 -2.0665439890201633e-20

R53_142 V53 V142 -136545.2381633988
L53_142 V53 V142 -5.496015055769542e-12
C53_142 V53 V142 -1.6620183305920374e-20

R53_143 V53 V143 -29264.900713620867
L53_143 V53 V143 -6.96627888758888e-12
C53_143 V53 V143 -1.2845777358525723e-20

R53_144 V53 V144 -21557.718945738532
L53_144 V53 V144 5.840148213210143e-12
C53_144 V53 V144 2.1132166017456203e-20

R54_54 V54 0 95.78347873057758
L54_54 V54 0 9.493777715496565e-14
C54_54 V54 0 7.10576155686652e-19

R54_55 V54 V55 -2009.1792654171245
L54_55 V54 V55 -1.957327941842859e-12
C54_55 V54 V55 -1.2888641354685628e-19

R54_56 V54 V56 -4702.938905861536
L54_56 V54 V56 -4.007195269655063e-12
C54_56 V54 V56 4.561006801018347e-21

R54_57 V54 V57 -252.8216973199543
L54_57 V54 V57 -4.797657342635619e-13
C54_57 V54 V57 4.540473396656912e-20

R54_58 V54 V58 -1986.0660747929992
L54_58 V54 V58 -8.540458806448287e-13
C54_58 V54 V58 -1.3025200493387918e-21

R54_59 V54 V59 -4107.625405239368
L54_59 V54 V59 -4.454161697134605e-12
C54_59 V54 V59 -7.161421150702869e-21

R54_60 V54 V60 -1086.408351104542
L54_60 V54 V60 -4.212363014929989e-12
C54_60 V54 V60 4.385128038501902e-21

R54_61 V54 V61 935.6853580484959
L54_61 V54 V61 2.083513201533864e-11
C54_61 V54 V61 -1.4416673000242343e-19

R54_62 V54 V62 979.2902019880011
L54_62 V54 V62 2.142243844899646e-11
C54_62 V54 V62 -1.1384643018917218e-19

R54_63 V54 V63 3920.013692665237
L54_63 V54 V63 -2.406091017418069e-11
C54_63 V54 V63 2.0453133945613352e-20

R54_64 V54 V64 -20881.228776436914
L54_64 V54 V64 -1.0621593816214663e-11
C54_64 V54 V64 6.086985156664019e-21

R54_65 V54 V65 -597.3855073882985
L54_65 V54 V65 -8.864613398581222e-13
C54_65 V54 V65 -1.4187862396128467e-20

R54_66 V54 V66 -652.3340849614168
L54_66 V54 V66 -6.613143376564865e-13
C54_66 V54 V66 -7.900504776035598e-20

R54_67 V54 V67 -2790.8271139822255
L54_67 V54 V67 -5.7928442929084804e-11
C54_67 V54 V67 -2.477992013155715e-22

R54_68 V54 V68 -6161.346707540352
L54_68 V54 V68 -1.3692871569066634e-11
C54_68 V54 V68 8.645120464934654e-21

R54_69 V54 V69 3080.85792703654
L54_69 V54 V69 4.019392526725432e-12
C54_69 V54 V69 2.731035062997503e-20

R54_70 V54 V70 3581.70846136417
L54_70 V54 V70 3.5532459347109397e-11
C54_70 V54 V70 -7.44560208759742e-20

R54_71 V54 V71 141206.46697009975
L54_71 V54 V71 -1.514300825029421e-11
C54_71 V54 V71 -1.084119451004224e-20

R54_72 V54 V72 2041.4454976199042
L54_72 V54 V72 2.902582085221116e-12
C54_72 V54 V72 -2.759806978545506e-20

R54_73 V54 V73 11981.526697485066
L54_73 V54 V73 -8.211807990695096e-11
C54_73 V54 V73 -3.58267735066324e-20

R54_74 V54 V74 2990.2425307694707
L54_74 V54 V74 4.19557574287918e-12
C54_74 V54 V74 1.6635895187657083e-20

R54_75 V54 V75 -3468.8205457181607
L54_75 V54 V75 -5.373509298115568e-12
C54_75 V54 V75 3.616165798040617e-20

R54_76 V54 V76 -3601.521130422825
L54_76 V54 V76 -2.0540950130240163e-12
C54_76 V54 V76 -6.769361129403286e-20

R54_77 V54 V77 -12391.501227315031
L54_77 V54 V77 -5.272550307488674e-12
C54_77 V54 V77 -1.9058601476176334e-20

R54_78 V54 V78 -41723.61667399625
L54_78 V54 V78 -3.197984502454684e-12
C54_78 V54 V78 -8.333700886291921e-20

R54_79 V54 V79 8234.046598650652
L54_79 V54 V79 1.144274355592611e-10
C54_79 V54 V79 -2.0899307679056974e-20

R54_80 V54 V80 9179.761068197511
L54_80 V54 V80 5.299805942920009e-12
C54_80 V54 V80 6.005150857266221e-20

R54_81 V54 V81 31898.88090290843
L54_81 V54 V81 1.2722268664989665e-11
C54_81 V54 V81 -1.0239842949111448e-20

R54_82 V54 V82 15314.754743149218
L54_82 V54 V82 2.1836763483282956e-12
C54_82 V54 V82 1.9129363376794495e-19

R54_83 V54 V83 29623.931987347147
L54_83 V54 V83 3.014907790313574e-12
C54_83 V54 V83 1.5007663675237184e-19

R54_84 V54 V84 40517.852519447464
L54_84 V54 V84 -2.2772828683656835e-08
C54_84 V54 V84 -2.12914848240211e-20

R54_85 V54 V85 11235.400574047739
L54_85 V54 V85 -9.929069392168407e-12
C54_85 V54 V85 -6.593565544356339e-20

R54_86 V54 V86 21667.166746872248
L54_86 V54 V86 -5.684472554554393e-12
C54_86 V54 V86 -4.5221121976317575e-20

R54_87 V54 V87 -19828.861957712736
L54_87 V54 V87 -3.698798827336503e-12
C54_87 V54 V87 -9.771103993430429e-20

R54_88 V54 V88 -155483.51941586673
L54_88 V54 V88 -1.6454013653356018e-11
C54_88 V54 V88 -1.593327680426822e-20

R54_89 V54 V89 -51195.006735345094
L54_89 V54 V89 4.898894024510236e-12
C54_89 V54 V89 9.132903682329895e-20

R54_90 V54 V90 88182.71234932046
L54_90 V54 V90 2.1709617967075476e-11
C54_90 V54 V90 3.1951295860235024e-20

R54_91 V54 V91 13809.019443863548
L54_91 V54 V91 2.230615935329852e-12
C54_91 V54 V91 1.6210149917220662e-19

R54_92 V54 V92 31895.927964946928
L54_92 V54 V92 6.489455229903141e-12
C54_92 V54 V92 9.079758176118863e-20

R54_93 V54 V93 4262.072049640313
L54_93 V54 V93 -2.4444032682972345e-11
C54_93 V54 V93 3.366494224066475e-21

R54_94 V54 V94 25013.864082691893
L54_94 V54 V94 -6.5782361870781895e-12
C54_94 V54 V94 -7.075701092606656e-20

R54_95 V54 V95 24925.926405146307
L54_95 V54 V95 4.469388778067984e-12
C54_95 V54 V95 1.0344721325427755e-19

R54_96 V54 V96 -28595.706975926212
L54_96 V54 V96 5.469395734092512e-09
C54_96 V54 V96 4.775567211637637e-20

R54_97 V54 V97 9575.091191568736
L54_97 V54 V97 -2.333153750157523e-11
C54_97 V54 V97 -2.925885826655714e-20

R54_98 V54 V98 6061.194215136845
L54_98 V54 V98 3.6205267046038924e-12
C54_98 V54 V98 9.035126324487053e-20

R54_99 V54 V99 27580.198986641437
L54_99 V54 V99 -2.601019407366634e-11
C54_99 V54 V99 -2.3863207864826853e-20

R54_100 V54 V100 -28667.16497371943
L54_100 V54 V100 -2.818059855907005e-11
C54_100 V54 V100 -2.559886941297163e-20

R54_101 V54 V101 8198.407794626315
L54_101 V54 V101 3.811461911877852e-12
C54_101 V54 V101 1.0682148076153893e-19

R54_102 V54 V102 8146.266205043544
L54_102 V54 V102 3.441551678761545e-12
C54_102 V54 V102 1.3332921494454576e-19

R54_103 V54 V103 18916.349111833773
L54_103 V54 V103 2.279185012156479e-11
C54_103 V54 V103 -7.039628072488943e-21

R54_104 V54 V104 -143907.54488836322
L54_104 V54 V104 -9.949106807694048e-12
C54_104 V54 V104 5.8973338797379715e-21

R54_105 V54 V105 -6968.984450381396
L54_105 V54 V105 -3.374344047285107e-12
C54_105 V54 V105 -1.2860670202698883e-19

R54_106 V54 V106 -30367.235349448136
L54_106 V54 V106 2.5262705986514466e-12
C54_106 V54 V106 1.99324016138381e-19

R54_107 V54 V107 20104.10810463581
L54_107 V54 V107 5.398264315493578e-12
C54_107 V54 V107 9.752583135428853e-20

R54_108 V54 V108 -21126.091969526
L54_108 V54 V108 -5.0450770563034584e-12
C54_108 V54 V108 -1.1499337125367416e-19

R54_109 V54 V109 267534.1174890564
L54_109 V54 V109 -1.084747298781425e-11
C54_109 V54 V109 -2.435459342518918e-20

R54_110 V54 V110 -17406.853160460352
L54_110 V54 V110 -2.4095503591551738e-12
C54_110 V54 V110 -1.8958951247663054e-19

R54_111 V54 V111 -11860.844560091256
L54_111 V54 V111 -9.073827372688333e-12
C54_111 V54 V111 -8.293158804334621e-20

R54_112 V54 V112 36200.877560773144
L54_112 V54 V112 3.0744902859660585e-12
C54_112 V54 V112 1.1903260417006007e-19

R54_113 V54 V113 -22656.32742271073
L54_113 V54 V113 6.1737839088034666e-12
C54_113 V54 V113 3.9257569657476965e-20

R54_114 V54 V114 10724.775106826793
L54_114 V54 V114 4.154931962359341e-12
C54_114 V54 V114 1.1933577524591094e-19

R54_115 V54 V115 12423.15905581549
L54_115 V54 V115 1.5762157386952095e-11
C54_115 V54 V115 4.2466650996972536e-20

R54_116 V54 V116 -76580.07029215671
L54_116 V54 V116 -7.698541822709137e-12
C54_116 V54 V116 -5.480582668073535e-20

R54_117 V54 V117 12214.11740914855
L54_117 V54 V117 -7.775885367851421e-12
C54_117 V54 V117 -4.3696503398536984e-20

R54_118 V54 V118 -8645.619169958343
L54_118 V54 V118 -4.11346048750992e-12
C54_118 V54 V118 -8.102327493052592e-20

R54_119 V54 V119 -5775.925699151919
L54_119 V54 V119 -4.637988845193232e-12
C54_119 V54 V119 -1.205494325325887e-19

R54_120 V54 V120 5942.494770344291
L54_120 V54 V120 -1.3637359023448955e-11
C54_120 V54 V120 -4.3725047043698556e-20

R54_121 V54 V121 -13537.509202185987
L54_121 V54 V121 5.653242429122016e-12
C54_121 V54 V121 2.5703448386140964e-20

R54_122 V54 V122 -62694.78446233502
L54_122 V54 V122 6.137180557414033e-12
C54_122 V54 V122 7.542903642135942e-23

R54_123 V54 V123 15757.09561751893
L54_123 V54 V123 -3.34569491601208e-11
C54_123 V54 V123 -3.82319849014902e-20

R54_124 V54 V124 46431.71811499648
L54_124 V54 V124 -1.756804758464945e-11
C54_124 V54 V124 -4.7791888685256163e-20

R54_125 V54 V125 5582.714249507536
L54_125 V54 V125 -6.313122513930744e-12
C54_125 V54 V125 -2.301479604855265e-21

R54_126 V54 V126 -28954.811155411917
L54_126 V54 V126 -1.2807883042102483e-11
C54_126 V54 V126 1.4894666054697056e-20

R54_127 V54 V127 8572.117606566539
L54_127 V54 V127 1.7934110211042965e-11
C54_127 V54 V127 -1.4556160904226588e-20

R54_128 V54 V128 37007.3815553381
L54_128 V54 V128 4.6585515391100694e-11
C54_128 V54 V128 -1.3101008380467938e-20

R54_129 V54 V129 8711.916199694548
L54_129 V54 V129 -6.299081011815348e-11
C54_129 V54 V129 -3.5633680892784885e-20

R54_130 V54 V130 -19336.908475326178
L54_130 V54 V130 -1.1497679231292354e-11
C54_130 V54 V130 -4.136932602238464e-20

R54_131 V54 V131 -64420.0074046072
L54_131 V54 V131 4.4901042481922936e-11
C54_131 V54 V131 3.395513721702965e-20

R54_132 V54 V132 -33250.18559608068
L54_132 V54 V132 -2.907664623544817e-10
C54_132 V54 V132 1.6706936455597187e-21

R54_133 V54 V133 -104713.83076404834
L54_133 V54 V133 8.062386696966241e-12
C54_133 V54 V133 6.515983446422195e-20

R54_134 V54 V134 -7941.311465062939
L54_134 V54 V134 -2.292366021820302e-11
C54_134 V54 V134 3.7497891472229736e-21

R54_135 V54 V135 27492.566880611328
L54_135 V54 V135 3.552866263445442e-11
C54_135 V54 V135 -1.4962725487531676e-20

R54_136 V54 V136 64674.08114668019
L54_136 V54 V136 -3.1972065134166065e-10
C54_136 V54 V136 -2.255031837198279e-22

R54_137 V54 V137 6821.05721266413
L54_137 V54 V137 -6.507956242796444e-12
C54_137 V54 V137 -5.083479281191273e-20

R54_138 V54 V138 -12110.66827265261
L54_138 V54 V138 -7.527397269270063e-12
C54_138 V54 V138 -3.941584726746403e-20

R54_139 V54 V139 4789.299384627147
L54_139 V54 V139 1.0186346453491205e-11
C54_139 V54 V139 1.8106997191538256e-20

R54_140 V54 V140 -7410.925431177244
L54_140 V54 V140 -1.4383049465151271e-11
C54_140 V54 V140 -3.980357702232409e-21

R54_141 V54 V141 15894.209868814041
L54_141 V54 V141 -2.0488975921421236e-11
C54_141 V54 V141 -1.0436833871030593e-20

R54_142 V54 V142 -5653.0129258744
L54_142 V54 V142 -7.846642439672383e-12
C54_142 V54 V142 -5.078049125800029e-20

R54_143 V54 V143 -14906.259179066772
L54_143 V54 V143 4.1933502233975077e-11
C54_143 V54 V143 1.2480168605491618e-20

R54_144 V54 V144 -15811.089360653736
L54_144 V54 V144 1.8465338857537785e-11
C54_144 V54 V144 -9.349084668117447e-22

R55_55 V55 0 84.37650775902459
L55_55 V55 0 5.768588032455053e-14
C55_55 V55 0 2.922366384660206e-18

R55_56 V55 V56 -2377.379133347873
L55_56 V55 V56 -1.7341150485396747e-12
C55_56 V55 V56 -2.570192970876531e-19

R55_57 V55 V57 -220.81905733923762
L55_57 V55 V57 -2.6357778914401885e-13
C55_57 V55 V57 1.1599813189494346e-19

R55_58 V55 V58 -597.5059619084766
L55_58 V55 V58 -1.1018629722828747e-12
C55_58 V55 V58 2.6003990377582247e-20

R55_59 V55 V59 853.5993765228659
L55_59 V55 V59 -3.220013216215501e-12
C55_59 V55 V59 2.2543943070390043e-20

R55_60 V55 V60 -2210.450485837651
L55_60 V55 V60 -1.5033727925306817e-12
C55_60 V55 V60 3.75566059067387e-21

R55_61 V55 V61 1005.3975814981125
L55_61 V55 V61 5.0490916462709894e-12
C55_61 V55 V61 -3.7545273309442706e-19

R55_62 V55 V62 573.114075683768
L55_62 V55 V62 9.554717793121494e-12
C55_62 V55 V62 -3.128981853079594e-19

R55_63 V55 V63 -46604.623419784206
L55_63 V55 V63 -1.767065777984653e-11
C55_63 V55 V63 -4.3638176079248363e-20

R55_64 V55 V64 27227.161263991507
L55_64 V55 V64 -1.4149065436135861e-11
C55_64 V55 V64 -1.0126833949207655e-19

R55_65 V55 V65 -549.3275531241671
L55_65 V55 V65 -5.534944996701415e-13
C55_65 V55 V65 -4.728336702221348e-20

R55_66 V55 V66 -473.0801888949298
L55_66 V55 V66 -4.986653919354105e-13
C55_66 V55 V66 -1.9992090833750877e-19

R55_67 V55 V67 -15318.003244879186
L55_67 V55 V67 -2.9717076307554568e-12
C55_67 V55 V67 -1.4096231844057376e-19

R55_68 V55 V68 -7804.6762817814
L55_68 V55 V68 -2.7611200171582614e-12
C55_68 V55 V68 -9.525213535934121e-21

R55_69 V55 V69 11114.983571861592
L55_69 V55 V69 4.8513839060675666e-12
C55_69 V55 V69 1.1177748182956702e-19

R55_70 V55 V70 2268.8339491902484
L55_70 V55 V70 4.377885822315145e-12
C55_70 V55 V70 -1.2890568058577299e-19

R55_71 V55 V71 -6067.169417437576
L55_71 V55 V71 -5.040695661764465e-12
C55_71 V55 V71 -6.335376033525817e-20

R55_72 V55 V72 1567.046710901544
L55_72 V55 V72 1.5295005799949683e-12
C55_72 V55 V72 -3.1985765009438455e-20

R55_73 V55 V73 8006.988340326901
L55_73 V55 V73 -3.8681052420890203e-11
C55_73 V55 V73 -3.961877261871602e-20

R55_74 V55 V74 2798.983893368335
L55_74 V55 V74 3.6431196172752875e-12
C55_74 V55 V74 9.311160996086803e-20

R55_75 V55 V75 -2757.213103702109
L55_75 V55 V75 -2.1055402975688747e-12
C55_75 V55 V75 2.1140943060919557e-20

R55_76 V55 V76 -2674.4990034562306
L55_76 V55 V76 -2.1277623144811217e-12
C55_76 V55 V76 -8.308902665534652e-20

R55_77 V55 V77 -6969.027637078285
L55_77 V55 V77 -3.4265808640557848e-12
C55_77 V55 V77 -2.980715297036816e-20

R55_78 V55 V78 1352583.4373028988
L55_78 V55 V78 -3.125400545075368e-12
C55_78 V55 V78 -1.5757759862495648e-19

R55_79 V55 V79 9790.950952607878
L55_79 V55 V79 1.524769260204944e-11
C55_79 V55 V79 -2.968442778351719e-20

R55_80 V55 V80 9791.247315070668
L55_80 V55 V80 8.065598849253966e-12
C55_80 V55 V80 5.945253084429301e-20

R55_81 V55 V81 17321.469034167203
L55_81 V55 V81 3.2638591147432e-12
C55_81 V55 V81 4.434660593541777e-20

R55_82 V55 V82 11834.470269915557
L55_82 V55 V82 4.9722266189744095e-12
C55_82 V55 V82 2.901803771898862e-19

R55_83 V55 V83 82223.47977302235
L55_83 V55 V83 1.91981251458531e-11
C55_83 V55 V83 2.1308774642710577e-19

R55_84 V55 V84 56835.090735698344
L55_84 V55 V84 1.1642454622959509e-11
C55_84 V55 V84 -3.2103940449527146e-21

R55_85 V55 V85 9404.65084235113
L55_85 V55 V85 1.1620675782411576e-11
C55_85 V55 V85 -6.716737983866919e-20

R55_86 V55 V86 11584.153273492206
L55_86 V55 V86 -1.5853860792629018e-11
C55_86 V55 V86 -7.789789075553962e-20

R55_87 V55 V87 -14200.719711257152
L55_87 V55 V87 -1.1588670725037701e-11
C55_87 V55 V87 -1.0854691673184118e-19

R55_88 V55 V88 -129597.35751429132
L55_88 V55 V88 2.4421092554470046e-11
C55_88 V55 V88 -2.2294355717175107e-20

R55_89 V55 V89 -35643.56630402254
L55_89 V55 V89 1.1811917147967466e-11
C55_89 V55 V89 9.436004136620564e-20

R55_90 V55 V90 -140749.42624777145
L55_90 V55 V90 3.3230822671562685e-11
C55_90 V55 V90 4.313602377283362e-20

R55_91 V55 V91 10046.11718690877
L55_91 V55 V91 3.4779149649406732e-12
C55_91 V55 V91 2.94017910408184e-19

R55_92 V55 V92 96243.16025172328
L55_92 V55 V92 -1.2457064046956642e-11
C55_92 V55 V92 9.977965456179356e-20

R55_93 V55 V93 4250.491060702151
L55_93 V55 V93 4.330136891088957e-11
C55_93 V55 V93 -5.4733064484352264e-21

R55_94 V55 V94 18287.225059832814
L55_94 V55 V94 -5.7082114762288284e-11
C55_94 V55 V94 -9.449909171073107e-20

R55_95 V55 V95 48776.02791262685
L55_95 V55 V95 9.707432876351007e-12
C55_95 V55 V95 1.5479091913383777e-19

R55_96 V55 V96 -24612.268950663823
L55_96 V55 V96 -5.298741644942828e-12
C55_96 V55 V96 5.809420503611979e-21

R55_97 V55 V97 6045.616230969463
L55_97 V55 V97 2.427330506833278e-11
C55_97 V55 V97 -5.3239550412106745e-20

R55_98 V55 V98 4765.600413836766
L55_98 V55 V98 2.044664015236041e-11
C55_98 V55 V98 1.1027618654858974e-19

R55_99 V55 V99 21192.559044979116
L55_99 V55 V99 1.7718526190799743e-10
C55_99 V55 V99 -1.703472648480964e-20

R55_100 V55 V100 -50787.43074449441
L55_100 V55 V100 1.2159676063665796e-11
C55_100 V55 V100 -7.257923320297237e-21

R55_101 V55 V101 7136.739429760413
L55_101 V55 V101 -7.317720487891394e-11
C55_101 V55 V101 9.079894270492773e-20

R55_102 V55 V102 12035.5994220391
L55_102 V55 V102 1.5520300813114484e-11
C55_102 V55 V102 1.4234086163942154e-19

R55_103 V55 V103 11422.787823258832
L55_103 V55 V103 9.345880937408035e-12
C55_103 V55 V103 7.069958578034051e-21

R55_104 V55 V104 -51859.43699882634
L55_104 V55 V104 -8.19846181922935e-12
C55_104 V55 V104 -2.801261104179915e-20

R55_105 V55 V105 -5402.204812114527
L55_105 V55 V105 -3.8409535289142685e-11
C55_105 V55 V105 -1.4601466990053252e-19

R55_106 V55 V106 -21488.243833694458
L55_106 V55 V106 1.1664870947331717e-10
C55_106 V55 V106 2.5654092925652034e-19

R55_107 V55 V107 11861.00412792416
L55_107 V55 V107 3.171661378861176e-11
C55_107 V55 V107 1.0093420243762647e-19

R55_108 V55 V108 -26533.30096223029
L55_108 V55 V108 2.209221313657921e-11
C55_108 V55 V108 -8.05405339831356e-20

R55_109 V55 V109 44629.83325357502
L55_109 V55 V109 -1.0819455512406596e-11
C55_109 V55 V109 -4.293698733625459e-20

R55_110 V55 V110 -6472.9247787800705
L55_110 V55 V110 -1.0100173733913922e-11
C55_110 V55 V110 -2.5571099332289336e-19

R55_111 V55 V111 -28448.139035401287
L55_111 V55 V111 2.132091695530105e-11
C55_111 V55 V111 -7.825256883699454e-20

R55_112 V55 V112 121393.96109102269
L55_112 V55 V112 6.715105920585138e-11
C55_112 V55 V112 1.1304623800791683e-19

R55_113 V55 V113 -14515.644892417087
L55_113 V55 V113 1.4868742796649082e-11
C55_113 V55 V113 5.565713810603738e-20

R55_114 V55 V114 6754.269297393503
L55_114 V55 V114 1.133664347810066e-09
C55_114 V55 V114 1.160130090740545e-19

R55_115 V55 V115 26742.66206056805
L55_115 V55 V115 3.8211793877532005e-11
C55_115 V55 V115 7.818035723272173e-20

R55_116 V55 V116 34405.66451456041
L55_116 V55 V116 2.7874767804768056e-10
C55_116 V55 V116 -7.730139335157875e-20

R55_117 V55 V117 9907.21423401656
L55_117 V55 V117 -1.6359221944118798e-11
C55_117 V55 V117 -6.760392019772036e-20

R55_118 V55 V118 -5775.462787857803
L55_118 V55 V118 -1.2454284619434907e-11
C55_118 V55 V118 -1.2021581250781102e-19

R55_119 V55 V119 -5678.1395426173685
L55_119 V55 V119 -7.578157321488846e-11
C55_119 V55 V119 -1.5297363492119225e-19

R55_120 V55 V120 15858.099563318321
L55_120 V55 V120 1.471130396984691e-10
C55_120 V55 V120 -3.3416915598168096e-20

R55_121 V55 V121 -46520.93657868699
L55_121 V55 V121 1.286298421531232e-11
C55_121 V55 V121 4.5328344798862776e-20

R55_122 V55 V122 -10962.073083275975
L55_122 V55 V122 1.4286683291134545e-11
C55_122 V55 V122 4.947250530605187e-21

R55_123 V55 V123 13940.50776764505
L55_123 V55 V123 -3.544483001368659e-11
C55_123 V55 V123 -6.397654798351478e-20

R55_124 V55 V124 26645.250458064467
L55_124 V55 V124 -2.6612571331336452e-11
C55_124 V55 V124 -5.263055988482441e-20

R55_125 V55 V125 9998.638597601537
L55_125 V55 V125 -4.0499947174770995e-11
C55_125 V55 V125 -5.341469436882611e-21

R55_126 V55 V126 8735.929126603778
L55_126 V55 V126 -2.3347954035256286e-11
C55_126 V55 V126 1.8121827756094976e-20

R55_127 V55 V127 -78789.82104321901
L55_127 V55 V127 -4.636524759118026e-10
C55_127 V55 V127 -3.20901044331936e-21

R55_128 V55 V128 -334558.00469940616
L55_128 V55 V128 3.93181011133197e-10
C55_128 V55 V128 -1.5933203578774177e-20

R55_129 V55 V129 11774.00757733774
L55_129 V55 V129 -6.862241845059833e-11
C55_129 V55 V129 -3.2614137938316827e-20

R55_130 V55 V130 -15930.127851656242
L55_130 V55 V130 -1.4663998638463862e-11
C55_130 V55 V130 -2.8930431778372273e-20

R55_131 V55 V131 -441894.2391299435
L55_131 V55 V131 -1.5063730753171224e-11
C55_131 V55 V131 1.751925259935755e-20

R55_132 V55 V132 -568590.3705389492
L55_132 V55 V132 4.9649648770146504e-11
C55_132 V55 V132 1.0353545992815652e-20

R55_133 V55 V133 -60452.319748572685
L55_133 V55 V133 3.247111504769869e-11
C55_133 V55 V133 9.815750063360407e-20

R55_134 V55 V134 -5961.976361068045
L55_134 V55 V134 -3.397181480589782e-11
C55_134 V55 V134 4.67907459747641e-21

R55_135 V55 V135 -36275.30830452433
L55_135 V55 V135 5.7233601445187207e-11
C55_135 V55 V135 -1.267708797348608e-20

R55_136 V55 V136 136840.25372133186
L55_136 V55 V136 4.539180549938419e-11
C55_136 V55 V136 2.439306145095275e-21

R55_137 V55 V137 9734.767939285583
L55_137 V55 V137 -1.9996700353493874e-11
C55_137 V55 V137 -4.335234363340688e-20

R55_138 V55 V138 -305250.7042089579
L55_138 V55 V138 -8.046193976535265e-12
C55_138 V55 V138 -4.837935067235964e-20

R55_139 V55 V139 17221.682817140372
L55_139 V55 V139 4.0929816762539813e-10
C55_139 V55 V139 1.1838303480372558e-20

R55_140 V55 V140 -6437.777634307009
L55_140 V55 V140 3.2084884430757286e-11
C55_140 V55 V140 7.587473967130076e-21

R55_141 V55 V141 9900.323418846338
L55_141 V55 V141 -4.096550475040744e-11
C55_141 V55 V141 -1.1148222607938313e-20

R55_142 V55 V142 -6488.194402844679
L55_142 V55 V142 -1.0386853907321281e-11
C55_142 V55 V142 -5.107232746793442e-20

R55_143 V55 V143 -34262.473142415045
L55_143 V55 V143 -2.529658010633166e-11
C55_143 V55 V143 -1.622385431616527e-20

R55_144 V55 V144 -21281.880836986053
L55_144 V55 V144 4.22389990628664e-11
C55_144 V55 V144 1.4522933826587694e-20

R56_56 V56 0 359.19931797950545
L56_56 V56 0 6.693575731120499e-14
C56_56 V56 0 4.020231606984418e-18

R56_57 V56 V57 -446.3518930691619
L56_57 V56 V57 -3.771536528858759e-13
C56_57 V56 V57 8.894831844458423e-20

R56_58 V56 V58 1509.4935928071372
L56_58 V56 V58 4.898071507887931e-12
C56_58 V56 V58 -4.085689686515741e-21

R56_59 V56 V59 -8815.077876874175
L56_59 V56 V59 -4.8062866444344e-12
C56_59 V56 V59 2.3656540433520236e-20

R56_60 V56 V60 503.4182310520048
L56_60 V56 V60 -7.438028954828541e-13
C56_60 V56 V60 1.9997295840600024e-20

R56_61 V56 V61 3925.172377915876
L56_61 V56 V61 1.0946666032514909e-11
C56_61 V56 V61 -3.646214083001214e-19

R56_62 V56 V62 1102.0985030340057
L56_62 V56 V62 4.082631136646415e-11
C56_62 V56 V62 -1.774544694781489e-19

R56_63 V56 V63 2506.4571806315453
L56_63 V56 V63 -3.82012569869389e-11
C56_63 V56 V63 -2.3626119274855885e-19

R56_64 V56 V64 -2229.149199338243
L56_64 V56 V64 -1.3617934275051465e-12
C56_64 V56 V64 -5.29656782801986e-19

R56_65 V56 V65 -1125.2694829292998
L56_65 V56 V65 -9.000327283505048e-13
C56_65 V56 V65 9.548647468752163e-21

R56_66 V56 V66 -1056.191960016245
L56_66 V56 V66 -7.750438729834389e-13
C56_66 V56 V66 -2.788081939993603e-19

R56_67 V56 V67 -2608.5680087699197
L56_67 V56 V67 -1.3458086012186563e-12
C56_67 V56 V67 -1.6853648953314536e-19

R56_68 V56 V68 1580.6782676199357
L56_68 V56 V68 -3.4307341056588963e-12
C56_68 V56 V68 -1.4114214584292578e-19

R56_69 V56 V69 -10246.614564788188
L56_69 V56 V69 7.765746881949471e-12
C56_69 V56 V69 5.08151208482752e-20

R56_70 V56 V70 5175.365216127146
L56_70 V56 V70 -2.0554060922308975e-11
C56_70 V56 V70 -2.1092068312723864e-19

R56_71 V56 V71 -5343.856408967254
L56_71 V56 V71 2.0214038347064847e-11
C56_71 V56 V71 -4.633753380212908e-20

R56_72 V56 V72 3679.9415396556115
L56_72 V56 V72 9.671330999371955e-12
C56_72 V56 V72 -6.938933565774263e-20

R56_73 V56 V73 3158.4812821995315
L56_73 V56 V73 -1.8911097727330936e-11
C56_73 V56 V73 -1.0205775154006316e-19

R56_74 V56 V74 3785.7514506767607
L56_74 V56 V74 5.204084896661946e-12
C56_74 V56 V74 4.040423572965176e-20

R56_75 V56 V75 -3493.5779379254404
L56_75 V56 V75 -5.376517015829065e-12
C56_75 V56 V75 4.817324765634596e-20

R56_76 V56 V76 -4782.227908436312
L56_76 V56 V76 -1.553987394376849e-12
C56_76 V56 V76 -1.9349856080440535e-19

R56_77 V56 V77 -24350.146035890877
L56_77 V56 V77 8.406963203176805e-12
C56_77 V56 V77 1.1505837197871321e-19

R56_78 V56 V78 129968.19134090625
L56_78 V56 V78 -2.9611715992195423e-12
C56_78 V56 V78 -1.2127725614995015e-19

R56_79 V56 V79 12475.224825329506
L56_79 V56 V79 -4.4515502266212284e-12
C56_79 V56 V79 -1.7092549740450382e-19

R56_80 V56 V80 9661.981328682346
L56_80 V56 V80 2.049842178173393e-12
C56_80 V56 V80 2.7435024024917007e-19

R56_81 V56 V81 -27427.127370222377
L56_81 V56 V81 -2.5902814648177554e-12
C56_81 V56 V81 -2.5872270885039475e-19

R56_82 V56 V82 10893.982591781765
L56_82 V56 V82 2.496021057998909e-12
C56_82 V56 V82 2.4345032637700855e-19

R56_83 V56 V83 56007.59900460511
L56_83 V56 V83 1.902484492606252e-12
C56_83 V56 V83 3.1498802608732237e-19

R56_84 V56 V84 20896.903862346313
L56_84 V56 V84 -1.0376473036119877e-11
C56_84 V56 V84 -4.9852849063449474e-20

R56_85 V56 V85 15159.01462301317
L56_85 V56 V85 -3.98775854612102e-12
C56_85 V56 V85 -2.0496552286208898e-19

R56_86 V56 V86 8340.503473525108
L56_86 V56 V86 -9.548003949674878e-12
C56_86 V56 V86 -9.597210972372763e-20

R56_87 V56 V87 -9942.8098772638
L56_87 V56 V87 -2.479358722353557e-12
C56_87 V56 V87 -2.1126624794400695e-19

R56_88 V56 V88 -15037.02418784518
L56_88 V56 V88 -7.514819070905885e-12
C56_88 V56 V88 -6.26567220984942e-20

R56_89 V56 V89 -83838.32421064498
L56_89 V56 V89 4.899574944144144e-12
C56_89 V56 V89 1.3111610041031638e-19

R56_90 V56 V90 28290.437831725423
L56_90 V56 V90 3.9939270971194365e-12
C56_90 V56 V90 1.5524940005276023e-19

R56_91 V56 V91 17013.221159107026
L56_91 V56 V91 3.449436942474114e-12
C56_91 V56 V91 1.6081644548860554e-19

R56_92 V56 V92 8541.397422294987
L56_92 V56 V92 1.850957316283648e-12
C56_92 V56 V92 3.321143153901288e-19

R56_93 V56 V93 8258.012891701508
L56_93 V56 V93 -9.615747304657583e-12
C56_93 V56 V93 -5.4053049995243297e-20

R56_94 V56 V94 -30277.173748833684
L56_94 V56 V94 -4.585283557225923e-12
C56_94 V56 V94 -1.1923583947343205e-19

R56_95 V56 V95 27110.271702279068
L56_95 V56 V95 5.440984671465517e-12
C56_95 V56 V95 1.255913645140136e-19

R56_96 V56 V96 22458.209341698646
L56_96 V56 V96 2.1451402212925123e-12
C56_96 V56 V96 3.0962857087581597e-19

R56_97 V56 V97 9943.33643356154
L56_97 V56 V97 -2.5229637619659237e-11
C56_97 V56 V97 -3.744375717308623e-20

R56_98 V56 V98 5078.8007704955035
L56_98 V56 V98 2.6376051182078456e-12
C56_98 V56 V98 2.2243143607507394e-19

R56_99 V56 V99 -90570.68340124981
L56_99 V56 V99 -7.266724284338677e-12
C56_99 V56 V99 -5.805270288173488e-20

R56_100 V56 V100 -12627.605343612186
L56_100 V56 V100 -7.638555465845257e-12
C56_100 V56 V100 -7.195624586681058e-20

R56_101 V56 V101 9703.655892654575
L56_101 V56 V101 3.4586124063463067e-12
C56_101 V56 V101 1.8173920525528913e-19

R56_102 V56 V102 5461.198284891534
L56_102 V56 V102 1.7511595973743061e-12
C56_102 V56 V102 4.02450392989445e-19

R56_103 V56 V103 -136579.12534498103
L56_103 V56 V103 -4.046488073006246e-12
C56_103 V56 V103 -2.0194533051970363e-19

R56_104 V56 V104 15993.155381072473
L56_104 V56 V104 4.689429264663371e-12
C56_104 V56 V104 1.597306821589053e-19

R56_105 V56 V105 -5108.541155793863
L56_105 V56 V105 -2.2362434547138415e-12
C56_105 V56 V105 -2.621085480309794e-19

R56_106 V56 V106 20445.861735721865
L56_106 V56 V106 1.6288363048199326e-12
C56_106 V56 V106 4.246755303192375e-19

R56_107 V56 V107 7824.768352423236
L56_107 V56 V107 2.0783615781775987e-12
C56_107 V56 V107 3.402293470019847e-19

R56_108 V56 V108 -8536.90821757713
L56_108 V56 V108 -1.941822829422576e-12
C56_108 V56 V108 -3.461476058045002e-19

R56_109 V56 V109 12013.164394117593
L56_109 V56 V109 -9.676875739053339e-11
C56_109 V56 V109 -2.4381696682845362e-20

R56_110 V56 V110 -13863.654858425665
L56_110 V56 V110 -2.1367862770137313e-12
C56_110 V56 V110 -3.2655917683453773e-19

R56_111 V56 V111 -8302.461433408376
L56_111 V56 V111 -3.043152172787745e-12
C56_111 V56 V111 -2.1317373465000372e-19

R56_112 V56 V112 6460.212564097721
L56_112 V56 V112 2.1449833095401498e-12
C56_112 V56 V112 2.841641117284422e-19

R56_113 V56 V113 -46539.293495252525
L56_113 V56 V113 4.790405219004355e-12
C56_113 V56 V113 1.3058668612076285e-19

R56_114 V56 V114 8401.633249553855
L56_114 V56 V114 3.64231097048863e-12
C56_114 V56 V114 1.8567462063409618e-19

R56_115 V56 V115 7403.689910149855
L56_115 V56 V115 3.946954177087699e-12
C56_115 V56 V115 1.925829721282886e-19

R56_116 V56 V116 -11678.086272930237
L56_116 V56 V116 -2.7000442385251182e-12
C56_116 V56 V116 -2.2388786655486847e-19

R56_117 V56 V117 18457.62506939989
L56_117 V56 V117 -6.179390314189999e-12
C56_117 V56 V117 -1.4909154233428683e-19

R56_118 V56 V118 -9054.5213797713
L56_118 V56 V118 -3.8849871729467095e-12
C56_118 V56 V118 -1.5269528971806136e-19

R56_119 V56 V119 -5479.460411618363
L56_119 V56 V119 -2.471807829573221e-12
C56_119 V56 V119 -2.421006248111251e-19

R56_120 V56 V120 8709.799628952009
L56_120 V56 V120 6.531313797325648e-11
C56_120 V56 V120 -9.697940238179383e-20

R56_121 V56 V121 29438.01081429526
L56_121 V56 V121 1.1090505791086942e-11
C56_121 V56 V121 2.1811542067597454e-20

R56_122 V56 V122 6055.321777738567
L56_122 V56 V122 4.175333612203001e-12
C56_122 V56 V122 4.489066084065888e-21

R56_123 V56 V123 12246.454163352026
L56_123 V56 V123 -4.905537726313466e-11
C56_123 V56 V123 -3.36018415536341e-20

R56_124 V56 V124 -37732.02170914889
L56_124 V56 V124 -5.8557533388457125e-12
C56_124 V56 V124 -9.010358886298595e-20

R56_125 V56 V125 13638.270255838344
L56_125 V56 V125 -1.1070567189375201e-11
C56_125 V56 V125 -5.347030735996334e-20

R56_126 V56 V126 -5594.332048357196
L56_126 V56 V126 -3.83458158425789e-12
C56_126 V56 V126 3.9506224000439324e-20

R56_127 V56 V127 5863.989104334844
L56_127 V56 V127 4.117662193367421e-12
C56_127 V56 V127 9.346408798985173e-21

R56_128 V56 V128 28400.437556074605
L56_128 V56 V128 1.2171855537817263e-09
C56_128 V56 V128 -1.2776994336390327e-20

R56_129 V56 V129 8433.701226502628
L56_129 V56 V129 3.2125239326113825e-11
C56_129 V56 V129 -1.4242360218630124e-20

R56_130 V56 V130 -10197.783447555496
L56_130 V56 V130 -5.513884517096627e-12
C56_130 V56 V130 -1.0343041671438414e-19

R56_131 V56 V131 -32236.859002667738
L56_131 V56 V131 1.803272541832511e-11
C56_131 V56 V131 8.098410968000825e-20

R56_132 V56 V132 -17293.15198096535
L56_132 V56 V132 -7.034367966974546e-12
C56_132 V56 V132 -5.1561816281618655e-20

R56_133 V56 V133 -98618.13982474536
L56_133 V56 V133 5.248674660770862e-12
C56_133 V56 V133 1.3423889042391335e-19

R56_134 V56 V134 -8641.687717745179
L56_134 V56 V134 -1.8671455874868598e-11
C56_134 V56 V134 1.2391143043948826e-21

R56_135 V56 V135 12822.480065480622
L56_135 V56 V135 7.851722001344624e-12
C56_135 V56 V135 -3.4342231949560434e-20

R56_136 V56 V136 -1757686.5233880193
L56_136 V56 V136 -4.719729899532577e-10
C56_136 V56 V136 -4.477709316057538e-21

R56_137 V56 V137 23637.497733356642
L56_137 V56 V137 -9.375924970221987e-12
C56_137 V56 V137 -5.0251938737647836e-20

R56_138 V56 V138 -4173.982662300232
L56_138 V56 V138 -3.750545312352263e-12
C56_138 V56 V138 -2.880106025695738e-20

R56_139 V56 V139 3399.9501079742445
L56_139 V56 V139 2.8674254888620626e-12
C56_139 V56 V139 4.811042806739308e-20

R56_140 V56 V140 -7196.244009141108
L56_140 V56 V140 -5.4136989399331595e-12
C56_140 V56 V140 -4.88777946724397e-20

R56_141 V56 V141 164067.46067702599
L56_141 V56 V141 -2.150220658427034e-11
C56_141 V56 V141 -2.1716833492576428e-21

R56_142 V56 V142 -5100.05872535269
L56_142 V56 V142 -7.1462525009132615e-12
C56_142 V56 V142 -3.958190173411672e-20

R56_143 V56 V143 -10218.652704642982
L56_143 V56 V143 -8.747219928324402e-12
C56_143 V56 V143 -7.179371401807938e-21

R56_144 V56 V144 -29648.96466148539
L56_144 V56 V144 8.299956830972281e-12
C56_144 V56 V144 4.2794368732459e-20

R57_57 V57 0 9.516562700760124
L57_57 V57 0 1.3309425986698781e-14
C57_57 V57 0 -1.7907296079547088e-18

R57_58 V57 V58 -95.8387766602777
L57_58 V57 V58 -2.4565623558953695e-13
C57_58 V57 V58 -2.4205435028087396e-20

R57_59 V57 V59 -471.6896853347919
L57_59 V57 V59 -3.3450722961639258e-12
C57_59 V57 V59 -3.148808963955398e-20

R57_60 V57 V60 -157.92209111862053
L57_60 V57 V60 -3.6804757725411225e-13
C57_60 V57 V60 -5.302031847462442e-21

R57_61 V57 V61 84.3876425220889
L57_61 V57 V61 9.498728150938697e-13
C57_61 V57 V61 2.9568631287968036e-19

R57_62 V57 V62 85.10791056270307
L57_62 V57 V62 7.510415514883948e-13
C57_62 V57 V62 1.902971962902535e-19

R57_63 V57 V63 757.7010494864179
L57_63 V57 V63 -1.2876988720449847e-12
C57_63 V57 V63 4.49852148678277e-20

R57_64 V57 V64 -2223.2323820350293
L57_64 V57 V64 -1.893077919915612e-12
C57_64 V57 V64 5.423704298288585e-20

R57_65 V57 V65 -59.59650862201645
L57_65 V57 V65 -1.3811047739022668e-13
C57_65 V57 V65 8.632128171265225e-20

R57_66 V57 V66 -67.00131680824968
L57_66 V57 V66 -1.70641277874381e-13
C57_66 V57 V66 1.346176063621652e-19

R57_67 V57 V67 -300.1012330487437
L57_67 V57 V67 -6.83705450409881e-13
C57_67 V57 V67 3.9631065410830776e-20

R57_68 V57 V68 -799.2852275860897
L57_68 V57 V68 -7.988003015626948e-13
C57_68 V57 V68 1.3767017382510453e-20

R57_69 V57 V69 568.8986142485022
L57_69 V57 V69 8.54924758822264e-13
C57_69 V57 V69 -2.6247462181651043e-20

R57_70 V57 V70 260.0700876552409
L57_70 V57 V70 -8.348357850054648e-12
C57_70 V57 V70 7.332829783365287e-20

R57_71 V57 V71 727.1795231192275
L57_71 V57 V71 -4.990941295427126e-12
C57_71 V57 V71 1.471672651649579e-20

R57_72 V57 V72 228.82828523755234
L57_72 V57 V72 1.1758090838124948e-12
C57_72 V57 V72 -1.2782562682695353e-20

R57_73 V57 V73 5484.262089565461
L57_73 V57 V73 -1.0486441699094738e-12
C57_73 V57 V73 2.93129655357315e-20

R57_74 V57 V74 422.33611689177695
L57_74 V57 V74 7.601183164136025e-13
C57_74 V57 V74 -4.5380538269200964e-20

R57_75 V57 V75 -339.18495876782646
L57_75 V57 V75 -8.759745377501267e-13
C57_75 V57 V75 3.801675157402884e-21

R57_76 V57 V76 -361.34132011647574
L57_76 V57 V76 -6.228675000427544e-13
C57_76 V57 V76 1.32638930474784e-19

R57_77 V57 V77 -1017.6113833251817
L57_77 V57 V77 -1.8671269641862127e-12
C57_77 V57 V77 2.1507488036677066e-20

R57_78 V57 V78 -109801.79329262707
L57_78 V57 V78 -3.4074618487184068e-12
C57_78 V57 V78 6.498189599274467e-20

R57_79 V57 V79 1256.7317246131545
L57_79 V57 V79 1.0223149220859115e-11
C57_79 V57 V79 6.700757423744932e-20

R57_80 V57 V80 1053.7702907543173
L57_80 V57 V80 3.0144528884514273e-12
C57_80 V57 V80 -1.435411887286867e-19

R57_81 V57 V81 2079.9426883985357
L57_81 V57 V81 -1.730378372312614e-11
C57_81 V57 V81 2.3463346667131686e-20

R57_82 V57 V82 -35664.088102705
L57_82 V57 V82 5.176876324351199e-12
C57_82 V57 V82 -1.5305232643286625e-19

R57_83 V57 V83 3856.1642953661412
L57_83 V57 V83 -3.22895503968071e-12
C57_83 V57 V83 -1.3751518792704457e-19

R57_84 V57 V84 -15717.023108436444
L57_84 V57 V84 -2.770019230069749e-12
C57_84 V57 V84 3.753887531361257e-20

R57_85 V57 V85 1063.0613160798405
L57_85 V57 V85 -4.1443122865205316e-12
C57_85 V57 V85 9.107265824765124e-20

R57_86 V57 V86 3579.5789683102403
L57_86 V57 V86 -8.618651711080301e-12
C57_86 V57 V86 5.412113230163003e-20

R57_87 V57 V87 -7432.537946937924
L57_87 V57 V87 -1.7150741209267286e-10
C57_87 V57 V87 1.260916610164826e-19

R57_88 V57 V88 6418.520963235742
L57_88 V57 V88 9.327759519516452e-12
C57_88 V57 V88 2.7688091337699984e-20

R57_89 V57 V89 -1560.4318919068978
L57_89 V57 V89 4.041273311055331e-12
C57_89 V57 V89 -9.385206552528349e-20

R57_90 V57 V90 8709.412706535988
L57_90 V57 V90 -1.516356415670537e-11
C57_90 V57 V90 -7.914678439910429e-20

R57_91 V57 V91 5117.237892841619
L57_91 V57 V91 -5.0085330879663045e-12
C57_91 V57 V91 -1.412688457930363e-19

R57_92 V57 V92 -9609.107603379865
L57_92 V57 V92 -1.1301612235271034e-11
C57_92 V57 V92 -1.1496833161265582e-19

R57_93 V57 V93 454.18467472908475
L57_93 V57 V93 7.22075291677627e-12
C57_93 V57 V93 4.341448725421583e-21

R57_94 V57 V94 1130.246010339969
L57_94 V57 V94 1.9246985192813648e-11
C57_94 V57 V94 4.9007559496324996e-20

R57_95 V57 V95 -27775.441370078534
L57_95 V57 V95 -1.5405409601540657e-11
C57_95 V57 V95 -8.363353407273829e-20

R57_96 V57 V96 -1657.5757884516247
L57_96 V57 V96 2.0835225146882774e-10
C57_96 V57 V96 -7.969390639271028e-20

R57_97 V57 V97 932.9680368690756
L57_97 V57 V97 -2.7354095293958202e-11
C57_97 V57 V97 -8.005666762508384e-21

R57_98 V57 V98 764.7727464339972
L57_98 V57 V98 -1.413655875097242e-11
C57_98 V57 V98 -1.0117640220401656e-19

R57_99 V57 V99 1511.0156036840092
L57_99 V57 V99 3.1342110052081225e-11
C57_99 V57 V99 2.2388139247178623e-20

R57_100 V57 V100 -3456.2010837284856
L57_100 V57 V100 8.326300257371981e-11
C57_100 V57 V100 2.2371262963663374e-20

R57_101 V57 V101 1225.063089512965
L57_101 V57 V101 1.436410881245353e-11
C57_101 V57 V101 -1.0390820084455823e-19

R57_102 V57 V102 1437.9227365698011
L57_102 V57 V102 -5.288758416834243e-12
C57_102 V57 V102 -2.0266698406500884e-19

R57_103 V57 V103 1889.534522229932
L57_103 V57 V103 7.346486473627279e-12
C57_103 V57 V103 9.381790949354347e-20

R57_104 V57 V104 -4553.440023829693
L57_104 V57 V104 2.687240910298535e-11
C57_104 V57 V104 -2.7705699326729655e-20

R57_105 V57 V105 -962.0042072421404
L57_105 V57 V105 6.559994845952727e-12
C57_105 V57 V105 1.1994581242721346e-19

R57_106 V57 V106 -846.8471238361577
L57_106 V57 V106 -4.507734958071031e-12
C57_106 V57 V106 -2.3515126479965798e-19

R57_107 V57 V107 3517.2997374661104
L57_107 V57 V107 -4.999268853103041e-12
C57_107 V57 V107 -1.6102172081478262e-19

R57_108 V57 V108 -13210.510551300613
L57_108 V57 V108 8.874368262857995e-12
C57_108 V57 V108 1.8572528036918103e-19

R57_109 V57 V109 6067.633538817988
L57_109 V57 V109 1.835601161097787e-11
C57_109 V57 V109 3.931473412651674e-20

R57_110 V57 V110 -7755.431563853621
L57_110 V57 V110 1.1417954098145441e-11
C57_110 V57 V110 1.8970471877347172e-19

R57_111 V57 V111 -2908.7452049341964
L57_111 V57 V111 9.637690712802817e-12
C57_111 V57 V111 9.853719214764307e-20

R57_112 V57 V112 -2842.9719183553384
L57_112 V57 V112 -5.709034842203646e-12
C57_112 V57 V112 -1.6049910175345942e-19

R57_113 V57 V113 -1565.640888729304
L57_113 V57 V113 -1.163592110580024e-11
C57_113 V57 V113 -6.093662853693876e-20

R57_114 V57 V114 7287.77589153946
L57_114 V57 V114 -1.2976621022645288e-11
C57_114 V57 V114 -1.1147936592952906e-19

R57_115 V57 V115 2278.5286799332425
L57_115 V57 V115 -6.879716278319758e-12
C57_115 V57 V115 -9.457421757459454e-20

R57_116 V57 V116 5233.983614390936
L57_116 V57 V116 6.955425987305699e-12
C57_116 V57 V116 1.129018900058397e-19

R57_117 V57 V117 1082.6682480989268
L57_117 V57 V117 1.4284845955841479e-11
C57_117 V57 V117 7.727154869202798e-20

R57_118 V57 V118 -1278.690250474565
L57_118 V57 V118 7.0502470654764455e-12
C57_118 V57 V118 1.0153780377274572e-19

R57_119 V57 V119 -1066.6459551574676
L57_119 V57 V119 6.510795632560252e-12
C57_119 V57 V119 1.4172671028406534e-19

R57_120 V57 V120 880.7367598451264
L57_120 V57 V120 -1.6255678626607412e-11
C57_120 V57 V120 5.3471044162889886e-20

R57_121 V57 V121 -1527.2819880840475
L57_121 V57 V121 -1.885103195952885e-11
C57_121 V57 V121 -1.1228197883867471e-20

R57_122 V57 V122 -1001.317868235516
L57_122 V57 V122 -7.688315715016065e-12
C57_122 V57 V122 -7.500785164528686e-21

R57_123 V57 V123 2985.9524344853085
L57_123 V57 V123 1.0945297039662313e-10
C57_123 V57 V123 2.3854562437698682e-20

R57_124 V57 V124 6590.4375245462425
L57_124 V57 V124 2.5033002075374595e-11
C57_124 V57 V124 4.516062775748101e-20

R57_125 V57 V125 711.1609255057407
L57_125 V57 V125 6.701017279217525e-11
C57_125 V57 V125 2.963130052312436e-20

R57_126 V57 V126 1359.9232754739794
L57_126 V57 V126 6.324201083366459e-12
C57_126 V57 V126 -1.5097691955011623e-20

R57_127 V57 V127 2727.0274811224645
L57_127 V57 V127 -6.995739258376924e-12
C57_127 V57 V127 4.987965080393728e-21

R57_128 V57 V128 1962.0649350935846
L57_128 V57 V128 -5.885806115168781e-11
C57_128 V57 V128 4.050625085736161e-21

R57_129 V57 V129 1508.4975945740584
L57_129 V57 V129 -1.722637905031359e-11
C57_129 V57 V129 8.206447246161057e-21

R57_130 V57 V130 3556.6231995632097
L57_130 V57 V130 1.7681138241785554e-11
C57_130 V57 V130 5.820039858502649e-20

R57_131 V57 V131 2801.372586345078
L57_131 V57 V131 -1.4167315173872174e-10
C57_131 V57 V131 -3.57583541550923e-20

R57_132 V57 V132 -9465.063583587975
L57_132 V57 V132 4.62360115722167e-11
C57_132 V57 V132 -1.720866951611798e-21

R57_133 V57 V133 -3506.025224275086
L57_133 V57 V133 -1.971516015326934e-11
C57_133 V57 V133 -7.433554984335136e-20

R57_134 V57 V134 -877.3489677545556
L57_134 V57 V134 2.2762252306019916e-10
C57_134 V57 V134 1.1503482910155709e-20

R57_135 V57 V135 -5230.687614988897
L57_135 V57 V135 -1.4180371606957176e-11
C57_135 V57 V135 1.9831899533350472e-20

R57_136 V57 V136 3632.907504072729
L57_136 V57 V136 -1.8245644146949226e-09
C57_136 V57 V136 9.343284738497765e-21

R57_137 V57 V137 689.3121205919167
L57_137 V57 V137 3.064772627340114e-11
C57_137 V57 V137 4.951355373433443e-20

R57_138 V57 V138 2059.2912047076984
L57_138 V57 V138 5.8190113937680886e-12
C57_138 V57 V138 3.046753018378072e-20

R57_139 V57 V139 1085.9740386503963
L57_139 V57 V139 -5.2653466553086526e-12
C57_139 V57 V139 -2.6989901058696127e-20

R57_140 V57 V140 -999.7901154649644
L57_140 V57 V140 1.18426669157371e-11
C57_140 V57 V140 1.302718511522906e-20

R57_141 V57 V141 1488.369574739889
L57_141 V57 V141 2.1526367874474033e-11
C57_141 V57 V141 1.339964891832837e-20

R57_142 V57 V142 -864.6664641628765
L57_142 V57 V142 9.491909711936455e-12
C57_142 V57 V142 9.611590202700623e-21

R57_143 V57 V143 -6109.779801605075
L57_143 V57 V143 1.3233259705346028e-11
C57_143 V57 V143 1.5515369559972357e-20

R57_144 V57 V144 -1261.5987252071097
L57_144 V57 V144 -3.652425499943917e-11
C57_144 V57 V144 -5.589315022514266e-21

R58_58 V58 0 34.98858332253161
L58_58 V58 0 5.250188643418587e-14
C58_58 V58 0 -3.265408575965038e-19

R58_59 V58 V59 6622.78763941663
L58_59 V58 V59 -5.5349927641251486e-12
C58_59 V58 V59 -7.20505443584491e-20

R58_60 V58 V60 -2433.614512537819
L58_60 V58 V60 -1.0209716796397239e-10
C58_60 V58 V60 -1.9810258293202765e-20

R58_61 V58 V61 277.4090686022621
L58_61 V58 V61 1.8032765550053046e-12
C58_61 V58 V61 7.954560653848541e-20

R58_62 V58 V62 261.41333252331935
L58_62 V58 V62 3.375460322504951e-12
C58_62 V58 V62 1.8790829978857508e-19

R58_63 V58 V63 -639.8623861636614
L58_63 V58 V63 -1.0934068397740256e-12
C58_63 V58 V63 -2.1409618002386427e-19

R58_64 V58 V64 4682.904566025398
L58_64 V58 V64 3.0423285466666634e-11
C58_64 V58 V64 -4.8599938949464176e-20

R58_65 V58 V65 -226.42271845941536
L58_65 V58 V65 -5.29734832368889e-13
C58_65 V58 V65 5.053551744049151e-20

R58_66 V58 V66 -164.30931550091898
L58_66 V58 V66 -4.267040151710453e-13
C58_66 V58 V66 7.292571559387833e-20

R58_67 V58 V67 437.7533741122281
L58_67 V58 V67 1.6013059677929818e-12
C58_67 V58 V67 -7.19369933609991e-20

R58_68 V58 V68 8360.905196367423
L58_68 V58 V68 -7.670052756028396e-12
C58_68 V58 V68 2.299265849697267e-21

R58_69 V58 V69 1273.7702000620052
L58_69 V58 V69 5.174354381139548e-12
C58_69 V58 V69 -2.5372157304582568e-20

R58_70 V58 V70 867.3403303033614
L58_70 V58 V70 5.8788277906525984e-12
C58_70 V58 V70 -1.9746359483406072e-20

R58_71 V58 V71 -1113.5278470710914
L58_71 V58 V71 1.7154481894262767e-12
C58_71 V58 V71 8.707426077594325e-20

R58_72 V58 V72 552.1368053539939
L58_72 V58 V72 3.053822361366366e-11
C58_72 V58 V72 -6.141002472238191e-20

R58_73 V58 V73 2607.7583016606454
L58_73 V58 V73 -1.8427103601789305e-12
C58_73 V58 V73 -3.139781799592219e-20

R58_74 V58 V74 1690.8278242687088
L58_74 V58 V74 9.145537945149324e-12
C58_74 V58 V74 1.1515593682440662e-20

R58_75 V58 V75 -1685.2536705389234
L58_75 V58 V75 -2.168706859693292e-11
C58_75 V58 V75 7.220868862750708e-21

R58_76 V58 V76 -791.9550154664233
L58_76 V58 V76 -1.2733006844254056e-12
C58_76 V58 V76 8.169245331892591e-20

R58_77 V58 V77 -1521.441416622505
L58_77 V58 V77 -3.800434251210232e-12
C58_77 V58 V77 6.346509063215922e-20

R58_78 V58 V78 -5344.5506733208995
L58_78 V58 V78 -2.766789131451101e-12
C58_78 V58 V78 -2.194444910983637e-20

R58_79 V58 V79 214976.40600054193
L58_79 V58 V79 -5.3393557651393956e-12
C58_79 V58 V79 7.324930089552048e-20

R58_80 V58 V80 3142.215387844759
L58_80 V58 V80 3.4933675631034665e-12
C58_80 V58 V80 -4.923615086256503e-20

R58_81 V58 V81 5889.224106813261
L58_81 V58 V81 -1.0411578671381665e-11
C58_81 V58 V81 -5.68750115499231e-20

R58_82 V58 V82 14598.322602684897
L58_82 V58 V82 3.583227022692903e-12
C58_82 V58 V82 5.922092761384284e-20

R58_83 V58 V83 -105843.5564068408
L58_83 V58 V83 2.029970089047803e-12
C58_83 V58 V83 7.284912179404149e-20

R58_84 V58 V84 -9071.42810281057
L58_84 V58 V84 -3.365866717132801e-12
C58_84 V58 V84 -2.76596219490449e-21

R58_85 V58 V85 5045.443616936655
L58_85 V58 V85 -3.37704098042766e-12
C58_85 V58 V85 -2.75873354295859e-20

R58_86 V58 V86 7207.054388902555
L58_86 V58 V86 -2.8792881362642524e-12
C58_86 V58 V86 -3.316426773800674e-20

R58_87 V58 V87 -10012.71658994423
L58_87 V58 V87 -5.874846796906737e-12
C58_87 V58 V87 -7.644574450794823e-21

R58_88 V58 V88 10158.989391105875
L58_88 V58 V88 -2.8136411615719753e-10
C58_88 V58 V88 -1.085268569973943e-20

R58_89 V58 V89 -8542.191039693953
L58_89 V58 V89 7.91534599280867e-12
C58_89 V58 V89 2.2416176785798812e-20

R58_90 V58 V90 17554.788360699218
L58_90 V58 V90 7.132006714305163e-12
C58_90 V58 V90 -2.713124426624348e-20

R58_91 V58 V91 9135.96327505806
L58_91 V58 V91 4.415865707669972e-12
C58_91 V58 V91 5.3455490792772393e-20

R58_92 V58 V92 -37099.02620020654
L58_92 V58 V92 5.218410999169314e-12
C58_92 V58 V92 4.284114606543176e-20

R58_93 V58 V93 2375.165074040087
L58_93 V58 V93 -4.423258037706092e-11
C58_93 V58 V93 -1.9515867202796678e-22

R58_94 V58 V94 3975.350380163783
L58_94 V58 V94 -1.215337123768456e-11
C58_94 V58 V94 -5.432985683581002e-20

R58_95 V58 V95 -6604.590186548176
L58_95 V58 V95 6.722768611938694e-12
C58_95 V58 V95 4.13295458214023e-20

R58_96 V58 V96 -5655.433936438376
L58_96 V58 V96 6.751876511098919e-12
C58_96 V58 V96 2.761369948865848e-20

R58_97 V58 V97 2833.1503861272545
L58_97 V58 V97 -8.607182546757992e-12
C58_97 V58 V97 -4.936481206249756e-20

R58_98 V58 V98 3737.683553884812
L58_98 V58 V98 5.457420769177377e-12
C58_98 V58 V98 3.0357561254482815e-20

R58_99 V58 V99 18960.989625258782
L58_99 V58 V99 -5.6251906263226295e-11
C58_99 V58 V99 -1.9437078029666452e-21

R58_100 V58 V100 -15892.21921999865
L58_100 V58 V100 -1.4477776723050999e-11
C58_100 V58 V100 -2.3732865114608163e-20

R58_101 V58 V101 3622.1421199530573
L58_101 V58 V101 5.234119012622229e-12
C58_101 V58 V101 3.957554247287355e-20

R58_102 V58 V102 10845.320800954194
L58_102 V58 V102 4.101945613176181e-12
C58_102 V58 V102 -3.570511206443949e-21

R58_103 V58 V103 3107.75774527365
L58_103 V58 V103 -1.5001002969309887e-11
C58_103 V58 V103 3.3657469502772564e-20

R58_104 V58 V104 -9137.80785880405
L58_104 V58 V104 3.766602643198916e-11
C58_104 V58 V104 9.904399077787801e-21

R58_105 V58 V105 -2279.909884137854
L58_105 V58 V105 -4.49626838851169e-12
C58_105 V58 V105 -5.007553652315376e-20

R58_106 V58 V106 -4014.6402486688207
L58_106 V58 V106 3.2628988899417143e-12
C58_106 V58 V106 5.081270452753021e-20

R58_107 V58 V107 17885.32342179006
L58_107 V58 V107 1.0276817457884709e-11
C58_107 V58 V107 -4.147757368384639e-20

R58_108 V58 V108 -3416.6829317578467
L58_108 V58 V108 -6.547498972983284e-12
C58_108 V58 V108 1.3111206316082344e-20

R58_109 V58 V109 161704.0211983515
L58_109 V58 V109 -3.438359306319594e-10
C58_109 V58 V109 2.180084481403757e-20

R58_110 V58 V110 -5527.301115918228
L58_110 V58 V110 -3.5737660698224324e-12
C58_110 V58 V110 -5.837096295894006e-20

R58_111 V58 V111 25445.68267088382
L58_111 V58 V111 -7.995156796559088e-12
C58_111 V58 V111 -1.1050366102444967e-20

R58_112 V58 V112 -5359.2289198408025
L58_112 V58 V112 6.079113986040671e-12
C58_112 V58 V112 7.433099611467065e-21

R58_113 V58 V113 -3834.1298431029413
L58_113 V58 V113 1.5727133249399772e-11
C58_113 V58 V113 7.660957556897336e-21

R58_114 V58 V114 13845.953210957414
L58_114 V58 V114 6.9430942380961085e-12
C58_114 V58 V114 3.2658127113445983e-20

R58_115 V58 V115 -6100.225589172786
L58_115 V58 V115 6.691125649091071e-11
C58_115 V58 V115 -3.079377281178596e-20

R58_116 V58 V116 -84635.9590531582
L58_116 V58 V116 -1.0173309695145774e-11
C58_116 V58 V116 -3.2451634111243224e-21

R58_117 V58 V117 3887.23604026656
L58_117 V58 V117 -1.851641537350625e-11
C58_117 V58 V117 9.201944558213287e-22

R58_118 V58 V118 -4077.676128635282
L58_118 V58 V118 -9.958769523052525e-12
C58_118 V58 V118 -1.4518048133914644e-20

R58_119 V58 V119 -4064.8936471349134
L58_119 V58 V119 -6.2657350477868555e-12
C58_119 V58 V119 -2.6907693481876364e-20

R58_120 V58 V120 2928.8473889168436
L58_120 V58 V120 -2.2726375877038442e-11
C58_120 V58 V120 1.3887192667833814e-21

R58_121 V58 V121 -6571.746497122314
L58_121 V58 V121 2.146688157578478e-11
C58_121 V58 V121 1.3158287894618665e-20

R58_122 V58 V122 -2542.978733089763
L58_122 V58 V122 -9.14956255583063e-11
C58_122 V58 V122 2.05993451357996e-21

R58_123 V58 V123 6529.518173392413
L58_123 V58 V123 -2.144056374364736e-11
C58_123 V58 V123 -1.3308321464842647e-20

R58_124 V58 V124 22704.76237995534
L58_124 V58 V124 -3.7166439710004913e-11
C58_124 V58 V124 -1.4072142750680715e-21

R58_125 V58 V125 3754.3720312126184
L58_125 V58 V125 -2.514250556153109e-11
C58_125 V58 V125 -2.6389089990437904e-21

R58_126 V58 V126 4968.469280250103
L58_126 V58 V126 1.9242317973126957e-11
C58_126 V58 V126 7.764176867097735e-21

R58_127 V58 V127 14102.987216708252
L58_127 V58 V127 1.1892460218994419e-10
C58_127 V58 V127 -1.271944680724431e-22

R58_128 V58 V128 6594.31345369474
L58_128 V58 V128 5.7039838951480805e-11
C58_128 V58 V128 -8.122976121447643e-21

R58_129 V58 V129 5563.011413464966
L58_129 V58 V129 -4.1861559708710836e-11
C58_129 V58 V129 -1.101881371896868e-20

R58_130 V58 V130 -56240.544837694426
L58_130 V58 V130 7.604368076971949e-11
C58_130 V58 V130 6.162588602433212e-21

R58_131 V58 V131 22939.06445690488
L58_131 V58 V131 1.321597000488945e-11
C58_131 V58 V131 1.0411243901351089e-20

R58_132 V58 V132 -180723.26764734875
L58_132 V58 V132 -3.5082888271901146e-11
C58_132 V58 V132 -9.781521355635448e-21

R58_133 V58 V133 -31349.417286846907
L58_133 V58 V133 9.783320414683635e-12
C58_133 V58 V133 1.424564043377912e-20

R58_134 V58 V134 -4163.162924669255
L58_134 V58 V134 2.247591552411009e-10
C58_134 V58 V134 2.5324366199273017e-21

R58_135 V58 V135 19849.205684826702
L58_135 V58 V135 3.0534023153456634e-09
C58_135 V58 V135 1.1251215025279999e-20

R58_136 V58 V136 13895.532034376973
L58_136 V58 V136 5.194604279175441e-11
C58_136 V58 V136 1.1299538998351413e-20

R58_137 V58 V137 2933.479760474319
L58_137 V58 V137 -1.4580608494580728e-10
C58_137 V58 V137 6.1503591701304e-21

R58_138 V58 V138 3329.1973850512054
L58_138 V58 V138 2.7888222133784006e-11
C58_138 V58 V138 -9.938863836142842e-21

R58_139 V58 V139 30827.320640737027
L58_139 V58 V139 -5.919591300048201e-10
C58_139 V58 V139 -6.16567073772707e-21

R58_140 V58 V140 -2417.4995200090234
L58_140 V58 V140 -2.922923500910796e-11
C58_140 V58 V140 -2.714941334095449e-21

R58_141 V58 V141 4994.847538136733
L58_141 V58 V141 -2.932913734355994e-10
C58_141 V58 V141 3.159625147536397e-21

R58_142 V58 V142 -2313.2259263476103
L58_142 V58 V142 -2.1390238633098387e-11
C58_142 V58 V142 -2.733390620362442e-20

R58_143 V58 V143 -12796.098201798477
L58_143 V58 V143 2.3009960939312922e-11
C58_143 V58 V143 1.026532611136869e-20

R58_144 V58 V144 38781.50079072405
L58_144 V58 V144 -1.4638250949201285e-10
C58_144 V58 V144 -1.7123897364814656e-20

R59_59 V59 0 148.91597563368703
L59_59 V59 0 2.1812963898662306e-13
C59_59 V59 0 -8.2694325342893e-19

R59_60 V59 V60 -3904.8410928748035
L59_60 V59 V60 -4.9329082023067745e-12
C59_60 V59 V60 -2.6680328771632116e-20

R59_61 V59 V61 912.2709152003845
L59_61 V59 V61 3.408239918948514e-12
C59_61 V59 V61 1.1179262034215708e-19

R59_62 V59 V62 -1533.8975624994378
L59_62 V59 V62 -1.288246714755358e-12
C59_62 V59 V62 1.8231662798695856e-19

R59_63 V59 V63 3886.117195057281
L59_63 V59 V63 -8.069897058456296e-12
C59_63 V59 V63 -7.231022539368313e-20

R59_64 V59 V64 -3161.0026693772784
L59_64 V59 V64 -4.331586932959562e-12
C59_64 V59 V64 8.333600380069068e-21

R59_65 V59 V65 -998.3259824174806
L59_65 V59 V65 -1.962665056092737e-11
C59_65 V59 V65 1.2823609987726017e-19

R59_66 V59 V66 -2229.0503544654116
L59_66 V59 V66 -3.190407347849252e-12
C59_66 V59 V66 -4.0130208325570166e-20

R59_67 V59 V67 -1692.5740508077463
L59_67 V59 V67 -1.3825966653654452e-12
C59_67 V59 V67 -6.307502503656723e-20

R59_68 V59 V68 2664.9326919870005
L59_68 V59 V68 3.1954150263625192e-12
C59_68 V59 V68 1.4177307841423967e-20

R59_69 V59 V69 995.6302029844618
L59_69 V59 V69 1.178521195678713e-12
C59_69 V59 V69 -6.113302361273299e-20

R59_70 V59 V70 -3984.503265462378
L59_70 V59 V70 -2.407313145534386e-12
C59_70 V59 V70 -5.371184516186762e-20

R59_71 V59 V71 7265.191440069346
L59_71 V59 V71 4.506755731424414e-12
C59_71 V59 V71 1.0995422771539113e-21

R59_72 V59 V72 -101406.13115015007
L59_72 V59 V72 -4.1559011457860034e-12
C59_72 V59 V72 -4.6549342570472824e-20

R59_73 V59 V73 8223.879892651037
L59_73 V59 V73 -1.2026409340582692e-11
C59_73 V59 V73 2.951977322770842e-21

R59_74 V59 V74 3107.1478741491705
L59_74 V59 V74 5.245914453641709e-12
C59_74 V59 V74 2.1881898017672033e-20

R59_75 V59 V75 -94771.99885567346
L59_75 V59 V75 5.928484095830172e-12
C59_75 V59 V75 8.473723886961117e-20

R59_76 V59 V76 -11912.53636886376
L59_76 V59 V76 -2.43538884461043e-11
C59_76 V59 V76 4.3929672869087834e-20

R59_77 V59 V77 -26187.297814544614
L59_77 V59 V77 -6.638556700638867e-11
C59_77 V59 V77 1.5388069722830428e-20

R59_78 V59 V78 -4379.17984329864
L59_78 V59 V78 -1.8121230640618435e-12
C59_78 V59 V78 -1.6213038062979463e-19

R59_79 V59 V79 15456.264086368132
L59_79 V59 V79 -3.306355075817169e-11
C59_79 V59 V79 1.3928199753081477e-20

R59_80 V59 V80 21341.596262223233
L59_80 V59 V80 1.376140644041453e-10
C59_80 V59 V80 -2.876734880604372e-20

R59_81 V59 V81 26528.32523941044
L59_81 V59 V81 6.350281818033419e-11
C59_81 V59 V81 1.587742311831967e-20

R59_82 V59 V82 5977.1183068150585
L59_82 V59 V82 1.897190595716819e-12
C59_82 V59 V82 2.5722005567795573e-19

R59_83 V59 V83 8878.68102229667
L59_83 V59 V83 2.0969105784772505e-12
C59_83 V59 V83 1.9382242012677502e-19

R59_84 V59 V84 1298827.1153535962
L59_84 V59 V84 -2.2008081267041177e-11
C59_84 V59 V84 -9.008274935787179e-21

R59_85 V59 V85 301294.9972063492
L59_85 V59 V85 -5.90470204684902e-12
C59_85 V59 V85 -8.296145095294418e-20

R59_86 V59 V86 -32882.308543633204
L59_86 V59 V86 -4.546686022656481e-12
C59_86 V59 V86 -7.202835324300685e-20

R59_87 V59 V87 87559.85709241411
L59_87 V59 V87 -4.720022573222791e-12
C59_87 V59 V87 -7.645361776270973e-20

R59_88 V59 V88 -124486.03108095913
L59_88 V59 V88 -1.60941498520022e-11
C59_88 V59 V88 -2.3055843654977825e-20

R59_89 V59 V89 -38972.844646672376
L59_89 V59 V89 1.0041627257281069e-11
C59_89 V59 V89 5.750870529727949e-20

R59_90 V59 V90 38383.1439878455
L59_90 V59 V90 1.65422838267682e-11
C59_90 V59 V90 2.839067580039582e-20

R59_91 V59 V91 12218.997328232803
L59_91 V59 V91 2.1548982335815217e-12
C59_91 V59 V91 2.1196559005189697e-19

R59_92 V59 V92 17170.646751876608
L59_92 V59 V92 5.99562814174155e-12
C59_92 V59 V92 6.053830656776544e-20

R59_93 V59 V93 16647.78526845034
L59_93 V59 V93 -1.9565031234695323e-11
C59_93 V59 V93 -2.516763298214665e-20

R59_94 V59 V94 73360.2406975455
L59_94 V59 V94 -6.174123735938177e-12
C59_94 V59 V94 -8.309716915776753e-20

R59_95 V59 V95 16980.35849280309
L59_95 V59 V95 3.846643258705258e-12
C59_95 V59 V95 1.268489737046728e-19

R59_96 V59 V96 -7358.907427727749
L59_96 V59 V96 3.678303094758492e-11
C59_96 V59 V96 -4.167722294515092e-21

R59_97 V59 V97 -15783.1932653084
L59_97 V59 V97 -7.158386605020976e-12
C59_97 V59 V97 -5.633193802353592e-20

R59_98 V59 V98 11950.925512132175
L59_98 V59 V98 5.274457201916008e-12
C59_98 V59 V98 8.895103290727626e-20

R59_99 V59 V99 17488.258576374585
L59_99 V59 V99 -4.4215217219958804e-11
C59_99 V59 V99 -1.1420782148861021e-20

R59_100 V59 V100 -14764.267389774282
L59_100 V59 V100 -1.966466459921096e-11
C59_100 V59 V100 -8.785469599180367e-21

R59_101 V59 V101 29163.737915670492
L59_101 V59 V101 5.787826543439267e-12
C59_101 V59 V101 7.861601568071203e-20

R59_102 V59 V102 5212.99106368611
L59_102 V59 V102 3.930852754203652e-12
C59_102 V59 V102 1.4979919348366378e-19

R59_103 V59 V103 37064.791861044585
L59_103 V59 V103 -4.1655164173057824e-11
C59_103 V59 V103 -1.187141443758104e-20

R59_104 V59 V104 -26021.39673676478
L59_104 V59 V104 -1.3820419754756098e-11
C59_104 V59 V104 -3.7053401338773294e-20

R59_105 V59 V105 -9421.00202916886
L59_105 V59 V105 -3.418814655568468e-12
C59_105 V59 V105 -1.4207429371131138e-19

R59_106 V59 V106 944029.9767836699
L59_106 V59 V106 2.1125394557114647e-12
C59_106 V59 V106 2.259767602628001e-19

R59_107 V59 V107 114484.75876237563
L59_107 V59 V107 6.789775390089694e-12
C59_107 V59 V107 8.480809544584665e-20

R59_108 V59 V108 -14631.331908866232
L59_108 V59 V108 -8.325163549157567e-12
C59_108 V59 V108 -5.561730053324619e-20

R59_109 V59 V109 -1234625.0129972626
L59_109 V59 V109 -1.1556021374080031e-11
C59_109 V59 V109 -6.646022132893376e-20

R59_110 V59 V110 20486.42821302434
L59_110 V59 V110 -2.173715145517395e-12
C59_110 V59 V110 -2.4770991041333945e-19

R59_111 V59 V111 -13655.409935098927
L59_111 V59 V111 -5.739843381141256e-12
C59_111 V59 V111 -8.440473369039935e-20

R59_112 V59 V112 10356.262910587506
L59_112 V59 V112 6.333765608973653e-12
C59_112 V59 V112 7.20945605555785e-20

R59_113 V59 V113 -50886.736034006164
L59_113 V59 V113 8.420756216464552e-12
C59_113 V59 V113 6.638349625589227e-20

R59_114 V59 V114 -24062.29429653065
L59_114 V59 V114 4.3946463127257964e-12
C59_114 V59 V114 1.2596251025169867e-19

R59_115 V59 V115 8404.369840883486
L59_115 V59 V115 1.6605765195808323e-11
C59_115 V59 V115 2.835506625858073e-20

R59_116 V59 V116 -9132.308352678965
L59_116 V59 V116 -7.77594402897019e-12
C59_116 V59 V116 -6.229762545478805e-20

R59_117 V59 V117 -36097.47528847169
L59_117 V59 V117 -9.753596220873483e-12
C59_117 V59 V117 -6.783543448291857e-20

R59_118 V59 V118 -147676.024948964
L59_118 V59 V118 -4.655019432510579e-12
C59_118 V59 V118 -1.0770340623280243e-19

R59_119 V59 V119 -15049.863275754784
L59_119 V59 V119 -3.975357479844632e-12
C59_119 V59 V119 -1.1520813084165232e-19

R59_120 V59 V120 9336.608260922934
L59_120 V59 V120 7.648002447888548e-11
C59_120 V59 V120 -6.658583541487282e-21

R59_121 V59 V121 44079.88850996226
L59_121 V59 V121 1.1542771521461986e-11
C59_121 V59 V121 5.124980481819485e-20

R59_122 V59 V122 39832.78725477499
L59_122 V59 V122 9.209969577375253e-11
C59_122 V59 V122 -1.0903829022628523e-20

R59_123 V59 V123 536267.2956688545
L59_123 V59 V123 -9.55965628253692e-12
C59_123 V59 V123 -5.733623663128054e-20

R59_124 V59 V124 22910.587375908806
L59_124 V59 V124 -1.4826218529093144e-11
C59_124 V59 V124 -1.5764809226297154e-20

R59_125 V59 V125 14122.813076869785
L59_125 V59 V125 -2.941042877875333e-11
C59_125 V59 V125 -2.5004186091955255e-20

R59_126 V59 V126 -12370.779562806505
L59_126 V59 V126 -9.236429632822301e-11
C59_126 V59 V126 2.2973968551868033e-20

R59_127 V59 V127 7455.880506586069
L59_127 V59 V127 1.8481854538504102e-11
C59_127 V59 V127 2.769578136799445e-21

R59_128 V59 V128 16674.58741049443
L59_128 V59 V128 -8.427917035309871e-10
C59_128 V59 V128 -2.384039166042109e-20

R59_129 V59 V129 9940.66826847145
L59_129 V59 V129 -2.099604814417846e-11
C59_129 V59 V129 -3.047440253523231e-20

R59_130 V59 V130 14655.918763595855
L59_130 V59 V130 3.665577313145174e-10
C59_130 V59 V130 -1.5076069314109715e-20

R59_131 V59 V131 33670.123910903836
L59_131 V59 V131 1.2289002241179147e-11
C59_131 V59 V131 4.1867479676606503e-20

R59_132 V59 V132 -49186.6953636898
L59_132 V59 V132 -6.096329079609051e-11
C59_132 V59 V132 -1.1251778825948694e-20

R59_133 V59 V133 -73731.47093035611
L59_133 V59 V133 8.743867365320498e-12
C59_133 V59 V133 3.639597327850594e-20

R59_134 V59 V134 28473.13288057782
L59_134 V59 V134 -1.3001090884305511e-08
C59_134 V59 V134 4.472879755816584e-21

R59_135 V59 V135 109666.2191698314
L59_135 V59 V135 4.15005016807082e-11
C59_135 V59 V135 6.378707835731297e-22

R59_136 V59 V136 56080.49769894393
L59_136 V59 V136 3.074249576024653e-11
C59_136 V59 V136 2.2592641159054726e-20

R59_137 V59 V137 7302.738082204011
L59_137 V59 V137 -8.692512698638714e-10
C59_137 V59 V137 1.2627714963868315e-20

R59_138 V59 V138 -27414.37096086376
L59_138 V59 V138 -1.9838502106075145e-11
C59_138 V59 V138 -3.37474905399717e-20

R59_139 V59 V139 9375.906172398783
L59_139 V59 V139 1.3947399809102214e-11
C59_139 V59 V139 -2.582229341683678e-21

R59_140 V59 V140 -15011.422373160178
L59_140 V59 V140 -1.1766350850256872e-10
C59_140 V59 V140 9.502553132055724e-22

R59_141 V59 V141 30917.011803877118
L59_141 V59 V141 -2.17666929065223e-11
C59_141 V59 V141 -1.2594703487466754e-20

R59_142 V59 V142 -6490.906017899364
L59_142 V59 V142 -9.267027514505328e-12
C59_142 V59 V142 -6.441903440708095e-20

R59_143 V59 V143 -27750.21626088232
L59_143 V59 V143 -4.658343471100732e-11
C59_143 V59 V143 -1.1474724266419525e-20

R59_144 V59 V144 -13626.443515675748
L59_144 V59 V144 -5.585169781951836e-11
C59_144 V59 V144 -9.47467420539101e-21

R60_60 V60 0 33.30987449310553
L60_60 V60 0 4.532131885109829e-14
C60_60 V60 0 -3.0418757187520924e-19

R60_61 V60 V61 447.00882410250415
L60_61 V60 V61 2.737221967690216e-12
C60_61 V60 V61 2.4920757394151183e-20

R60_62 V60 V62 3003.3921003704427
L60_62 V60 V62 -1.7651359671691223e-12
C60_62 V60 V62 4.085303548181719e-20

R60_63 V60 V63 5520.882351577397
L60_63 V60 V63 -4.115360045257228e-12
C60_63 V60 V63 -2.8850018686928214e-21

R60_64 V60 V64 3577.944955627205
L60_64 V60 V64 -1.037937978805232e-12
C60_64 V60 V64 -2.792472784332992e-20

R60_65 V60 V65 -346.8986909196164
L60_65 V60 V65 -8.109888210939208e-13
C60_65 V60 V65 2.3806724965300295e-20

R60_66 V60 V66 -456.6146948914421
L60_66 V60 V66 -7.06551132835331e-13
C60_66 V60 V66 -1.4157968412036782e-21

R60_67 V60 V67 -1318.247573423893
L60_67 V60 V67 -1.789812887395553e-12
C60_67 V60 V67 -9.268951126598032e-22

R60_68 V60 V68 -361.69540545613427
L60_68 V60 V68 -5.40881371355329e-13
C60_68 V60 V68 2.821434853045491e-20

R60_69 V60 V69 744.0443041622215
L60_69 V60 V69 1.0730373636189756e-12
C60_69 V60 V69 -3.093619962304601e-20

R60_70 V60 V70 8824.141802221464
L60_70 V60 V70 -5.288572221329336e-12
C60_70 V60 V70 -1.9540426299479413e-20

R60_71 V60 V71 4229.502486392565
L60_71 V60 V71 -8.893141820569142e-12
C60_71 V60 V71 -2.5982392583870423e-20

R60_72 V60 V72 1071.0618529879887
L60_72 V60 V72 2.509131539058489e-12
C60_72 V60 V72 -4.847634590298665e-21

R60_73 V60 V73 -1798.8519721040689
L60_73 V60 V73 -2.663965883155725e-12
C60_73 V60 V73 7.161698163869685e-21

R60_74 V60 V74 2135.1461910471608
L60_74 V60 V74 3.1399428147467543e-12
C60_74 V60 V74 -1.118483761567118e-21

R60_75 V60 V75 -4067.159166128837
L60_75 V60 V75 -8.766292984974686e-12
C60_75 V60 V75 4.10320441818135e-20

R60_76 V60 V76 -2561.9656906962864
L60_76 V60 V76 -1.992409905798584e-12
C60_76 V60 V76 -2.129461563575031e-20

R60_77 V60 V77 6825.421731219262
L60_77 V60 V77 4.163119618217644e-12
C60_77 V60 V77 1.7874545047370503e-20

R60_78 V60 V78 -15384.538638178981
L60_78 V60 V78 -4.095985633592845e-12
C60_78 V60 V78 -1.7398316974042865e-20

R60_79 V60 V79 8767.20197679362
L60_79 V60 V79 -1.2789926710528146e-11
C60_79 V60 V79 -4.956087924979305e-20

R60_80 V60 V80 4383.053711216148
L60_80 V60 V80 3.223359829827469e-12
C60_80 V60 V80 7.761379090851762e-20

R60_81 V60 V81 -11541.700091013681
L60_81 V60 V81 -3.3706293018559955e-12
C60_81 V60 V81 -3.50892420016246e-20

R60_82 V60 V82 1154761.1163508904
L60_82 V60 V82 9.408442727331538e-12
C60_82 V60 V82 5.131961758244746e-20

R60_83 V60 V83 9132.054256291252
L60_83 V60 V83 5.370857021248536e-12
C60_83 V60 V83 7.057333404567186e-20

R60_84 V60 V84 8375.541026792584
L60_84 V60 V84 1.139996579497422e-10
C60_84 V60 V84 -2.566999034849369e-22

R60_85 V60 V85 15657.504288319005
L60_85 V60 V85 -1.1058388278515493e-11
C60_85 V60 V85 -4.17617976795239e-20

R60_86 V60 V86 -6462.030938842008
L60_86 V60 V86 -4.892309877030567e-11
C60_86 V60 V86 -2.2380240199326703e-20

R60_87 V60 V87 237167.78201951398
L60_87 V60 V87 -9.449659155018945e-12
C60_87 V60 V87 -2.5527062459649595e-20

R60_88 V60 V88 18908.473160664504
L60_88 V60 V88 -3.1222465016572355e-11
C60_88 V60 V88 6.718801636728116e-21

R60_89 V60 V89 -28861.104037588844
L60_89 V60 V89 8.816314058459398e-12
C60_89 V60 V89 4.058094715182638e-20

R60_90 V60 V90 -88847.37013460428
L60_90 V60 V90 1.1555405998452827e-11
C60_90 V60 V90 5.788306601207973e-20

R60_91 V60 V91 22942.463758510938
L60_91 V60 V91 5.472406576470825e-11
C60_91 V60 V91 5.205766773391494e-20

R60_92 V60 V92 -95153.83197167453
L60_92 V60 V92 3.6279665814406593e-12
C60_92 V60 V92 6.868645102086232e-20

R60_93 V60 V93 3502.3339502123863
L60_93 V60 V93 -3.728552527454686e-11
C60_93 V60 V93 -8.537730638819719e-21

R60_94 V60 V94 8694.360205554121
L60_94 V60 V94 -8.913450683668445e-12
C60_94 V60 V94 -2.733011308961106e-20

R60_95 V60 V95 20259.314913206497
L60_95 V60 V95 3.5111929461709403e-11
C60_95 V60 V95 2.770204998610807e-20

R60_96 V60 V96 29817.886799678112
L60_96 V60 V96 3.5019863939138474e-12
C60_96 V60 V96 4.246021078214553e-20

R60_97 V60 V97 9106.979823873486
L60_97 V60 V97 -4.0776358891808594e-11
C60_97 V60 V97 1.0818220731145095e-20

R60_98 V60 V98 4319.102317442757
L60_98 V60 V98 7.110763069362556e-12
C60_98 V60 V98 4.731979698495567e-20

R60_99 V60 V99 9462.557824691447
L60_99 V60 V99 -1.7531702648553586e-11
C60_99 V60 V99 -1.5738486345214804e-20

R60_100 V60 V100 13052.510685945166
L60_100 V60 V100 -1.545883397479187e-11
C60_100 V60 V100 -3.497446301829412e-22

R60_101 V60 V101 8911.737358142822
L60_101 V60 V101 9.693682670084287e-12
C60_101 V60 V101 3.3740758488417704e-20

R60_102 V60 V102 5145.12358066489
L60_102 V60 V102 6.3342423278202864e-12
C60_102 V60 V102 1.1132417934918721e-19

R60_103 V60 V103 141020.51255512235
L60_103 V60 V103 -1.961108215181775e-11
C60_103 V60 V103 -3.6598596360654144e-20

R60_104 V60 V104 -14079.940370167664
L60_104 V60 V104 5.056603342315219e-12
C60_104 V60 V104 4.7075204350293875e-20

R60_105 V60 V105 -36347.1785498741
L60_105 V60 V105 -6.36713846632822e-12
C60_105 V60 V105 -7.292754773953484e-20

R60_106 V60 V106 -8710.629427913836
L60_106 V60 V106 6.422677203998671e-12
C60_106 V60 V106 1.0060099308473679e-19

R60_107 V60 V107 10029.86199350314
L60_107 V60 V107 6.712244174941055e-12
C60_107 V60 V107 9.532587009578459e-20

R60_108 V60 V108 8749.064115486162
L60_108 V60 V108 -5.2438041376181304e-12
C60_108 V60 V108 -9.088737883667264e-20

R60_109 V60 V109 -5699.404286230251
L60_109 V60 V109 1.27647603899532e-11
C60_109 V60 V109 -1.4827913920550618e-20

R60_110 V60 V110 -19535.527913430542
L60_110 V60 V110 -7.124520732345288e-12
C60_110 V60 V110 -7.838776930159589e-20

R60_111 V60 V111 -12191.883354513982
L60_111 V60 V111 -1.175531656464764e-11
C60_111 V60 V111 -3.8362063933190693e-20

R60_112 V60 V112 279177.7116078079
L60_112 V60 V112 8.113391958742892e-12
C60_112 V60 V112 4.88151482521367e-20

R60_113 V60 V113 10610.917238139093
L60_113 V60 V113 2.0160266350176336e-11
C60_113 V60 V113 5.453336532222092e-20

R60_114 V60 V114 10072.657540305125
L60_114 V60 V114 1.8081821298665856e-11
C60_114 V60 V114 1.545757602850771e-20

R60_115 V60 V115 8443.288769473598
L60_115 V60 V115 1.2609407238592132e-11
C60_115 V60 V115 4.95925667763181e-20

R60_116 V60 V116 23128.54099639024
L60_116 V60 V116 -7.467634571950599e-12
C60_116 V60 V116 -5.409775891956271e-20

R60_117 V60 V117 92245.00196069639
L60_117 V60 V117 -2.068656435005813e-11
C60_117 V60 V117 -6.535374704574723e-20

R60_118 V60 V118 -5878.881961740932
L60_118 V60 V118 -1.961915972374484e-11
C60_118 V60 V118 -5.1306833920715306e-20

R60_119 V60 V119 -8311.99869706143
L60_119 V60 V119 -8.464710888694655e-12
C60_119 V60 V119 -3.4192886317172e-20

R60_120 V60 V120 5915.721595076974
L60_120 V60 V120 -3.424181967262735e-11
C60_120 V60 V120 -1.1922196144153826e-20

R60_121 V60 V121 -9226.194593201448
L60_121 V60 V121 6.705852608367361e-11
C60_121 V60 V121 5.4407875776587435e-21

R60_122 V60 V122 -13351.231516963466
L60_122 V60 V122 1.6907589792409882e-11
C60_122 V60 V122 -2.7712081208148033e-21

R60_123 V60 V123 19517.23414036099
L60_123 V60 V123 -1.231237403434356e-10
C60_123 V60 V123 -1.2060752886572432e-20

R60_124 V60 V124 7756.122480720046
L60_124 V60 V124 -1.2744620297579014e-11
C60_124 V60 V124 -2.891972479712733e-20

R60_125 V60 V125 6619.372010503734
L60_125 V60 V125 -2.7870404889253784e-11
C60_125 V60 V125 -1.5122172808769576e-20

R60_126 V60 V126 8994.743340104074
L60_126 V60 V126 -1.523322783146528e-11
C60_126 V60 V126 4.8006002559820166e-21

R60_127 V60 V127 10651.396624197661
L60_127 V60 V127 1.937290884895109e-11
C60_127 V60 V127 5.0814125409884846e-21

R60_128 V60 V128 21819.66368354027
L60_128 V60 V128 -2.9595845099305054e-11
C60_128 V60 V128 -2.773312181404364e-20

R60_129 V60 V129 7284.556735609485
L60_129 V60 V129 -1.592223711040612e-10
C60_129 V60 V129 -8.292272054298756e-21

R60_130 V60 V130 -29305.58187986719
L60_130 V60 V130 -1.2455742080357238e-11
C60_130 V60 V130 -5.0538892709366445e-20

R60_131 V60 V131 -184878.1429215219
L60_131 V60 V131 -6.517755180502209e-10
C60_131 V60 V131 6.583340727378902e-21

R60_132 V60 V132 -20118.210871258474
L60_132 V60 V132 -1.0996619315958874e-11
C60_132 V60 V132 -2.0648073252979577e-20

R60_133 V60 V133 -65200.833948199615
L60_133 V60 V133 1.4455144855708423e-11
C60_133 V60 V133 4.621816958572404e-20

R60_134 V60 V134 -5741.791110718361
L60_134 V60 V134 -6.755465712544692e-11
C60_134 V60 V134 4.78339409489611e-21

R60_135 V60 V135 -75527.29194495545
L60_135 V60 V135 5.493941090331976e-11
C60_135 V60 V135 -1.6589106601675496e-20

R60_136 V60 V136 28562.35924370134
L60_136 V60 V136 5.407330644460698e-11
C60_136 V60 V136 1.5393424330381968e-20

R60_137 V60 V137 3988.7166077160546
L60_137 V60 V137 -2.3439623043991e-11
C60_137 V60 V137 -1.5897876298169938e-20

R60_138 V60 V138 29975.089151476466
L60_138 V60 V138 -1.7724064200305002e-11
C60_138 V60 V138 1.0080563121890175e-20

R60_139 V60 V139 6770.243254126943
L60_139 V60 V139 1.2806897532868716e-11
C60_139 V60 V139 1.3286253750790388e-20

R60_140 V60 V140 -8454.541962784491
L60_140 V60 V140 -2.0137560412168555e-11
C60_140 V60 V140 -7.291662515097919e-21

R60_141 V60 V141 15209.903465324407
L60_141 V60 V141 6.384511259146412e-11
C60_141 V60 V141 1.5989229674022133e-20

R60_142 V60 V142 -17138.663210709004
L60_142 V60 V142 -2.4232787767031043e-11
C60_142 V60 V142 -2.0219841252149407e-20

R60_143 V60 V143 73607.68972807947
L60_143 V60 V143 -2.7569137376218937e-11
C60_143 V60 V143 -7.704447724529039e-21

R60_144 V60 V144 -26159.462336678585
L60_144 V60 V144 1.7753914945271386e-11
C60_144 V60 V144 4.415168785342551e-22

R61_61 V61 0 -33.87314349699966
L61_61 V61 0 -3.486601778089126e-13
C61_61 V61 0 5.681448029970274e-18

R61_62 V61 V62 -299.1059443627253
L61_62 V61 V62 7.99997709514971e-11
C61_62 V61 V62 -6.098036285267093e-19

R61_63 V61 V63 -2898.347884076738
L61_63 V61 V63 2.770976170985923e-12
C61_63 V61 V63 -1.5707874457816814e-19

R61_64 V61 V64 12398.627766900463
L61_64 V61 V64 -5.23574533011767e-12
C61_64 V61 V64 -1.943607765782683e-19

R61_65 V61 V65 202.22905681480304
L61_65 V61 V65 -1.1220205802111401e-11
C61_65 V61 V65 -2.326172796105689e-19

R61_66 V61 V66 231.24413367661543
L61_66 V61 V66 -1.3820527628939594e-12
C61_66 V61 V66 -3.754080836096254e-19

R61_67 V61 V67 1007.8030893829537
L61_67 V61 V67 -1.2280062566539708e-11
C61_67 V61 V67 -1.463988398956344e-19

R61_68 V61 V68 2326.6184935857113
L61_68 V61 V68 5.578313023612296e-12
C61_68 V61 V68 -7.711971428252547e-20

R61_69 V61 V69 -1525.279039499732
L61_69 V61 V69 -4.44175163263017e-12
C61_69 V61 V69 3.0940818321243266e-20

R61_70 V61 V70 -756.6365047915658
L61_70 V61 V70 5.894237995673863e-12
C61_70 V61 V70 -2.270095144958873e-19

R61_71 V61 V71 -1274.9667119893647
L61_71 V61 V71 2.509561583886766e-11
C61_71 V61 V71 -6.923911947967437e-20

R61_72 V61 V72 -755.6982426250713
L61_72 V61 V72 2.4474822667901497e-12
C61_72 V61 V72 3.757455061559556e-21

R61_73 V61 V73 -22307.2007682998
L61_73 V61 V73 4.1551500641259485e-12
C61_73 V61 V73 -1.245519860549263e-19

R61_74 V61 V74 -1520.8312940747317
L61_74 V61 V74 1.6719542236047473e-11
C61_74 V61 V74 1.386311481764382e-19

R61_75 V61 V75 1177.0301362833236
L61_75 V61 V75 -4.4548134172910397e-11
C61_75 V61 V75 8.478180216939037e-21

R61_76 V61 V76 1252.3020836132819
L61_76 V61 V76 -2.074816758822525e-12
C61_76 V61 V76 -3.29230177284357e-19

R61_77 V61 V77 3134.8982675865927
L61_77 V61 V77 -1.134243681479022e-11
C61_77 V61 V77 -3.506397899325761e-20

R61_78 V61 V78 51450.2969404404
L61_78 V61 V78 -3.0922033640340578e-12
C61_78 V61 V78 -2.2333203530561216e-19

R61_79 V61 V79 -3793.5666850219695
L61_79 V61 V79 -6.2611319604106984e-12
C61_79 V61 V79 -1.5187523556142864e-19

R61_80 V61 V80 -4891.1038366631055
L61_80 V61 V80 2.0302210931727404e-12
C61_80 V61 V80 3.294648858690168e-19

R61_81 V61 V81 -4565.320049600324
L61_81 V61 V81 -1.7363568519321214e-11
C61_81 V61 V81 -9.101942870836694e-20

R61_82 V61 V82 4815.190445080664
L61_82 V61 V82 2.634375617783486e-12
C61_82 V61 V82 3.7357544017610376e-19

R61_83 V61 V83 -7820.017662619296
L61_83 V61 V83 1.6515086024528762e-12
C61_83 V61 V83 3.3461538753720405e-19

R61_84 V61 V84 -18516.360867872827
L61_84 V61 V84 -1.6323898289334908e-10
C61_84 V61 V84 -1.1398272087101927e-19

R61_85 V61 V85 -2540.477527994383
L61_85 V61 V85 -5.435673328052661e-12
C61_85 V61 V85 -2.33189509393489e-19

R61_86 V61 V86 -12577.233771533256
L61_86 V61 V86 -7.736406337780535e-12
C61_86 V61 V86 -1.2420210897155652e-19

R61_87 V61 V87 -12064.950549273906
L61_87 V61 V87 -2.2683913453088247e-12
C61_87 V61 V87 -2.953511448276016e-19

R61_88 V61 V88 -16634.71492097216
L61_88 V61 V88 -6.657670515100438e-12
C61_88 V61 V88 -7.041910961680111e-20

R61_89 V61 V89 2717.5544602142786
L61_89 V61 V89 3.4841569859973806e-12
C61_89 V61 V89 2.697628281516876e-19

R61_90 V61 V90 138016.80423236146
L61_90 V61 V90 2.7192542740910785e-12
C61_90 V61 V90 2.040700702099471e-19

R61_91 V61 V91 36829.05747514679
L61_91 V61 V91 2.1677916817666187e-12
C61_91 V61 V91 2.922350997790585e-19

R61_92 V61 V92 8615.92533871958
L61_92 V61 V92 2.383847843492934e-12
C61_92 V61 V92 2.805115900100069e-19

R61_93 V61 V93 -1666.0158552057
L61_93 V61 V93 -8.887509794523274e-12
C61_93 V61 V93 2.4823251810108158e-20

R61_94 V61 V94 -3097.9446654912435
L61_94 V61 V94 -3.981622241164469e-12
C61_94 V61 V94 -1.3068891461950596e-19

R61_95 V61 V95 13798.470857090437
L61_95 V61 V95 3.9706205607096405e-12
C61_95 V61 V95 2.1106191612402e-19

R61_96 V61 V96 4123.111494436167
L61_96 V61 V96 3.6300901571183456e-12
C61_96 V61 V96 2.184423984604068e-19

R61_97 V61 V97 -3712.2350344589536
L61_97 V61 V97 8.047650649868312e-12
C61_97 V61 V97 -7.77599667071662e-21

R61_98 V61 V98 -3633.8771863189845
L61_98 V61 V98 1.7169372593323013e-12
C61_98 V61 V98 2.6094783099707083e-19

R61_99 V61 V99 -4496.553631024639
L61_99 V61 V99 -5.829741061680579e-12
C61_99 V61 V99 -6.275411267961639e-20

R61_100 V61 V100 15050.887328702767
L61_100 V61 V100 -1.300695122047358e-11
C61_100 V61 V100 -5.2265422458998583e-20

R61_101 V61 V101 -11787.369118539538
L61_101 V61 V101 2.1589819413454137e-12
C61_101 V61 V101 3.3282500980062425e-19

R61_102 V61 V102 -32811.815222921854
L61_102 V61 V102 1.0805585811928633e-12
C61_102 V61 V102 5.221952871150575e-19

R61_103 V61 V103 -5044.682648592972
L61_103 V61 V103 -3.2042278092084887e-12
C61_103 V61 V103 -2.294253664590159e-19

R61_104 V61 V104 8921.03103942344
L61_104 V61 V104 1.2977647984807921e-11
C61_104 V61 V104 1.131122501050807e-19

R61_105 V61 V105 4745.019540578288
L61_105 V61 V105 -1.734485813390492e-12
C61_105 V61 V105 -3.034548722282705e-19

R61_106 V61 V106 1925.4661035086501
L61_106 V61 V106 1.3604112069993906e-12
C61_106 V61 V106 5.65183634408828e-19

R61_107 V61 V107 33088.02772222675
L61_107 V61 V107 1.4647677306779034e-12
C61_107 V61 V107 3.83865784339689e-19

R61_108 V61 V108 -7015.725202584801
L61_108 V61 V108 -1.550409383499916e-12
C61_108 V61 V108 -4.3054822667817083e-19

R61_109 V61 V109 -13998.80710012054
L61_109 V61 V109 -7.607559417201563e-12
C61_109 V61 V109 -8.232464365823149e-20

R61_110 V61 V110 -8510.631389760694
L61_110 V61 V110 -1.5830922050714281e-12
C61_110 V61 V110 -4.721920749458637e-19

R61_111 V61 V111 33627.28297817931
L61_111 V61 V111 -2.9843516457359583e-12
C61_111 V61 V111 -2.422922090773778e-19

R61_112 V61 V112 3742.997559689872
L61_112 V61 V112 1.1501277542135734e-12
C61_112 V61 V112 4.116901212285346e-19

R61_113 V61 V113 4139.146810287148
L61_113 V61 V113 2.849923832297183e-12
C61_113 V61 V113 1.5125815030352719e-19

R61_114 V61 V114 11780.35334447062
L61_114 V61 V114 2.3156169184775492e-12
C61_114 V61 V114 2.9744574785646834e-19

R61_115 V61 V115 -19379.540999282806
L61_115 V61 V115 2.8026842291761113e-12
C61_115 V61 V115 2.2918426318374687e-19

R61_116 V61 V116 -7059.189295383686
L61_116 V61 V116 -2.208022239487868e-12
C61_116 V61 V116 -2.4294766475492846e-19

R61_117 V61 V117 -2971.8522338809403
L61_117 V61 V117 -3.3051064352084357e-12
C61_117 V61 V117 -2.0538888027147994e-19

R61_118 V61 V118 6770.458978067701
L61_118 V61 V118 -2.5733484716685584e-12
C61_118 V61 V118 -1.969721918061799e-19

R61_119 V61 V119 6368.716433910063
L61_119 V61 V119 -2.3341890510723403e-12
C61_119 V61 V119 -3.116658057259371e-19

R61_120 V61 V120 -2741.9392398175864
L61_120 V61 V120 -2.4731716861093864e-11
C61_120 V61 V120 -1.4133862979011763e-19

R61_121 V61 V121 4886.8644986495165
L61_121 V61 V121 2.8808198086916307e-12
C61_121 V61 V121 3.7025494211265496e-20

R61_122 V61 V122 2793.7204602832044
L61_122 V61 V122 1.5845131820018412e-12
C61_122 V61 V122 4.23138636285162e-20

R61_123 V61 V123 -11813.191917876951
L61_123 V61 V123 1.9482770323798587e-11
C61_123 V61 V123 -4.823277066462678e-20

R61_124 V61 V124 -13744.749551784169
L61_124 V61 V124 -7.1399849723643e-12
C61_124 V61 V124 -1.145126969071201e-19

R61_125 V61 V125 -2393.385187067529
L61_125 V61 V125 -3.755112516326085e-12
C61_125 V61 V125 -1.7237560682676366e-20

R61_126 V61 V126 -4135.037870008213
L61_126 V61 V126 -2.182976773473523e-12
C61_126 V61 V126 6.156067604130666e-20

R61_127 V61 V127 -11105.514100153487
L61_127 V61 V127 2.7495360106532e-12
C61_127 V61 V127 -2.2876290882996406e-20

R61_128 V61 V128 -5837.847715991812
L61_128 V61 V128 4.03412407530926e-11
C61_128 V61 V128 -3.551754465069845e-20

R61_129 V61 V129 -5020.4364182443605
L61_129 V61 V129 1.0069264607642844e-10
C61_129 V61 V129 -9.995141256342132e-20

R61_130 V61 V130 -5540.418230156522
L61_130 V61 V130 -3.1494579682102275e-12
C61_130 V61 V130 -1.450840454675537e-19

R61_131 V61 V131 -9433.672406225422
L61_131 V61 V131 2.8886417600223904e-11
C61_131 V61 V131 1.1244954869720745e-19

R61_132 V61 V132 59904.94534889061
L61_132 V61 V132 -5.709433286190472e-12
C61_132 V61 V132 -3.1311339554817306e-20

R61_133 V61 V133 7858.5754753425135
L61_133 V61 V133 6.555428824490569e-12
C61_133 V61 V133 1.5629605312327123e-19

R61_134 V61 V134 3166.1743634798645
L61_134 V61 V134 -1.1760657771307163e-11
C61_134 V61 V134 1.1907009027749824e-20

R61_135 V61 V135 16047.021392776136
L61_135 V61 V135 4.532375885452672e-12
C61_135 V61 V135 -4.4072876549024554e-20

R61_136 V61 V136 -11120.627052620272
L61_136 V61 V136 -8.475095694608121e-10
C61_136 V61 V136 -5.598678522686187e-21

R61_137 V61 V137 -2088.231690824213
L61_137 V61 V137 -3.3272889099396137e-12
C61_137 V61 V137 -1.2191132101271765e-19

R61_138 V61 V138 -4175.298854187251
L61_138 V61 V138 -1.685638305174909e-12
C61_138 V61 V138 -1.101524864478674e-19

R61_139 V61 V139 -5172.336416297483
L61_139 V61 V139 1.7855725638775761e-12
C61_139 V61 V139 8.784546777351734e-20

R61_140 V61 V140 3774.5827372437375
L61_140 V61 V140 -3.748708718430317e-12
C61_140 V61 V140 -1.1816982494494049e-20

R61_141 V61 V141 -4853.39545413168
L61_141 V61 V141 -6.659239028005702e-12
C61_141 V61 V141 -2.518618660155372e-20

R61_142 V61 V142 3405.9214846703153
L61_142 V61 V142 -3.2458172336187906e-12
C61_142 V61 V142 -6.741890690674675e-20

R61_143 V61 V143 41014.93322360827
L61_143 V61 V143 -9.62653139921225e-12
C61_143 V61 V143 2.5408387390019365e-21

R61_144 V61 V144 4078.8194726711768
L61_144 V61 V144 4.249180610527954e-12
C61_144 V61 V144 2.8436228474215036e-20

R62_62 V62 0 -40.22964407522362
L62_62 V62 0 -2.964705352090374e-13
C62_62 V62 0 4.021955969858981e-18

R62_63 V62 V63 -3099.507165045764
L62_63 V62 V63 6.868063656569618e-12
C62_63 V62 V63 1.4301168545213922e-19

R62_64 V62 V64 9906.640802653348
L62_64 V62 V64 -5.650145312512394e-12
C62_64 V62 V64 -1.2993297169792512e-21

R62_65 V62 V65 209.853795054656
L62_65 V62 V65 2.8924023289761177e-12
C62_65 V62 V65 -1.8241894408335778e-19

R62_66 V62 V66 207.2060639161051
L62_66 V62 V66 -1.305424246198355e-11
C62_66 V62 V66 -2.9415007715864363e-19

R62_67 V62 V67 2993.10072202887
L62_67 V62 V67 -5.2245925741308725e-11
C62_67 V62 V67 -6.414078559295034e-20

R62_68 V62 V68 -19863.683035809325
L62_68 V62 V68 -2.5729453849078124e-11
C62_68 V62 V68 -3.00381749202179e-20

R62_69 V62 V69 -4879.230994511095
L62_69 V62 V69 1.970028025445663e-12
C62_69 V62 V69 4.999724271429926e-20

R62_70 V62 V70 -743.4977130344716
L62_70 V62 V70 -1.2550644537225241e-11
C62_70 V62 V70 -3.062221276329108e-20

R62_71 V62 V71 19699.379219356797
L62_71 V62 V71 -3.259022588238859e-11
C62_71 V62 V71 -7.121835874351716e-20

R62_72 V62 V72 -613.7352499171408
L62_72 V62 V72 7.783330265920339e-12
C62_72 V62 V72 5.197046954784657e-20

R62_73 V62 V73 -2398.570709766322
L62_73 V62 V73 5.889318600030598e-12
C62_73 V62 V73 -6.053945085730746e-20

R62_74 V62 V74 -1360.170308929042
L62_74 V62 V74 5.22549701978923e-12
C62_74 V62 V74 1.1371764032668291e-19

R62_75 V62 V75 1032.3134625613595
L62_75 V62 V75 1.527056895789405e-11
C62_75 V62 V75 -4.421704415397218e-20

R62_76 V62 V76 1160.501374054488
L62_76 V62 V76 1.604040231645674e-11
C62_76 V62 V76 -1.7046734779471922e-19

R62_77 V62 V77 2696.6863470903754
L62_77 V62 V77 8.628862231195919e-12
C62_77 V62 V77 -5.319831309644217e-20

R62_78 V62 V78 -10349.489151840708
L62_78 V62 V78 -4.503088745428257e-12
C62_78 V62 V78 -1.500770614002185e-19

R62_79 V62 V79 -3409.0764203200165
L62_79 V62 V79 4.797446132055573e-12
C62_79 V62 V79 2.98240524362009e-20

R62_80 V62 V80 -3833.0709869942816
L62_80 V62 V80 -2.1313936710827212e-11
C62_80 V62 V80 3.0213244420638397e-20

R62_81 V62 V81 -5691.141363273311
L62_81 V62 V81 -9.347523205066957e-12
C62_81 V62 V81 -5.423009707814342e-21

R62_82 V62 V82 12515.518033512502
L62_82 V62 V82 5.879366978907501e-12
C62_82 V62 V82 1.330095698543671e-19

R62_83 V62 V83 37008.55960306166
L62_83 V62 V83 5.618121093938179e-12
C62_83 V62 V83 5.3268451721031057e-20

R62_84 V62 V84 -11449.017054272033
L62_84 V62 V84 4.4478206423462895e-12
C62_84 V62 V84 3.441393100871566e-20

R62_85 V62 V85 -2603.3432320186853
L62_85 V62 V85 8.245924738069713e-12
C62_85 V62 V85 -5.6196473000269406e-21

R62_86 V62 V86 -4317.213951596985
L62_86 V62 V86 -8.298259008761416e-11
C62_86 V62 V86 -1.9081257459801612e-20

R62_87 V62 V87 15877.648908115689
L62_87 V62 V87 -1.1246277273041347e-10
C62_87 V62 V87 -3.962537541927067e-20

R62_88 V62 V88 -50483.85433264159
L62_88 V62 V88 -9.80982277622761e-12
C62_88 V62 V88 -3.859566107332875e-20

R62_89 V62 V89 4150.979906604029
L62_89 V62 V89 2.4359679573994527e-11
C62_89 V62 V89 6.309487367759098e-20

R62_90 V62 V90 -90952.60074331063
L62_90 V62 V90 -5.310782285628948e-12
C62_90 V62 V90 -3.800786359503176e-20

R62_91 V62 V91 -26751.904112669923
L62_91 V62 V91 5.7459343880356266e-12
C62_91 V62 V91 9.425002555886312e-20

R62_92 V62 V92 26086.095229830185
L62_92 V62 V92 7.01599005455149e-12
C62_92 V62 V92 3.6517525909963386e-20

R62_93 V62 V93 -1557.4085001163119
L62_93 V62 V93 1.3490814641466852e-10
C62_93 V62 V93 2.738347490239369e-20

R62_94 V62 V94 -3889.0761420570893
L62_94 V62 V94 -6.713406044718181e-12
C62_94 V62 V94 -6.003774580364858e-20

R62_95 V62 V95 19061.314782501868
L62_95 V62 V95 1.005222657859719e-11
C62_95 V62 V95 6.418629577938649e-20

R62_96 V62 V96 6432.024732329411
L62_96 V62 V96 1.0847532722716012e-11
C62_96 V62 V96 3.631105726290272e-20

R62_97 V62 V97 -2616.2332080907263
L62_97 V62 V97 -5.040641553725324e-12
C62_97 V62 V97 -4.661478573770968e-20

R62_98 V62 V98 -2682.334006957538
L62_98 V62 V98 1.4757741281591303e-11
C62_98 V62 V98 3.598889213603132e-20

R62_99 V62 V99 -7114.630216746748
L62_99 V62 V99 1.798770773276746e-11
C62_99 V62 V99 -2.6232057498837603e-21

R62_100 V62 V100 10692.988242021725
L62_100 V62 V100 -1.1866323243924469e-11
C62_100 V62 V100 -2.15501897589201e-20

R62_101 V62 V101 -4369.920738946273
L62_101 V62 V101 9.436015763420882e-12
C62_101 V62 V101 6.289405858408518e-20

R62_102 V62 V102 -6226.034168363732
L62_102 V62 V102 -3.971260618023756e-12
C62_102 V62 V102 -5.763611227234617e-20

R62_103 V62 V103 -5884.891177390809
L62_103 V62 V103 4.922847557365377e-12
C62_103 V62 V103 5.0308723416832885e-20

R62_104 V62 V104 16882.33284550064
L62_104 V62 V104 1.311964484278654e-11
C62_104 V62 V104 4.337237618997234e-20

R62_105 V62 V105 2837.0395541090293
L62_105 V62 V105 -1.1899026517255454e-11
C62_105 V62 V105 -4.8990201907691603e-20

R62_106 V62 V106 2892.328907418235
L62_106 V62 V106 1.169926232147009e-11
C62_106 V62 V106 8.494829060105516e-20

R62_107 V62 V107 -8575.032499597268
L62_107 V62 V107 -4.440454710258724e-12
C62_107 V62 V107 -5.967219823180788e-20

R62_108 V62 V108 12862.66346372047
L62_108 V62 V108 7.385352837056e-12
C62_108 V62 V108 3.9921678552866164e-20

R62_109 V62 V109 -16582.16415717109
L62_109 V62 V109 6.0012071488987754e-12
C62_109 V62 V109 5.219845449890218e-20

R62_110 V62 V110 18303.973318040717
L62_110 V62 V110 -4.9059136050853954e-12
C62_110 V62 V110 -1.081353441664748e-19

R62_111 V62 V111 8792.692352655575
L62_111 V62 V111 8.812215858698973e-12
C62_111 V62 V111 4.4676046292512115e-21

R62_112 V62 V112 8377.511464475427
L62_112 V62 V112 -1.1105694680114317e-11
C62_112 V62 V112 -7.541885827559666e-21

R62_113 V62 V113 4886.835977722011
L62_113 V62 V113 -2.8914775251237148e-11
C62_113 V62 V113 2.0493604347031855e-20

R62_114 V62 V114 -16696.59319751926
L62_114 V62 V114 3.5489880062176924e-11
C62_114 V62 V114 5.823739259218678e-20

R62_115 V62 V115 -10577.547660760843
L62_115 V62 V115 -8.047856557482526e-12
C62_115 V62 V115 -2.7919119454103414e-20

R62_116 V62 V116 -21330.478326079374
L62_116 V62 V116 1.3797022474756787e-11
C62_116 V62 V116 3.453439142479308e-20

R62_117 V62 V117 -3149.4683766656553
L62_117 V62 V117 8.440318061261356e-11
C62_117 V62 V117 -2.3521474054592073e-21

R62_118 V62 V118 3844.506773640056
L62_118 V62 V118 -6.242123706589942e-11
C62_118 V62 V118 -3.197609627891212e-20

R62_119 V62 V119 3303.608189827069
L62_119 V62 V119 -9.410068196890943e-11
C62_119 V62 V119 -3.37287048096425e-20

R62_120 V62 V120 -2423.522005977902
L62_120 V62 V120 -5.9053466003459725e-12
C62_120 V62 V120 -7.339749543028889e-21

R62_121 V62 V121 4959.641160410023
L62_121 V62 V121 3.513206369655768e-11
C62_121 V62 V121 4.88976006734917e-21

R62_122 V62 V122 4091.640532959347
L62_122 V62 V122 -6.418450718896534e-12
C62_122 V62 V122 2.3727916167820493e-20

R62_123 V62 V123 -7965.067675189132
L62_123 V62 V123 -1.2610572536969967e-11
C62_123 V62 V123 -1.6222927928661152e-20

R62_124 V62 V124 188707.18572923826
L62_124 V62 V124 -4.139390968417587e-11
C62_124 V62 V124 -3.3742864507689556e-20

R62_125 V62 V125 -2316.350332635058
L62_125 V62 V125 -1.8907190527477834e-11
C62_125 V62 V125 1.6762703617734536e-20

R62_126 V62 V126 -9039.416703606825
L62_126 V62 V126 3.740312059878422e-12
C62_126 V62 V126 3.864846354647731e-21

R62_127 V62 V127 -5547.523313411143
L62_127 V62 V127 -4.764266570572778e-12
C62_127 V62 V127 -1.856735935621772e-20

R62_128 V62 V128 -6117.957347957921
L62_128 V62 V128 -2.3428010786390752e-11
C62_128 V62 V128 -4.2909830007525896e-20

R62_129 V62 V129 -4987.274291455246
L62_129 V62 V129 -7.543113302261272e-12
C62_129 V62 V129 -4.5526197745160025e-20

R62_130 V62 V130 -29570.926272737288
L62_130 V62 V130 8.637345615464117e-12
C62_130 V62 V130 -2.9112244453089667e-20

R62_131 V62 V131 -10690.39435263134
L62_131 V62 V131 2.6354545179401608e-11
C62_131 V62 V131 -1.2491667470276345e-20

R62_132 V62 V132 22838.91469661195
L62_132 V62 V132 5.6209821455449935e-11
C62_132 V62 V132 -1.1761336547003917e-20

R62_133 V62 V133 12956.825766018193
L62_133 V62 V133 1.6698630644196237e-11
C62_133 V62 V133 3.2573116019309645e-20

R62_134 V62 V134 2695.1530498303127
L62_134 V62 V134 2.8898539662058058e-11
C62_134 V62 V134 -1.279483636981835e-20

R62_135 V62 V135 -45651.20659373127
L62_135 V62 V135 -7.783148775895698e-12
C62_135 V62 V135 1.6491987202843886e-21

R62_136 V62 V136 -11219.26173898423
L62_136 V62 V136 3.185538523042121e-11
C62_136 V62 V136 2.3896872454762788e-20

R62_137 V62 V137 -2493.494402880417
L62_137 V62 V137 -1.5194769502825253e-11
C62_137 V62 V137 -4.8909639898457444e-20

R62_138 V62 V138 -13589.28010114951
L62_138 V62 V138 4.439242856802847e-12
C62_138 V62 V138 -3.864312936351827e-20

R62_139 V62 V139 -2643.747489459638
L62_139 V62 V139 -3.7755961786439265e-12
C62_139 V62 V139 2.327760093763113e-20

R62_140 V62 V140 2834.7704793850667
L62_140 V62 V140 9.940700112535378e-12
C62_140 V62 V140 2.9903926062326027e-20

R62_141 V62 V141 -5890.202846152507
L62_141 V62 V141 1.6368684921634748e-11
C62_141 V62 V141 1.3871828400882124e-21

R62_142 V62 V142 2654.461169318482
L62_142 V62 V142 1.4489657624793098e-11
C62_142 V62 V142 1.4567113380998917e-21

R62_143 V62 V143 10045.410124783662
L62_143 V62 V143 8.98096057843081e-12
C62_143 V62 V143 3.124594013473797e-21

R62_144 V62 V144 5466.91807185404
L62_144 V62 V144 -2.1580443857595877e-11
C62_144 V62 V144 -2.9815143697325114e-20

R63_63 V63 0 -345.4979394607971
L63_63 V63 0 3.179362871149792e-13
C63_63 V63 0 2.4648102019359836e-18

R63_64 V63 V64 10133.720066734231
L63_64 V63 V64 1.4935555065565006e-11
C63_64 V63 V64 -1.943780059538278e-19

R63_65 V63 V65 2316.969987238833
L63_65 V63 V65 1.6205163387447406e-11
C63_65 V63 V65 -9.013854766308754e-20

R63_66 V63 V66 -3744.512050684619
L63_66 V63 V66 1.1208441781481186e-12
C63_66 V63 V66 2.693759032130753e-19

R63_67 V63 V67 784.3834830390522
L63_67 V63 V67 -2.364090791922303e-12
C63_67 V63 V67 -2.1504408621595935e-19

R63_68 V63 V68 6730.78764532412
L63_68 V63 V68 -4.069750816559617e-12
C63_68 V63 V68 -6.255683871470058e-20

R63_69 V63 V69 3643.61786826602
L63_69 V63 V69 -6.9355855704792675e-12
C63_69 V63 V69 1.9298801885730323e-20

R63_70 V63 V70 -3865.272994637878
L63_70 V63 V70 8.479631672392855e-12
C63_70 V63 V70 7.985831509564596e-20

R63_71 V63 V71 -923.0377337753526
L63_71 V63 V71 1.1296736757015357e-12
C63_71 V63 V71 2.627894790481126e-19

R63_72 V63 V72 3316.8799638607406
L63_72 V63 V72 -1.5054254751781282e-12
C63_72 V63 V72 -1.0511717391278717e-19

R63_73 V63 V73 3048.9027517328254
L63_73 V63 V73 -1.9561220369569203e-12
C63_73 V63 V73 -6.223692909304298e-20

R63_74 V63 V74 8295.142214322967
L63_74 V63 V74 -3.010141424757765e-12
C63_74 V63 V74 3.86116118891927e-21

R63_75 V63 V75 34514.88649786554
L63_75 V63 V75 1.4078704369936613e-11
C63_75 V63 V75 -1.9572521906934455e-19

R63_76 V63 V76 -417675.35710988304
L63_76 V63 V76 3.4633916310792e-12
C63_76 V63 V76 2.1316524240378454e-19

R63_77 V63 V77 -15945.744952729394
L63_77 V63 V77 5.2896657863032496e-11
C63_77 V63 V77 6.917757460671645e-20

R63_78 V63 V78 13133.409177851689
L63_78 V63 V78 4.118884927279417e-12
C63_78 V63 V78 2.234130927645602e-19

R63_79 V63 V79 15015.40353190186
L63_79 V63 V79 -9.130357436535695e-12
C63_79 V63 V79 1.1017262483050936e-19

R63_80 V63 V80 -7001.455214245947
L63_80 V63 V80 -3.1750141661846342e-12
C63_80 V63 V80 -2.2250087872357387e-19

R63_81 V63 V81 -86290.8581899798
L63_81 V63 V81 3.901906677029047e-12
C63_81 V63 V81 1.4652614827058358e-19

R63_82 V63 V82 -22144.409955692692
L63_82 V63 V82 -2.2979459642910435e-12
C63_82 V63 V82 -3.710591814526543e-19

R63_83 V63 V83 -3095.395618438707
L63_83 V63 V83 -4.488426030889407e-12
C63_83 V63 V83 -2.4254591602986753e-19

R63_84 V63 V84 7881.1255948588805
L63_84 V63 V84 -3.894428330787054e-12
C63_84 V63 V84 -1.2747894591665832e-20

R63_85 V63 V85 12077.797589722973
L63_85 V63 V85 4.108383402934611e-11
C63_85 V63 V85 1.243031776824416e-19

R63_86 V63 V86 5757.82665104932
L63_86 V63 V86 -2.7661776584190642e-11
C63_86 V63 V86 8.131604961433565e-20

R63_87 V63 V87 18316.66458791723
L63_87 V63 V87 2.965059080941959e-12
C63_87 V63 V87 2.2466702782073826e-19

R63_88 V63 V88 -840597.9767100606
L63_88 V63 V88 4.786334497828423e-12
C63_88 V63 V88 1.0779347575026602e-19

R63_89 V63 V89 -25706.861560043944
L63_89 V63 V89 -3.646213488150979e-12
C63_89 V63 V89 -1.8760298321018108e-19

R63_90 V63 V90 -12654.928760922014
L63_90 V63 V90 -9.620924061822555e-11
C63_90 V63 V90 -4.833026687712019e-20

R63_91 V63 V91 -10994.78851816067
L63_91 V63 V91 -2.8006148433970123e-12
C63_91 V63 V91 -2.844788545883008e-19

R63_92 V63 V92 -12369.936994059004
L63_92 V63 V92 -2.294324018457363e-12
C63_92 V63 V92 -2.757235315168861e-19

R63_93 V63 V93 -7613.874356081119
L63_93 V63 V93 1.0997267683964713e-11
C63_93 V63 V93 2.714249068378555e-20

R63_94 V63 V94 -15039.76684644155
L63_94 V63 V94 3.611290828227768e-12
C63_94 V63 V94 1.2397679005850235e-19

R63_95 V63 V95 -11037.009811823698
L63_95 V63 V95 -5.307756044644498e-12
C63_95 V63 V95 -1.5514799014034965e-19

R63_96 V63 V96 -30540.141465106895
L63_96 V63 V96 -2.9462669354631816e-12
C63_96 V63 V96 -2.107121692053646e-19

R63_97 V63 V97 20860.70081801448
L63_97 V63 V97 2.025782028370926e-11
C63_97 V63 V97 9.02932777823012e-20

R63_98 V63 V98 -12891.299815679717
L63_98 V63 V98 -2.483164475183664e-12
C63_98 V63 V98 -1.8721780877570572e-19

R63_99 V63 V99 -6785.063760994942
L63_99 V63 V99 1.4166614851585809e-11
C63_99 V63 V99 2.6163126906786006e-20

R63_100 V63 V100 54163.57296199228
L63_100 V63 V100 7.47240374457234e-12
C63_100 V63 V100 8.027465125611453e-20

R63_101 V63 V101 -7516.515088548409
L63_101 V63 V101 -2.5854487662905234e-12
C63_101 V63 V101 -2.5074747588500454e-19

R63_102 V63 V102 -5788.717961140246
L63_102 V63 V102 -2.97778565317898e-12
C63_102 V63 V102 -1.9309207441893958e-19

R63_103 V63 V103 8719.853828641208
L63_103 V63 V103 2.435231885009465e-11
C63_103 V63 V103 4.419752983106278e-20

R63_104 V63 V104 -15293.710069629145
L63_104 V63 V104 -5.07746336201392e-12
C63_104 V63 V104 -1.2774057079245565e-19

R63_105 V63 V105 15721.392281245164
L63_105 V63 V105 2.3602975587944103e-12
C63_105 V63 V105 2.779219080369082e-19

R63_106 V63 V106 -6615.277466967749
L63_106 V63 V106 -1.9870566819242804e-12
C63_106 V63 V106 -4.17874412732948e-19

R63_107 V63 V107 -8781.414646464933
L63_107 V63 V107 -4.311906046032681e-12
C63_107 V63 V107 -1.3321097996164535e-19

R63_108 V63 V108 8507.971834544564
L63_108 V63 V108 2.7109886155058107e-12
C63_108 V63 V108 2.4888021136158674e-19

R63_109 V63 V109 156529.09473211368
L63_109 V63 V109 -8.590613863277612e-12
C63_109 V63 V109 -5.874359077832765e-20

R63_110 V63 V110 4233.3916234314665
L63_110 V63 V110 1.793706421511623e-12
C63_110 V63 V110 3.97853959424275e-19

R63_111 V63 V111 127779.70050959144
L63_111 V63 V111 7.228404745552985e-12
C63_111 V63 V111 1.2238302888627303e-19

R63_112 V63 V112 287617.5886939377
L63_112 V63 V112 -2.1613524358792e-12
C63_112 V63 V112 -1.945873623702388e-19

R63_113 V63 V113 19719.568085452163
L63_113 V63 V113 -5.9506705876237314e-12
C63_113 V63 V113 -5.270294664997046e-20

R63_114 V63 V114 -27760.220755199694
L63_114 V63 V114 -3.5791346447627845e-12
C63_114 V63 V114 -2.1008342090205308e-19

R63_115 V63 V115 -12712.157093159092
L63_115 V63 V115 -9.310546083898272e-12
C63_115 V63 V115 -7.113332899697223e-20

R63_116 V63 V116 -406722.7831407133
L63_116 V63 V116 3.1291919010094514e-12
C63_116 V63 V116 1.6690239193980923e-19

R63_117 V63 V117 9236.385096544838
L63_117 V63 V117 5.5454419255269174e-12
C63_117 V63 V117 9.968817238867392e-20

R63_118 V63 V118 48544.21558200065
L63_118 V63 V118 3.896673877530454e-12
C63_118 V63 V118 1.4626601150261917e-19

R63_119 V63 V119 18098.741850330938
L63_119 V63 V119 3.0918115365908053e-12
C63_119 V63 V119 2.648848136283259e-19

R63_120 V63 V120 2572.2691908936654
L63_120 V63 V120 6.174037162952828e-12
C63_120 V63 V120 7.983039446469126e-20

R63_121 V63 V121 11508.833811269182
L63_121 V63 V121 -4.1243784622742465e-12
C63_121 V63 V121 -4.063505347787718e-20

R63_122 V63 V122 1763.1176778433717
L63_122 V63 V122 -3.521303584485976e-12
C63_122 V63 V122 -1.8606611063346266e-21

R63_123 V63 V123 7633.181855666088
L63_123 V63 V123 1.309803183506687e-10
C63_123 V63 V123 2.743113109963405e-20

R63_124 V63 V124 -46397.26206887012
L63_124 V63 V124 6.815647691756901e-12
C63_124 V63 V124 9.838483594371018e-20

R63_125 V63 V125 -93200.48022434229
L63_125 V63 V125 3.578887733188413e-12
C63_125 V63 V125 3.8925547523438635e-20

R63_126 V63 V126 -1326.6689109720583
L63_126 V63 V126 8.233160511210731e-12
C63_126 V63 V126 -4.9241138955284203e-20

R63_127 V63 V127 1941.6202519203405
L63_127 V63 V127 -1.6549700033057777e-11
C63_127 V63 V127 2.6872351016548048e-20

R63_128 V63 V128 20214.689030154233
L63_128 V63 V128 2.916668895766503e-10
C63_128 V63 V128 2.642818466144805e-20

R63_129 V63 V129 5476.642309961214
L63_129 V63 V129 1.2530541515801572e-11
C63_129 V63 V129 6.303917055945892e-20

R63_130 V63 V130 -7080.2465016082315
L63_130 V63 V130 7.401475034288892e-12
C63_130 V63 V130 8.322734048010116e-20

R63_131 V63 V131 -4621.475290307793
L63_131 V63 V131 -5.266692753613726e-11
C63_131 V63 V131 -4.125507666168087e-20

R63_132 V63 V132 -8570.13681595261
L63_132 V63 V132 9.98261608859442e-12
C63_132 V63 V132 2.76331926127764e-20

R63_133 V63 V133 -15868.068461928742
L63_133 V63 V133 -8.10289902341234e-12
C63_133 V63 V133 -1.2802654348144666e-19

R63_134 V63 V134 -16747.538020520464
L63_134 V63 V134 1.1872371121463567e-11
C63_134 V63 V134 1.5952328784503573e-20

R63_135 V63 V135 2410.6248042420675
L63_135 V63 V135 -1.4042180507621026e-11
C63_135 V63 V135 -5.940573562939102e-23

R63_136 V63 V136 -316127.53822767775
L63_136 V63 V136 -4.0865489652977174e-11
C63_136 V63 V136 -1.2678731731516439e-20

R63_137 V63 V137 -21413.548078994612
L63_137 V63 V137 4.342776883777394e-12
C63_137 V63 V137 8.17060066534606e-20

R63_138 V63 V138 -1798.0773538453575
L63_138 V63 V138 4.296201497416227e-12
C63_138 V63 V138 4.517581325589172e-20

R63_139 V63 V139 1698.2572894502414
L63_139 V63 V139 -6.8868025240250585e-12
C63_139 V63 V139 -2.0813347346149875e-20

R63_140 V63 V140 -5873.64835142908
L63_140 V63 V140 1.056740596637586e-11
C63_140 V63 V140 1.5302826515579898e-20

R63_141 V63 V141 -6172.830309725458
L63_141 V63 V141 1.527619954759298e-11
C63_141 V63 V141 -2.1351818907317212e-21

R63_142 V63 V142 -7023.831770288349
L63_142 V63 V142 9.477140352499862e-12
C63_142 V63 V142 4.618809582619364e-20

R63_143 V63 V143 -4549.908725373056
L63_143 V63 V143 2.8425153122730868e-11
C63_143 V63 V143 1.8401802757549232e-20

R63_144 V63 V144 5242.231820256171
L63_144 V63 V144 -1.1663079059487728e-11
C63_144 V63 V144 -1.449140313086255e-20

R64_64 V64 0 1202.1445198272393
L64_64 V64 0 1.3731385560481563e-13
C64_64 V64 0 1.6485194408255933e-18

R64_65 V64 V65 -5335.181707695749
L64_65 V64 V65 -2.621044422058755e-12
C64_65 V64 V65 8.007556413345344e-20

R64_66 V64 V66 -2181.1981930449865
L64_66 V64 V66 -1.00740291801354e-12
C64_66 V64 V66 -2.344180182931866e-19

R64_67 V64 V67 20445.13858152194
L64_67 V64 V67 -2.757893346507144e-12
C64_67 V64 V67 -1.3043551916556128e-19

R64_68 V64 V68 10657.736683931598
L64_68 V64 V68 -1.9397945736776084e-12
C64_68 V64 V68 -5.1809439286989664e-20

R64_69 V64 V69 7625.143350940367
L64_69 V64 V69 1.150060786934175e-11
C64_69 V64 V69 -4.8093563257569704e-20

R64_70 V64 V70 -10484.621596296249
L64_70 V64 V70 -5.05355082742633e-12
C64_70 V64 V70 -1.839088902698126e-19

R64_71 V64 V71 -2947.847716341745
L64_71 V64 V71 1.7769316177549762e-11
C64_71 V64 V71 -6.301154323954585e-20

R64_72 V64 V72 4816.483264696806
L64_72 V64 V72 3.3046012611848703e-12
C64_72 V64 V72 -2.5172080912767774e-20

R64_73 V64 V73 7013.705032079988
L64_73 V64 V73 -2.479669643702127e-12
C64_73 V64 V73 -1.1650943560476094e-19

R64_74 V64 V74 8626.721766044202
L64_74 V64 V74 2.4600643177753973e-11
C64_74 V64 V74 5.384205906594056e-20

R64_75 V64 V75 -18578.431197806774
L64_75 V64 V75 6.3979666043024856e-12
C64_75 V64 V75 1.4267369980474355e-19

R64_76 V64 V76 -14482.005685098717
L64_76 V64 V76 -2.110275656552073e-12
C64_76 V64 V76 -1.4088237324225537e-19

R64_77 V64 V77 -55905.32795739342
L64_77 V64 V77 8.952008106289505e-12
C64_77 V64 V77 1.0369807808783679e-19

R64_78 V64 V78 -13945.74154965952
L64_78 V64 V78 -2.160887159115897e-12
C64_78 V64 V78 -1.9256203006154427e-19

R64_79 V64 V79 196601.67072213124
L64_79 V64 V79 -3.1029660844494086e-12
C64_79 V64 V79 -1.7251565071026407e-19

R64_80 V64 V80 11311.417894677217
L64_80 V64 V80 1.4542939085347563e-12
C64_80 V64 V80 2.6572190774555423e-19

R64_81 V64 V81 -23518.976500332974
L64_81 V64 V81 -1.6593168505050776e-12
C64_81 V64 V81 -1.8378754416860929e-19

R64_82 V64 V82 6959.211626879186
L64_82 V64 V82 1.736764015436325e-12
C64_82 V64 V82 3.058519384583487e-19

R64_83 V64 V83 36783.2888966182
L64_83 V64 V83 1.159407621331687e-12
C64_83 V64 V83 3.3943235581676967e-19

R64_84 V64 V84 19568.83627399314
L64_84 V64 V84 -7.425012676861285e-11
C64_84 V64 V84 -4.879820057096681e-20

R64_85 V64 V85 -35211.518274163274
L64_85 V64 V85 -2.1458708259412347e-12
C64_85 V64 V85 -2.582894651504798e-19

R64_86 V64 V86 81683.78002906972
L64_86 V64 V86 -2.7635448418131194e-12
C64_86 V64 V86 -1.7153041742986049e-19

R64_87 V64 V87 -9707.151001725562
L64_87 V64 V87 -2.0247384016919608e-12
C64_87 V64 V87 -1.9464875144549107e-19

R64_88 V64 V88 -28623.815087150273
L64_88 V64 V88 -5.712476648662531e-12
C64_88 V64 V88 -3.4493725488219065e-20

R64_89 V64 V89 17159.226568622515
L64_89 V64 V89 3.0746794251864174e-12
C64_89 V64 V89 1.7701508014369162e-19

R64_90 V64 V90 27048.845610927146
L64_90 V64 V90 2.5678204763797786e-12
C64_90 V64 V90 2.0468602742626946e-19

R64_91 V64 V91 9848.935683749709
L64_91 V64 V91 1.904879446444246e-12
C64_91 V64 V91 2.833347031467895e-19

R64_92 V64 V92 10788.598336000712
L64_92 V64 V92 1.3085232125353797e-12
C64_92 V64 V92 2.4270939135342747e-19

R64_93 V64 V93 47816.36476520184
L64_93 V64 V93 -5.682387652041095e-12
C64_93 V64 V93 -4.1368233660527976e-20

R64_94 V64 V94 -22541.00940327585
L64_94 V64 V94 -2.353026906308917e-12
C64_94 V64 V94 -1.2812561050417045e-19

R64_95 V64 V95 18015.04229600981
L64_95 V64 V95 3.1611985199780393e-12
C64_95 V64 V95 1.6715771894747007e-19

R64_96 V64 V96 17745.934293489147
L64_96 V64 V96 1.367170785104429e-12
C64_96 V64 V96 2.082910507156165e-19

R64_97 V64 V97 47405.303836526946
L64_97 V64 V97 -1.467093117805256e-11
C64_97 V64 V97 3.5686687505011924e-22

R64_98 V64 V98 9477.779631972047
L64_98 V64 V98 1.5851186791770521e-12
C64_98 V64 V98 2.2743208255147274e-19

R64_99 V64 V99 -33178.56530645424
L64_99 V64 V99 -4.4169230522770476e-12
C64_99 V64 V99 -6.100694999237054e-20

R64_100 V64 V100 -30646.620142140287
L64_100 V64 V100 -4.671503614401311e-12
C64_100 V64 V100 -1.1819360662923706e-20

R64_101 V64 V101 10429.303865982029
L64_101 V64 V101 1.864579546919729e-12
C64_101 V64 V101 2.277338630945923e-19

R64_102 V64 V102 5134.613783421513
L64_102 V64 V102 1.095316084999078e-12
C64_102 V64 V102 5.078530612218456e-19

R64_103 V64 V103 -21959.621823543905
L64_103 V64 V103 -2.4676089758283907e-12
C64_103 V64 V103 -2.3448723014006435e-19

R64_104 V64 V104 30547.273692799303
L64_104 V64 V104 2.179111605607417e-12
C64_104 V64 V104 1.6272014795065448e-19

R64_105 V64 V105 -7447.572022558151
L64_105 V64 V105 -1.2355010513490449e-12
C64_105 V64 V105 -3.367328455541791e-19

R64_106 V64 V106 6220.500426843354
L64_106 V64 V106 9.437832416250303e-13
C64_106 V64 V106 5.430800382254702e-19

R64_107 V64 V107 7566.182415591393
L64_107 V64 V107 1.3645803176569947e-12
C64_107 V64 V107 3.8903931289338234e-19

R64_108 V64 V108 -6356.582506724402
L64_108 V64 V108 -1.180190876620311e-12
C64_108 V64 V108 -3.890357047916448e-19

R64_109 V64 V109 -30524.12802047816
L64_109 V64 V109 7.946374320631502e-12
C64_109 V64 V109 -6.146901375137885e-20

R64_110 V64 V110 -8819.015023957092
L64_110 V64 V110 -1.19291393928736e-12
C64_110 V64 V110 -4.317712990230769e-19

R64_111 V64 V111 -10380.654475872465
L64_111 V64 V111 -1.9672057920354196e-12
C64_111 V64 V111 -2.233648145037334e-19

R64_112 V64 V112 6897.986243573865
L64_112 V64 V112 1.2619054520421264e-12
C64_112 V64 V112 3.086417861679931e-19

R64_113 V64 V113 22639.75949956842
L64_113 V64 V113 3.772611633882191e-12
C64_113 V64 V113 1.626655462481098e-19

R64_114 V64 V114 9210.678037871488
L64_114 V64 V114 2.1872634099813446e-12
C64_114 V64 V114 1.93272659895037e-19

R64_115 V64 V115 9918.796843904833
L64_115 V64 V115 2.563283001194949e-12
C64_115 V64 V115 2.0722998921504168e-19

R64_116 V64 V116 -8909.768241127105
L64_116 V64 V116 -1.6677264072929083e-12
C64_116 V64 V116 -2.539563176775879e-19

R64_117 V64 V117 -23492.131747650445
L64_117 V64 V117 -3.5154345127205392e-12
C64_117 V64 V117 -2.269988676202014e-19

R64_118 V64 V118 -12929.56788760478
L64_118 V64 V118 -2.49483609433153e-12
C64_118 V64 V118 -2.0370447129820466e-19

R64_119 V64 V119 -6855.494246874871
L64_119 V64 V119 -1.6539938729141416e-12
C64_119 V64 V119 -2.3531219937385074e-19

R64_120 V64 V120 21836.681355629236
L64_120 V64 V120 -3.743089638324677e-11
C64_120 V64 V120 -7.780326733152154e-20

R64_121 V64 V121 98418.87324404556
L64_121 V64 V121 4.67765987845129e-12
C64_121 V64 V121 5.008179757553157e-20

R64_122 V64 V122 13452.080805519641
L64_122 V64 V122 2.317400709003556e-12
C64_122 V64 V122 2.009600161911918e-20

R64_123 V64 V123 25298.592605295264
L64_123 V64 V123 9.813724491239716e-11
C64_123 V64 V123 -3.000069262020106e-20

R64_124 V64 V124 -997466.6664239718
L64_124 V64 V124 -4.072673715833382e-12
C64_124 V64 V124 -6.331410836670858e-20

R64_125 V64 V125 39411.59543715092
L64_125 V64 V125 -5.224160311069749e-12
C64_125 V64 V125 -6.548698095230574e-20

R64_126 V64 V126 -11353.755326437871
L64_126 V64 V126 -2.717222929558956e-12
C64_126 V64 V126 5.354761551602195e-20

R64_127 V64 V127 10974.557903737461
L64_127 V64 V127 2.7951756624092356e-12
C64_127 V64 V127 2.3689680954626543e-20

R64_128 V64 V128 -57797.69908416357
L64_128 V64 V128 -5.162487030331974e-11
C64_128 V64 V128 -6.78327754353418e-20

R64_129 V64 V129 15053.629886341574
L64_129 V64 V129 8.457594041648702e-11
C64_129 V64 V129 -3.3812397152812756e-20

R64_130 V64 V130 -9316.637199273884
L64_130 V64 V130 -2.9482385515907123e-12
C64_130 V64 V130 -1.8713474708808197e-19

R64_131 V64 V131 -49548.89795094815
L64_131 V64 V131 1.4991027072364878e-11
C64_131 V64 V131 6.483945621996014e-20

R64_132 V64 V132 -21450.578676858226
L64_132 V64 V132 -4.2685443247645225e-12
C64_132 V64 V132 -6.427386641601781e-20

R64_133 V64 V133 24476.14360203503
L64_133 V64 V133 3.0634367763331044e-12
C64_133 V64 V133 1.9435053464228652e-19

R64_134 V64 V134 -45177.158039469476
L64_134 V64 V134 -1.3761111543776118e-11
C64_134 V64 V134 6.532122471838389e-21

R64_135 V64 V135 23479.67935657973
L64_135 V64 V135 5.965385355084346e-12
C64_135 V64 V135 -4.2608800020560106e-20

R64_136 V64 V136 74665.60389132994
L64_136 V64 V136 8.199710077122755e-12
C64_136 V64 V136 8.437935152323613e-20

R64_137 V64 V137 107362.3974204522
L64_137 V64 V137 -4.540021486803235e-12
C64_137 V64 V137 -6.285882124222803e-20

R64_138 V64 V138 -8183.994827349577
L64_138 V64 V138 -2.8402131075108297e-12
C64_138 V64 V138 2.1854522885306527e-20

R64_139 V64 V139 7334.466509704868
L64_139 V64 V139 1.7897148032359091e-12
C64_139 V64 V139 8.391530637608333e-20

R64_140 V64 V140 -12209.396137110363
L64_140 V64 V140 -4.992483333562564e-12
C64_140 V64 V140 -1.492771978458993e-20

R64_141 V64 V141 50699.056704451985
L64_141 V64 V141 -1.1536965103357545e-11
C64_141 V64 V141 2.679152036596709e-20

R64_142 V64 V142 -9145.920469404695
L64_142 V64 V142 -4.8849398222115025e-12
C64_142 V64 V142 -4.6520003243447065e-20

R64_143 V64 V143 -17198.969001635745
L64_143 V64 V143 -7.164741912808552e-12
C64_143 V64 V143 -1.0409695761198832e-20

R64_144 V64 V144 58768.0294522255
L64_144 V64 V144 6.835290230808188e-12
C64_144 V64 V144 -6.7051018199127495e-21

R65_65 V65 0 23.14687911273628
L65_65 V65 0 2.6521992285775858e-14
C65_65 V65 0 1.5515709561072032e-18

R65_66 V65 V66 -158.47013432727456
L65_66 V65 V66 -1.9846642552249524e-13
C65_66 V65 V66 -4.922623984630233e-20

R65_67 V65 V67 -835.240183479372
L65_67 V65 V67 -9.809847449730177e-13
C65_67 V65 V67 -5.168225306287954e-20

R65_68 V65 V68 -1708.8988178233774
L65_68 V65 V68 -1.7371113792477191e-12
C65_68 V65 V68 -2.47563658435855e-20

R65_69 V65 V69 1100.426296578495
L65_69 V65 V69 1.058718760511203e-12
C65_69 V65 V69 2.4339954413002257e-20

R65_70 V65 V70 670.4272772185968
L65_70 V65 V70 8.480382485384479e-13
C65_70 V65 V70 6.537055917585627e-20

R65_71 V65 V71 2992.7290719742646
L65_71 V65 V71 1.2947118554982387e-12
C65_71 V65 V71 7.690069363104528e-20

R65_72 V65 V72 526.5919929670692
L65_72 V65 V72 5.285463727053384e-13
C65_72 V65 V72 1.8880221652851498e-20

R65_73 V65 V73 5858.064363421343
L65_73 V65 V73 4.107984164893579e-12
C65_73 V65 V73 -1.0688646727036461e-20

R65_74 V65 V74 991.4843211186452
L65_74 V65 V74 9.190880385847756e-13
C65_74 V65 V74 1.2578946006155395e-20

R65_75 V65 V75 -831.5523219737419
L65_75 V65 V75 -7.021646650127139e-13
C65_75 V65 V75 -1.4043357134248154e-19

R65_76 V65 V76 -935.6615608569551
L65_76 V65 V76 -6.626195565372339e-13
C65_76 V65 V76 1.417805216976838e-22

R65_77 V65 V77 -2642.309586180004
L65_77 V65 V77 -1.587376356525156e-12
C65_77 V65 V77 -4.236200847803311e-20

R65_78 V65 V78 -45359.11304408757
L65_78 V65 V78 -2.2286949662645877e-12
C65_78 V65 V78 1.6012113471452267e-20

R65_79 V65 V79 2678.515376735831
L65_79 V65 V79 1.9496196555095533e-12
C65_79 V65 V79 8.561576418305755e-20

R65_80 V65 V80 2890.3232319158137
L65_80 V65 V80 2.6862876847771352e-12
C65_80 V65 V80 -6.768982739355845e-20

R65_81 V65 V81 5326.951582396464
L65_81 V65 V81 2.404405340705522e-12
C65_81 V65 V81 7.420302997081694e-20

R65_82 V65 V82 213622.9627661782
L65_82 V65 V82 -1.8826445602744907e-12
C65_82 V65 V82 -1.1165357380804602e-19

R65_83 V65 V83 47145.70076542325
L65_83 V65 V83 -1.4396370842683877e-11
C65_83 V65 V83 -1.4814515739759823e-19

R65_84 V65 V84 114375.8512990239
L65_84 V65 V84 3.113196947998449e-12
C65_84 V65 V84 -1.0463640248141351e-20

R65_85 V65 V85 2497.0168383589394
L65_85 V65 V85 1.980380373956709e-12
C65_85 V65 V85 6.187810273666247e-20

R65_86 V65 V86 6654.486106241007
L65_86 V65 V86 7.482184235368982e-12
C65_86 V65 V86 3.234652335478287e-20

R65_87 V65 V87 -18820.967142059686
L65_87 V65 V87 -8.997021303347677e-10
C65_87 V65 V87 4.008462528799112e-20

R65_88 V65 V88 14097.865741910284
L65_88 V65 V88 -8.498583039324269e-12
C65_88 V65 V88 6.696372451735012e-21

R65_89 V65 V89 -4517.533417804272
L65_89 V65 V89 -7.644928068049551e-12
C65_89 V65 V89 -1.5558400056836652e-20

R65_90 V65 V90 114284.4363879082
L65_90 V65 V90 -5.65773314403571e-12
C65_90 V65 V90 -7.786467096653629e-20

R65_91 V65 V91 14439.01966426528
L65_91 V65 V91 -3.5904117673007362e-12
C65_91 V65 V91 -1.198250333181192e-19

R65_92 V65 V92 -17721.84886075795
L65_92 V65 V92 -5.486598235854324e-12
C65_92 V65 V92 -1.1014921618791261e-19

R65_93 V65 V93 1089.189710188033
L65_93 V65 V93 7.733432585620998e-12
C65_93 V65 V93 5.617878128471257e-20

R65_94 V65 V94 2870.419866274626
L65_94 V65 V94 1.1190095473495673e-11
C65_94 V65 V94 3.977521476417693e-20

R65_95 V65 V95 -50734.198443905014
L65_95 V65 V95 -6.334878179208542e-12
C65_95 V65 V95 -5.467164256783182e-20

R65_96 V65 V96 -3749.419460293381
L65_96 V65 V96 -8.200267139831597e-12
C65_96 V65 V96 -7.837410637628465e-20

R65_97 V65 V97 2251.962478842669
L65_97 V65 V97 8.934977588639381e-12
C65_97 V65 V97 1.920172308209985e-20

R65_98 V65 V98 1892.5893449089058
L65_98 V65 V98 3.463146485288306e-11
C65_98 V65 V98 -5.646847328611295e-20

R65_99 V65 V99 3812.2821729481566
L65_99 V65 V99 1.2717564896597694e-11
C65_99 V65 V99 1.370552186750687e-20

R65_100 V65 V100 -8789.043141257218
L65_100 V65 V100 4.184631128327759e-11
C65_100 V65 V100 1.9727976564915675e-20

R65_101 V65 V101 2763.9665512212314
L65_101 V65 V101 -4.468123576208221e-11
C65_101 V65 V101 -2.8855115738583656e-20

R65_102 V65 V102 3886.2595920606122
L65_102 V65 V102 -2.737059647933184e-12
C65_102 V65 V102 -1.7886142039054315e-19

R65_103 V65 V103 3832.6800298777666
L65_103 V65 V103 5.948158771153927e-12
C65_103 V65 V103 5.683018501643263e-20

R65_104 V65 V104 -10885.428033653889
L65_104 V65 V104 -2.109884536413573e-11
C65_104 V65 V104 -5.731373845585395e-20

R65_105 V65 V105 -2475.6074755232553
L65_105 V65 V105 4.253724834284461e-12
C65_105 V65 V105 1.4092602491007543e-19

R65_106 V65 V106 -1944.7890455185147
L65_106 V65 V106 -1.9787069919289048e-12
C65_106 V65 V106 -1.8140352800598533e-19

R65_107 V65 V107 14582.13068844468
L65_107 V65 V107 -3.5920353665106376e-12
C65_107 V65 V107 -1.5105259811723308e-19

R65_108 V65 V108 -20957.377943912554
L65_108 V65 V108 4.983325585396559e-12
C65_108 V65 V108 9.939224978883057e-20

R65_109 V65 V109 17143.07981029167
L65_109 V65 V109 8.582961115467555e-12
C65_109 V65 V109 1.0800563103018776e-21

R65_110 V65 V110 -32979.014284766614
L65_110 V65 V110 4.61139830841288e-12
C65_110 V65 V110 1.45004392764567e-19

R65_111 V65 V111 -7775.400796945257
L65_111 V65 V111 3.496191680758376e-12
C65_111 V65 V111 8.309681997676367e-20

R65_112 V65 V112 -7084.1138059009145
L65_112 V65 V112 -2.162083608985387e-11
C65_112 V65 V112 -6.105470792164605e-20

R65_113 V65 V113 -3806.888474558475
L65_113 V65 V113 -1.070526319760918e-11
C65_113 V65 V113 -3.978439518778737e-20

R65_114 V65 V114 15503.233942963665
L65_114 V65 V114 -7.834976562402999e-12
C65_114 V65 V114 -6.100679022581736e-20

R65_115 V65 V115 6277.82909610506
L65_115 V65 V115 -4.76804879550943e-12
C65_115 V65 V115 -7.392133122652199e-20

R65_116 V65 V116 13566.409088281065
L65_116 V65 V116 7.830528160834567e-12
C65_116 V65 V116 7.010388639253948e-20

R65_117 V65 V117 2672.2262690385246
L65_117 V65 V117 1.0854722098403128e-11
C65_117 V65 V117 6.125198574690808e-20

R65_118 V65 V118 -3211.6457765495975
L65_118 V65 V118 7.399296225586009e-12
C65_118 V65 V118 7.880321019096684e-20

R65_119 V65 V119 -2569.4677719547053
L65_119 V65 V119 3.586844782158727e-12
C65_119 V65 V119 9.97307324701685e-20

R65_120 V65 V120 1954.7518515038048
L65_120 V65 V120 -5.0828131966823325e-12
C65_120 V65 V120 2.2283309178108925e-20

R65_121 V65 V121 -3397.8328371387965
L65_121 V65 V121 1.0017724111907696e-11
C65_121 V65 V121 -4.3190451770092724e-20

R65_122 V65 V122 -2586.1853909926604
L65_122 V65 V122 3.355384211835253e-11
C65_122 V65 V122 1.4119647064589073e-20

R65_123 V65 V123 6508.664745036054
L65_123 V65 V123 8.540120970628441e-12
C65_123 V65 V123 4.0601947837035375e-20

R65_124 V65 V124 14487.20535626662
L65_124 V65 V124 8.768007870413848e-12
C65_124 V65 V124 3.6027368869754274e-20

R65_125 V65 V125 1641.7869812163397
L65_125 V65 V125 -4.3790394905134565e-12
C65_125 V65 V125 1.836774713135286e-20

R65_126 V65 V126 4002.8015888831887
L65_126 V65 V126 6.867926440980119e-12
C65_126 V65 V126 -1.6229218222911332e-20

R65_127 V65 V127 5306.039498877778
L65_127 V65 V127 -4.6063750953804204e-12
C65_127 V65 V127 -2.0860071229691163e-21

R65_128 V65 V128 4830.042028825698
L65_128 V65 V128 5.420720607241452e-11
C65_128 V65 V128 2.3943496005469314e-20

R65_129 V65 V129 3529.0069137843093
L65_129 V65 V129 -5.7487543243843956e-11
C65_129 V65 V129 2.1738361232855024e-20

R65_130 V65 V130 10275.214936739092
L65_130 V65 V130 1.5707983137444588e-11
C65_130 V65 V130 4.8468962561085835e-20

R65_131 V65 V131 8467.426557083565
L65_131 V65 V131 -1.2148817239826912e-11
C65_131 V65 V131 -3.521696450969654e-20

R65_132 V65 V132 -21761.60855363249
L65_132 V65 V132 2.0345274196240527e-11
C65_132 V65 V132 2.534785114462916e-20

R65_133 V65 V133 -8006.348877502798
L65_133 V65 V133 -4.398045858241013e-12
C65_133 V65 V133 -6.664395149096124e-20

R65_134 V65 V134 -2167.02114526033
L65_134 V65 V134 -1.2405729078042872e-11
C65_134 V65 V134 -1.5685267036249176e-21

R65_135 V65 V135 -23824.181380845497
L65_135 V65 V135 -1.0412077914117392e-11
C65_135 V65 V135 1.484011580036218e-20

R65_136 V65 V136 9059.132329790526
L65_136 V65 V136 -1.5639712587025885e-11
C65_136 V65 V136 -3.431360208701641e-20

R65_137 V65 V137 1644.7373960972639
L65_137 V65 V137 -1.0506119008273628e-11
C65_137 V65 V137 1.1914168188628904e-22

R65_138 V65 V138 6534.745053612745
L65_138 V65 V138 1.2576117302335825e-11
C65_138 V65 V138 1.0743197244128868e-22

R65_139 V65 V139 2418.3381349070323
L65_139 V65 V139 -3.82466070727448e-12
C65_139 V65 V139 -1.4455579398849332e-20

R65_140 V65 V140 -2334.830286356742
L65_140 V65 V140 1.24660107449694e-10
C65_140 V65 V140 5.687935643376447e-21

R65_141 V65 V141 3678.048389880202
L65_141 V65 V141 6.479998911269103e-11
C65_141 V65 V141 -1.539295568806097e-20

R65_142 V65 V142 -2081.3202170857826
L65_142 V65 V142 9.461046981820933e-12
C65_142 V65 V142 5.237117168932757e-20

R65_143 V65 V143 -11187.489442573178
L65_143 V65 V143 1.1871580406099594e-11
C65_143 V65 V143 3.659510268366489e-21

R65_144 V65 V144 -3221.562791285255
L65_144 V65 V144 -2.2872233284563867e-11
C65_144 V65 V144 -1.3171379638070528e-20

R66_66 V66 0 25.28694752691845
L66_66 V66 0 2.7971024645330376e-14
C66_66 V66 0 1.764699935442787e-18

R66_67 V66 V67 -6095.6462274792875
L66_67 V66 V67 5.0716216247829134e-12
C66_67 V66 V67 4.637610692262515e-20

R66_68 V66 V68 -2825.8879836818464
L66_68 V66 V68 -5.469613135074337e-12
C66_68 V66 V68 2.5390604127460392e-21

R66_69 V66 V69 957.027881812557
L66_69 V66 V69 5.66598119599531e-13
C66_69 V66 V69 1.8085041532491073e-20

R66_70 V66 V70 888.4355185758587
L66_70 V66 V70 5.088509255846901e-12
C66_70 V66 V70 -3.169670247239856e-19

R66_71 V66 V71 -2751.475926993962
L66_71 V66 V71 -1.3373923856792624e-12
C66_71 V66 V71 -2.2806026735870387e-19

R66_72 V66 V72 510.4888510740271
L66_72 V66 V72 4.075802052638757e-13
C66_72 V66 V72 4.3128805001239033e-20

R66_73 V66 V73 2696.450305157113
L66_73 V66 V73 1.3714742243683113e-12
C66_73 V66 V73 -6.88248207878804e-20

R66_74 V66 V74 870.4051154233565
L66_74 V66 V74 5.654916121215519e-13
C66_74 V66 V74 8.104746814865664e-20

R66_75 V66 V75 -1026.155090129512
L66_75 V66 V75 -1.4325146015519315e-12
C66_75 V66 V75 2.4044793367973604e-19

R66_76 V66 V76 -863.8849642941503
L66_76 V66 V76 -3.9097551346292613e-13
C66_76 V66 V76 -4.608130324887103e-19

R66_77 V66 V77 -2967.0469435839314
L66_77 V66 V77 -1.6584037033531925e-12
C66_77 V66 V77 8.55662535153224e-21

R66_78 V66 V78 30890.432043425244
L66_78 V66 V78 -1.0167439684489495e-12
C66_78 V66 V78 -3.0115593662125866e-19

R66_79 V66 V79 3576.384995614652
L66_79 V66 V79 1.7495708049928795e-11
C66_79 V66 V79 -2.7389153610147578e-19

R66_80 V66 V80 1964.6884093990452
L66_80 V66 V80 7.16827851182846e-13
C66_80 V66 V80 5.1211531959688e-19

R66_81 V66 V81 19629.21956163173
L66_81 V66 V81 -3.4816174737888525e-12
C66_81 V66 V81 -2.5779720672547873e-19

R66_82 V66 V82 4998.059808347108
L66_82 V66 V82 1.148333448278392e-12
C66_82 V66 V82 5.652629936256333e-19

R66_83 V66 V83 10895.286469734388
L66_83 V66 V83 8.855658685636689e-13
C66_83 V66 V83 4.868837675452535e-19

R66_84 V66 V84 -19161.1784686709
L66_84 V66 V84 3.3860280452433015e-12
C66_84 V66 V84 -1.4278034096871573e-19

R66_85 V66 V85 4853.5602543275345
L66_85 V66 V85 -3.764847477461479e-12
C66_85 V66 V85 -4.0752850297762338e-19

R66_86 V66 V86 5372.248494423528
L66_86 V66 V86 -9.718114178085368e-12
C66_86 V66 V86 -2.042147410933913e-19

R66_87 V66 V87 -4853.631938605243
L66_87 V66 V87 -1.0233908519962058e-12
C66_87 V66 V87 -4.410931257030582e-19

R66_88 V66 V88 17778.464898635157
L66_88 V66 V88 -2.0222638808231796e-12
C66_88 V66 V88 -1.26131865762741e-19

R66_89 V66 V89 -121344.46208723086
L66_89 V66 V89 1.7912873984043438e-12
C66_89 V66 V89 3.7714453151539105e-19

R66_90 V66 V90 9066.229590138932
L66_90 V66 V90 2.035514737938818e-12
C66_90 V66 V90 3.0578604589737214e-19

R66_91 V66 V91 5110.428921621083
L66_91 V66 V91 1.1293387612502089e-12
C66_91 V66 V91 4.273614754773945e-19

R66_92 V66 V92 7523.8229898764175
L66_92 V66 V92 9.795924984152957e-13
C66_92 V66 V92 4.56896935180355e-19

R66_93 V66 V93 1174.5125156073818
L66_93 V66 V93 -4.716220047797124e-12
C66_93 V66 V93 -2.629688227797088e-20

R66_94 V66 V94 3718.1045882793633
L66_94 V66 V94 -1.8447922823600834e-12
C66_94 V66 V94 -1.6002058569195859e-19

R66_95 V66 V95 24173.545578968442
L66_95 V66 V95 2.0281099464989265e-12
C66_95 V66 V95 2.7814566317829935e-19

R66_96 V66 V96 -13483.955274484424
L66_96 V66 V96 1.247577224275981e-12
C66_96 V66 V96 3.6936176998702794e-19

R66_97 V66 V97 2289.35353867684
L66_97 V66 V97 6.708284893819555e-12
C66_97 V66 V97 -6.878266474358102e-21

R66_98 V66 V98 1794.660631704662
L66_98 V66 V98 8.383100121377445e-13
C66_98 V66 V98 3.9209381838725445e-19

R66_99 V66 V99 4929.3645637127
L66_99 V66 V99 -3.1200532927115655e-12
C66_99 V66 V99 -7.789305522442833e-20

R66_100 V66 V100 -7711.681584612325
L66_100 V66 V100 -3.0994435932561952e-12
C66_100 V66 V100 -1.0753092646942275e-19

R66_101 V66 V101 1775.7029179736378
L66_101 V66 V101 9.982664014257727e-13
C66_101 V66 V101 4.913647444904323e-19

R66_102 V66 V102 1769.179328083265
L66_102 V66 V102 5.921506938071704e-13
C66_102 V66 V102 8.64856906455514e-19

R66_103 V66 V103 9437.055584574273
L66_103 V66 V103 -1.7262767614831999e-12
C66_103 V66 V103 -3.9417299319806324e-19

R66_104 V66 V104 1105442.8395741314
L66_104 V66 V104 2.990012107831197e-12
C66_104 V66 V104 2.236083365570369e-19

R66_105 V66 V105 -1676.348778476842
L66_105 V66 V105 -7.688297027257351e-13
C66_105 V66 V105 -5.492486919330926e-19

R66_106 V66 V106 -36255.37464226713
L66_106 V66 V106 6.036439871402368e-13
C66_106 V66 V106 9.317038635194304e-19

R66_107 V66 V107 2843.6703298246925
L66_107 V66 V107 8.046264795727996e-13
C66_107 V66 V107 6.055711931922487e-19

R66_108 V66 V108 -1996.939611857285
L66_108 V66 V108 -7.274980324983168e-13
C66_108 V66 V108 -7.287234392920107e-19

R66_109 V66 V109 -14358.223207058742
L66_109 V66 V109 -1.5016424154854632e-11
C66_109 V66 V109 -1.0187260061186256e-19

R66_110 V66 V110 -2279.741464734413
L66_110 V66 V110 -6.857332623810092e-13
C66_110 V66 V110 -7.363728834283412e-19

R66_111 V66 V111 -4696.068226946719
L66_111 V66 V111 -1.3516459607115657e-12
C66_111 V66 V111 -3.8788100423642333e-19

R66_112 V66 V112 55754.781061988084
L66_112 V66 V112 5.932254287878768e-13
C66_112 V66 V112 6.256001001454678e-19

R66_113 V66 V113 -4975.180011947192
L66_113 V66 V113 1.5199139737581212e-12
C66_113 V66 V113 2.4515242302774144e-19

R66_114 V66 V114 4559.812930069519
L66_114 V66 V114 1.0525450633649995e-12
C66_114 V66 V114 4.339137527459037e-19

R66_115 V66 V115 5051.786356168948
L66_115 V66 V115 1.737687327562044e-12
C66_115 V66 V115 3.2056831081186045e-19

R66_116 V66 V116 -8658.45249441958
L66_116 V66 V116 -1.0264644526305289e-12
C66_116 V66 V116 -4.174565970228868e-19

R66_117 V66 V117 6290.327772534267
L66_117 V66 V117 -1.7755819641758684e-12
C66_117 V66 V117 -3.466264156206034e-19

R66_118 V66 V118 -2474.0768694962753
L66_118 V66 V118 -1.1647020388980518e-12
C66_118 V66 V118 -3.2672271431132177e-19

R66_119 V66 V119 -1850.854559934573
L66_119 V66 V119 -1.0285866169396692e-12
C66_119 V66 V119 -4.87392170848675e-19

R66_120 V66 V120 4103.429094253902
L66_120 V66 V120 -9.542262588709124e-12
C66_120 V66 V120 -1.7936509431314893e-19

R66_121 V66 V121 -2823.9339407730013
L66_121 V66 V121 1.4501662952992474e-12
C66_121 V66 V121 7.583522966828956e-20

R66_122 V66 V122 -1375.2185613040585
L66_122 V66 V122 8.970152480330268e-13
C66_122 V66 V122 3.027533089403751e-20

R66_123 V66 V123 13961.886132680344
L66_123 V66 V123 1.0894725564106778e-11
C66_123 V66 V123 -5.761818952259821e-20

R66_124 V66 V124 96871.891112324
L66_124 V66 V124 -3.395590597241777e-12
C66_124 V66 V124 -1.3526209980612632e-19

R66_125 V66 V125 1848.4340258777233
L66_125 V66 V125 -1.5023162991966268e-12
C66_125 V66 V125 -9.080302638844156e-20

R66_126 V66 V126 1510.7657071100778
L66_126 V66 V126 -1.226610223901927e-12
C66_126 V66 V126 1.0719374833952836e-19

R66_127 V66 V127 -9270.772151098827
L66_127 V66 V127 1.5576359413742681e-12
C66_127 V66 V127 -1.4741161908920373e-20

R66_128 V66 V128 6339.838989212094
L66_128 V66 V128 4.955774694839705e-11
C66_128 V66 V128 -6.308405846439549e-20

R66_129 V66 V129 7735.98619112976
L66_129 V66 V129 2.8375691963242243e-11
C66_129 V66 V129 -9.9593354416859e-20

R66_130 V66 V130 -321438.7842976258
L66_130 V66 V130 -1.5269438301021845e-12
C66_130 V66 V130 -2.6369435543768017e-19

R66_131 V66 V131 3855.3861748868717
L66_131 V66 V131 8.971936944028204e-12
C66_131 V66 V131 1.8354924023938828e-19

R66_132 V66 V132 87050.31455759928
L66_132 V66 V132 -3.0652320475144505e-12
C66_132 V66 V132 -6.625558705969115e-20

R66_133 V66 V133 17062.04212147391
L66_133 V66 V133 2.525696076885991e-12
C66_133 V66 V133 2.733115463778943e-19

R66_134 V66 V134 -3013.5347506022163
L66_134 V66 V134 -3.802927487978693e-12
C66_134 V66 V134 1.1693177732755831e-21

R66_135 V66 V135 -4267.85979974696
L66_135 V66 V135 2.5450004867195135e-12
C66_135 V66 V135 -5.504679037120611e-20

R66_136 V66 V136 9372.532971039178
L66_136 V66 V136 1.6149156140382933e-11
C66_136 V66 V136 4.795246198843781e-20

R66_137 V66 V137 1941.4372762076084
L66_137 V66 V137 -1.6794299016307993e-12
C66_137 V66 V137 -1.5644989214173582e-19

R66_138 V66 V138 1959.54773253968
L66_138 V66 V138 -1.008212616433462e-12
C66_138 V66 V138 -8.79673124922135e-20

R66_139 V66 V139 23173.83186737292
L66_139 V66 V139 9.576369351024554e-13
C66_139 V66 V139 1.2239204384175194e-19

R66_140 V66 V140 -2894.6504252818163
L66_140 V66 V140 -1.855107626380497e-12
C66_140 V66 V140 -5.565328045240509e-20

R66_141 V66 V141 3116.7095626889495
L66_141 V66 V141 -3.5964226970828128e-12
C66_141 V66 V141 -1.2495426429213313e-20

R66_142 V66 V142 -2191.2132092470206
L66_142 V66 V142 -2.0734089981419383e-12
C66_142 V66 V142 -1.0415964630629206e-19

R66_143 V66 V143 165113.12682771124
L66_143 V66 V143 -5.1844145983234446e-12
C66_143 V66 V143 5.352316358515911e-21

R66_144 V66 V144 -3821.160146142428
L66_144 V66 V144 3.282577313563414e-12
C66_144 V66 V144 -1.2204433149168617e-21

R67_67 V67 0 162.90240596345157
L67_67 V67 0 8.496235305362165e-14
C67_67 V67 0 1.6583953673959353e-18

R67_68 V67 V68 -4143.378280894969
L67_68 V67 V68 -2.386539818852452e-12
C67_68 V67 V68 -1.536900258093888e-20

R67_69 V67 V69 -7184.34254307945
L67_69 V67 V69 -1.173654850244657e-11
C67_69 V67 V69 2.6424292046695494e-20

R67_70 V67 V70 2314.227830512593
L67_70 V67 V70 1.731920976762458e-12
C67_70 V67 V70 2.301469644555036e-20

R67_71 V67 V71 840.0273056018921
L67_71 V67 V71 4.664429642837283e-13
C67_71 V67 V71 8.53627187663917e-20

R67_72 V67 V72 -5618.975084929181
L67_72 V67 V72 -2.335835896224625e-12
C67_72 V67 V72 -4.566859649335006e-20

R67_73 V67 V73 -2946.387682377671
L67_73 V67 V73 -1.4074137709745685e-12
C67_73 V67 V73 -4.3413039323506647e-20

R67_74 V67 V74 -16003.360386957856
L67_74 V67 V74 9.559557438870143e-12
C67_74 V67 V74 1.2803864633442678e-19

R67_75 V67 V75 -9133.610831637394
L67_75 V67 V75 -3.963874016507144e-12
C67_75 V67 V75 -5.092694368665367e-20

R67_76 V67 V76 -7326.337606647982
L67_76 V67 V76 1.2749586326111801e-11
C67_76 V67 V76 1.2340677427011465e-19

R67_77 V67 V77 -27672.764535367045
L67_77 V67 V77 1.3077589253832442e-11
C67_77 V67 V77 5.3322422742516656e-20

R67_78 V67 V78 -11523.552797080423
L67_78 V67 V78 -3.887281157746034e-12
C67_78 V67 V78 -4.861695577271652e-20

R67_79 V67 V79 -105529.09954408066
L67_79 V67 V79 3.491875557678992e-12
C67_79 V67 V79 1.733870109669447e-19

R67_80 V67 V80 9432.323133232092
L67_80 V67 V80 -1.2938903417876992e-11
C67_80 V67 V80 -1.4186997946228993e-19

R67_81 V67 V81 12177.639914466286
L67_81 V67 V81 9.88141111445479e-12
C67_81 V67 V81 2.5857472029489222e-20

R67_82 V67 V82 105674.25141861486
L67_82 V67 V82 -6.61911070672408e-11
C67_82 V67 V82 8.106400989631778e-20

R67_83 V67 V83 4352.004659162097
L67_83 V67 V83 1.8048535073948042e-12
C67_83 V67 V83 2.365792432343904e-20

R67_84 V67 V84 -9675.732344558897
L67_84 V67 V84 -7.228606247576214e-12
C67_84 V67 V84 4.096366869636108e-20

R67_85 V67 V85 31256.235091037433
L67_85 V67 V85 4.5453741284302775e-11
C67_85 V67 V85 4.4718427198126886e-20

R67_86 V67 V86 -6160.163549204472
L67_86 V67 V86 -2.51385591074372e-12
C67_86 V67 V86 -4.719153145778296e-20

R67_87 V67 V87 827319.4800519424
L67_87 V67 V87 8.321585826035e-12
C67_87 V67 V87 6.613610575753422e-20

R67_88 V67 V88 -165821.44807901225
L67_88 V67 V88 5.511986126497487e-11
C67_88 V67 V88 1.1520466396838648e-20

R67_89 V67 V89 -19410.021758031537
L67_89 V67 V89 1.249546570414286e-11
C67_89 V67 V89 3.1956747572023204e-20

R67_90 V67 V90 16547.92591371011
L67_90 V67 V90 -1.3275279992078948e-11
C67_90 V67 V90 -9.488488380310158e-20

R67_91 V67 V91 15623.87494809297
L67_91 V67 V91 4.32890971129867e-12
C67_91 V67 V91 9.828950315655208e-20

R67_92 V67 V92 -99180.8766012326
L67_92 V67 V92 1.2005279337566228e-10
C67_92 V67 V92 -3.691807309835464e-20

R67_93 V67 V93 4241.975101456614
L67_93 V67 V93 1.2585049031197713e-11
C67_93 V67 V93 2.6555464144036364e-20

R67_94 V67 V94 17223.508774907754
L67_94 V67 V94 -4.640922516050107e-12
C67_94 V67 V94 -1.1296272716796536e-19

R67_95 V67 V95 10397.38800291478
L67_95 V67 V95 8.423286378703704e-12
C67_95 V67 V95 4.751589934080727e-20

R67_96 V67 V96 -14957.18920263363
L67_96 V67 V96 -1.0290356376367826e-11
C67_96 V67 V96 -7.609344361059043e-20

R67_97 V67 V97 71215.45814999494
L67_97 V67 V97 -4.846597541030407e-12
C67_97 V67 V97 -7.831674082586712e-20

R67_98 V67 V98 7331.888422207927
L67_98 V67 V98 1.7413990019051834e-11
C67_98 V67 V98 -2.465220645415399e-20

R67_99 V67 V99 13464.919325047349
L67_99 V67 V99 6.734949400405747e-12
C67_99 V67 V99 1.6987202456131303e-20

R67_100 V67 V100 -31791.028598321507
L67_100 V67 V100 -4.4509877912096586e-11
C67_100 V67 V100 1.0110750144556824e-20

R67_101 V67 V101 22261.178863490197
L67_101 V67 V101 8.9790871695725e-12
C67_101 V67 V101 -3.405780061300013e-21

R67_102 V67 V102 16177.225540882615
L67_102 V67 V102 -2.49932732716861e-12
C67_102 V67 V102 -2.2351589959366024e-19

R67_103 V67 V103 36656.08188981609
L67_103 V67 V103 2.7671333390297365e-12
C67_103 V67 V103 2.0334570895893482e-19

R67_104 V67 V104 -38830.08289886132
L67_104 V67 V104 -2.1148069930414475e-11
C67_104 V67 V104 -4.137006501523601e-20

R67_105 V67 V105 -54704.124349664715
L67_105 V67 V105 1.3950804378186126e-11
C67_105 V67 V105 3.601185738176445e-20

R67_106 V67 V106 -8820.469278325618
L67_106 V67 V106 -6.836494403266621e-12
C67_106 V67 V106 -7.141954772384868e-20

R67_107 V67 V107 -12120.828045123475
L67_107 V67 V107 -2.1437284941899e-12
C67_107 V67 V107 -2.2839198387062626e-19

R67_108 V67 V108 5657.551703182001
L67_108 V67 V108 2.7618228827169506e-12
C67_108 V67 V108 2.003338966843957e-19

R67_109 V67 V109 24756.7012590499
L67_109 V67 V109 5.9034738375601155e-12
C67_109 V67 V109 4.1182908628528066e-20

R67_110 V67 V110 8727.584737163314
L67_110 V67 V110 -5.1742280361956314e-12
C67_110 V67 V110 -4.392488895597171e-20

R67_111 V67 V111 -9179.205089252517
L67_111 V67 V111 3.1113376611678905e-12
C67_111 V67 V111 1.0365894472817454e-19

R67_112 V67 V112 162180.57425141317
L67_112 V67 V112 -3.648924202792289e-12
C67_112 V67 V112 -1.6375036641243164e-19

R67_113 V67 V113 -135565.56622005254
L67_113 V67 V113 -1.2728471391486921e-11
C67_113 V67 V113 -1.5864391215632466e-20

R67_114 V67 V114 23828.10741635005
L67_114 V67 V114 -1.4172389853533652e-11
C67_114 V67 V114 -1.5372987425611338e-20

R67_115 V67 V115 7145.905877850943
L67_115 V67 V115 -3.671183851903214e-12
C67_115 V67 V115 -1.1870222620697208e-19

R67_116 V67 V116 23112.73785375112
L67_116 V67 V116 6.7053560861324865e-12
C67_116 V67 V116 7.407542191487506e-20

R67_117 V67 V117 8387.762901878505
L67_117 V67 V117 1.2249505166712415e-10
C67_117 V67 V117 2.784735742836291e-20

R67_118 V67 V118 -22775.290084387405
L67_118 V67 V118 2.0145837561199435e-10
C67_118 V67 V118 -1.3436158743481861e-20

R67_119 V67 V119 -6709.560457430475
L67_119 V67 V119 8.257636169966443e-12
C67_119 V67 V119 2.804457093462981e-20

R67_120 V67 V120 3197.0050318861263
L67_120 V67 V120 -3.171978845400243e-12
C67_120 V67 V120 4.7934067858252556e-20

R67_121 V67 V121 -12044.223830225505
L67_121 V67 V121 1.2788290270512474e-11
C67_121 V67 V121 8.69222320478669e-21

R67_122 V67 V122 4839.723446170063
L67_122 V67 V122 -3.506852786401784e-12
C67_122 V67 V122 1.4984903042750685e-20

R67_123 V67 V123 14352.629512650305
L67_123 V67 V123 -7.766772531661896e-12
C67_123 V67 V123 -2.767625450285377e-20

R67_124 V67 V124 53937.941462830044
L67_124 V67 V124 1.5521303266773717e-11
C67_124 V67 V124 2.0119918918358285e-20

R67_125 V67 V125 3739.1520723113363
L67_125 V67 V125 -5.1412309890097424e-12
C67_125 V67 V125 2.3715951157939458e-21

R67_126 V67 V126 -3332.923328129302
L67_126 V67 V126 2.205417534994086e-12
C67_126 V67 V126 -3.528123437453092e-20

R67_127 V67 V127 3273.498991605343
L67_127 V67 V127 -2.479360433331267e-12
C67_127 V67 V127 7.689883917419604e-21

R67_128 V67 V128 22748.076897016603
L67_128 V67 V128 -1.8965393308482744e-11
C67_128 V67 V128 -3.3592855280938884e-20

R67_129 V67 V129 5570.497593107772
L67_129 V67 V129 -6.018479590719279e-12
C67_129 V67 V129 -1.383587231783744e-20

R67_130 V67 V130 -39635.46359701381
L67_130 V67 V130 3.327698803323893e-12
C67_130 V67 V130 6.095370105375981e-20

R67_131 V67 V131 -10849.024257512096
L67_131 V67 V131 -9.576633187866753e-11
C67_131 V67 V131 -6.3760026028647e-20

R67_132 V67 V132 -13023.39638381452
L67_132 V67 V132 1.4399809569525425e-11
C67_132 V67 V132 -1.3651390565730917e-20

R67_133 V67 V133 -19969.770095241278
L67_133 V67 V133 -1.196024624400344e-11
C67_133 V67 V133 -3.7384554578005984e-20

R67_134 V67 V134 -7098.911978182967
L67_134 V67 V134 7.916092931574967e-11
C67_134 V67 V134 -3.60437747743364e-21

R67_135 V67 V135 7335.264845541198
L67_135 V67 V135 -3.783559445102979e-12
C67_135 V67 V135 2.6583443093481613e-20

R67_136 V67 V136 60709.60217888301
L67_136 V67 V136 3.41062890574433e-11
C67_136 V67 V136 3.194670851989016e-20

R67_137 V67 V137 5569.844255039804
L67_137 V67 V137 3.6318360972083566e-11
C67_137 V67 V137 5.132913135393579e-20

R67_138 V67 V138 -3070.6753856561563
L67_138 V67 V138 2.137800797093846e-12
C67_138 V67 V138 2.1816782102499598e-20

R67_139 V67 V139 2045.58847934054
L67_139 V67 V139 -1.6847522007538575e-12
C67_139 V67 V139 -4.517524619465873e-20

R67_140 V67 V140 -11224.576012596986
L67_140 V67 V140 4.670792089601579e-12
C67_140 V67 V140 4.371953640000059e-20

R67_141 V67 V141 269106.5401299418
L67_141 V67 V141 8.927969193808371e-12
C67_141 V67 V141 1.1387837134527862e-20

R67_142 V67 V142 -6018.510696844464
L67_142 V67 V142 6.897039972261666e-12
C67_142 V67 V142 -3.335047393418623e-21

R67_143 V67 V143 -8075.699632068353
L67_143 V67 V143 7.054013656891689e-12
C67_143 V67 V143 -3.5317794916431255e-20

R67_144 V67 V144 -7615.222811596671
L67_144 V67 V144 -8.020379788302225e-12
C67_144 V67 V144 -8.377510492266581e-21

R68_68 V68 0 135.47397630335686
L68_68 V68 0 1.1316302230849204e-13
C68_68 V68 0 9.450296569538209e-19

R68_69 V68 V69 7266.051990312037
L68_69 V68 V69 4.756716785834782e-12
C68_69 V68 V69 -2.538718701441633e-20

R68_70 V68 V70 9025.773467589504
L68_70 V68 V70 7.439911257416892e-12
C68_70 V68 V70 1.1447753355062749e-20

R68_71 V68 V71 4662.457946035465
L68_71 V68 V71 2.6023820928011155e-12
C68_71 V68 V71 1.3702668945121155e-20

R68_72 V68 V72 5034.971435503033
L68_72 V68 V72 -1.859312465160046e-11
C68_72 V68 V72 2.796647589730953e-20

R68_73 V68 V73 -3653.326132177311
L68_73 V68 V73 -5.435286182777803e-12
C68_73 V68 V73 -4.893573347164501e-20

R68_74 V68 V74 -42181.178542973284
L68_74 V68 V74 8.660539598135388e-12
C68_74 V68 V74 -2.4934134943019657e-20

R68_75 V68 V75 -21397.424810874076
L68_75 V68 V75 -1.15638479709183e-11
C68_75 V68 V75 -3.8205890233918336e-20

R68_76 V68 V76 -8232.359600105292
L68_76 V68 V76 -7.468098549070744e-12
C68_76 V68 V76 -1.387417964142149e-20

R68_77 V68 V77 14391.748314735827
L68_77 V68 V77 5.91480490229807e-12
C68_77 V68 V77 5.385254302824937e-20

R68_78 V68 V78 207438.34276290674
L68_78 V68 V78 9.98591629922831e-12
C68_78 V68 V78 4.854477701538712e-20

R68_79 V68 V79 -34881.753349050436
L68_79 V68 V79 1.6285918881899516e-09
C68_79 V68 V79 -2.5424081088678542e-20

R68_80 V68 V80 9048.988985274787
L68_80 V68 V80 2.16364726665502e-11
C68_80 V68 V80 1.0516951019849143e-19

R68_81 V68 V81 -10416.012551237203
L68_81 V68 V81 -6.7675135301900645e-12
C68_81 V68 V81 -2.1727940657518916e-19

R68_82 V68 V82 -12624.136126831783
L68_82 V68 V82 -2.4630572657807217e-12
C68_82 V68 V82 -1.7116885582453576e-19

R68_83 V68 V83 19738.769320959564
L68_83 V68 V83 -8.193262414573283e-12
C68_83 V68 V83 -2.6772456945068487e-20

R68_84 V68 V84 65655.62924149034
L68_84 V68 V84 -7.535646569346232e-12
C68_84 V68 V84 -3.752882671260059e-20

R68_85 V68 V85 293190.7020942575
L68_85 V68 V85 1.3777707079059051e-11
C68_85 V68 V85 8.483557561955925e-21

R68_86 V68 V86 -16287.77234791362
L68_86 V68 V86 5.012565756800973e-12
C68_86 V68 V86 1.2926999009580973e-19

R68_87 V68 V87 -1400610.5847564614
L68_87 V68 V87 5.077481479739367e-12
C68_87 V68 V87 3.312316113665778e-20

R68_88 V68 V88 267870.92486198596
L68_88 V68 V88 6.393660569717457e-11
C68_88 V68 V88 -3.973329897077407e-20

R68_89 V68 V89 -87614.21418001207
L68_89 V68 V89 -1.2853308854514004e-11
C68_89 V68 V89 -1.1928056753173986e-20

R68_90 V68 V90 66132.13044270818
L68_90 V68 V90 6.370896632441846e-11
C68_90 V68 V90 2.810492116529752e-20

R68_91 V68 V91 -15773.898058301016
L68_91 V68 V91 -2.2235353587475297e-12
C68_91 V68 V91 -2.6389716673544005e-19

R68_92 V68 V92 29533.00908571655
L68_92 V68 V92 -1.164976119130722e-10
C68_92 V68 V92 1.520803997152734e-19

R68_93 V68 V93 17050.422259524308
L68_93 V68 V93 1.7921813389421033e-11
C68_93 V68 V93 6.922790542442451e-22

R68_94 V68 V94 35021.337664878985
L68_94 V68 V94 1.3301151701793826e-11
C68_94 V68 V94 -2.638227303791211e-20

R68_95 V68 V95 -81649.54301951456
L68_95 V68 V95 -5.2004440697970395e-12
C68_95 V68 V95 -9.88066319701104e-20

R68_96 V68 V96 9997.294722561734
L68_96 V68 V96 7.375490342843494e-12
C68_96 V68 V96 2.434230908871159e-19

R68_97 V68 V97 68074.74580641955
L68_97 V68 V97 6.008485807408298e-11
C68_97 V68 V97 -2.036514525921084e-20

R68_98 V68 V98 21233.35669689184
L68_98 V68 V98 -6.978966848200264e-12
C68_98 V68 V98 -2.548747979169397e-21

R68_99 V68 V99 65701.44454583073
L68_99 V68 V99 2.6032621551574198e-11
C68_99 V68 V99 -1.3983456175457857e-20

R68_100 V68 V100 85101.19030508093
L68_100 V68 V100 -1.9291451150968694e-10
C68_100 V68 V100 -1.0033863367269587e-19

R68_101 V68 V101 42486.78550846458
L68_101 V68 V101 -7.957920524444623e-12
C68_101 V68 V101 4.972128335884116e-21

R68_102 V68 V102 73942.9108248106
L68_102 V68 V102 -5.482050481911174e-12
C68_102 V68 V102 -1.321395186812166e-20

R68_103 V68 V103 -26906.147551569225
L68_103 V68 V103 -1.188067187339942e-10
C68_103 V68 V103 -5.084278452385038e-20

R68_104 V68 V104 20765.90196169822
L68_104 V68 V104 6.873074455643891e-12
C68_104 V68 V104 1.9289946067329868e-19

R68_105 V68 V105 36788.07731012315
L68_105 V68 V105 4.060716369775327e-12
C68_105 V68 V105 2.9484566500003425e-20

R68_106 V68 V106 -16986.951938284394
L68_106 V68 V106 -2.4661350181168425e-12
C68_106 V68 V106 -1.3667414709355629e-19

R68_107 V68 V107 88348.06413419511
L68_107 V68 V107 -6.0473452660120786e-12
C68_107 V68 V107 -1.901856653986706e-20

R68_108 V68 V108 25943.08715504829
L68_108 V68 V108 7.277292608048536e-12
C68_108 V68 V108 -7.993292293412806e-20

R68_109 V68 V109 -199454.2554304519
L68_109 V68 V109 7.936477434691379e-12
C68_109 V68 V109 1.6901882399317784e-19

R68_110 V68 V110 35837.272369975886
L68_110 V68 V110 3.2749827780464204e-12
C68_110 V68 V110 1.0683393038767371e-19

R68_111 V68 V111 -36955.10664384141
L68_111 V68 V111 7.715789273004083e-12
C68_111 V68 V111 -4.770221109663266e-21

R68_112 V68 V112 -208784.6373355306
L68_112 V68 V112 -5.42985557061774e-12
C68_112 V68 V112 2.235481241470627e-20

R68_113 V68 V113 39663.20879016232
L68_113 V68 V113 -6.140619492515399e-12
C68_113 V68 V113 -1.2206670225853578e-19

R68_114 V68 V114 -54465.474101426604
L68_114 V68 V114 -6.144068258802517e-12
C68_114 V68 V114 -2.587173705410826e-20

R68_115 V68 V115 42544.26845787154
L68_115 V68 V115 -1.7882251877512082e-11
C68_115 V68 V115 2.662423220579506e-20

R68_116 V68 V116 93592.24216076931
L68_116 V68 V116 1.2660167571915397e-11
C68_116 V68 V116 -6.605931122723635e-20

R68_117 V68 V117 54721.792322629175
L68_117 V68 V117 7.667175462680293e-12
C68_117 V68 V117 8.84128205669579e-20

R68_118 V68 V118 -613417.9873955938
L68_118 V68 V118 4.176045398664045e-12
C68_118 V68 V118 1.401225737383852e-19

R68_119 V68 V119 -135704.6151712498
L68_119 V68 V119 6.028344282570265e-12
C68_119 V68 V119 -1.6036680490727753e-20

R68_120 V68 V120 19355.6751801292
L68_120 V68 V120 -1.8288481672094944e-11
C68_120 V68 V120 -6.657056637964707e-20

R68_121 V68 V121 -21049.311791336942
L68_121 V68 V121 -1.09939424152601e-11
C68_121 V68 V121 -2.1306157910701752e-20

R68_122 V68 V122 82014.11370445247
L68_122 V68 V122 -1.1164989262846874e-11
C68_122 V68 V122 9.331089603895486e-21

R68_123 V68 V123 -96177.84209609406
L68_123 V68 V123 2.1653426752268472e-10
C68_123 V68 V123 1.4387610111754726e-20

R68_124 V68 V124 -313839.8227101687
L68_124 V68 V124 2.905690396584203e-11
C68_124 V68 V124 -4.5978935869234264e-20

R68_125 V68 V125 25782.71306197745
L68_125 V68 V125 1.2715271342403855e-11
C68_125 V68 V125 2.7640778486310044e-20

R68_126 V68 V126 -86315.5038299171
L68_126 V68 V126 8.856209313041898e-12
C68_126 V68 V126 3.145604016736847e-22

R68_127 V68 V127 19241.51743724231
L68_127 V68 V127 -9.64314125664474e-12
C68_127 V68 V127 -2.554545580535339e-20

R68_128 V68 V128 191408.58648586468
L68_128 V68 V128 2.65633921886114e-11
C68_128 V68 V128 5.51234171253351e-20

R68_129 V68 V129 470003.5057012731
L68_129 V68 V129 -2.6457636027998006e-11
C68_129 V68 V129 -1.920314081256522e-20

R68_130 V68 V130 64048.652232982124
L68_130 V68 V130 8.471112470875843e-12
C68_130 V68 V130 6.175699525291152e-20

R68_131 V68 V131 67513.076737524
L68_131 V68 V131 3.449298077956431e-10
C68_131 V68 V131 3.1726716169605005e-20

R68_132 V68 V132 -30081.85619634411
L68_132 V68 V132 4.3377847004848404e-10
C68_132 V68 V132 -3.4309275046124735e-20

R68_133 V68 V133 -89818.42429894717
L68_133 V68 V133 -5.880117665325733e-12
C68_133 V68 V133 -9.179092466907164e-20

R68_134 V68 V134 -19431.929101950227
L68_134 V68 V134 2.8006512390303842e-11
C68_134 V68 V134 1.832382177414931e-20

R68_135 V68 V135 54603.69151154066
L68_135 V68 V135 -2.8053424002720676e-11
C68_135 V68 V135 3.3856859274423726e-21

R68_136 V68 V136 53850.173138979306
L68_136 V68 V136 -3.591298819544248e-11
C68_136 V68 V136 -2.2627926701192998e-20

R68_137 V68 V137 21857.469648556285
L68_137 V68 V137 1.017633371406988e-11
C68_137 V68 V137 2.093119654495982e-20

R68_138 V68 V138 -518390.0504799774
L68_138 V68 V138 1.9642251518105223e-11
C68_138 V68 V138 -6.672946385056144e-20

R68_139 V68 V139 11148.47749887841
L68_139 V68 V139 -6.290749601855947e-12
C68_139 V68 V139 -2.923816438641912e-20

R68_140 V68 V140 -48299.081040694145
L68_140 V68 V140 1.8400261380378172e-11
C68_140 V68 V140 -5.826223573776203e-21

R68_141 V68 V141 -225586.3021091102
L68_141 V68 V141 4.556647035174726e-11
C68_141 V68 V141 -1.1279950625294624e-20

R68_142 V68 V142 26290.36987961111
L68_142 V68 V142 1.1523050758687963e-11
C68_142 V68 V142 -3.110563749557351e-21

R68_143 V68 V143 261707.35451474402
L68_143 V68 V143 7.528187315979302e-11
C68_143 V68 V143 -2.112053537433897e-20

R68_144 V68 V144 780750.1747642037
L68_144 V68 V144 2.5022885883867315e-11
C68_144 V68 V144 4.510394071104482e-20

R69_69 V69 0 -132.16161384195487
L69_69 V69 0 -1.2675572063810448e-13
C69_69 V69 0 -3.1600763942436535e-19

R69_70 V69 V70 5798.404806121902
L69_70 V69 V70 -7.313149189399385e-12
C69_70 V69 V70 4.741459724220932e-20

R69_71 V69 V71 2204.5525129783946
L69_71 V69 V71 2.664540821619124e-12
C69_71 V69 V71 -1.0284997624515844e-19

R69_72 V69 V72 -2595.240547651989
L69_72 V69 V72 -1.2903748046457571e-12
C69_72 V69 V72 8.024910675508362e-20

R69_73 V69 V73 -4228.526040773437
L69_73 V69 V73 -2.194151968159615e-12
C69_73 V69 V73 -1.5653092118454914e-20

R69_74 V69 V74 -2090.0512789102077
L69_74 V69 V74 -3.449800110564249e-12
C69_74 V69 V74 -1.2159862086089862e-20

R69_75 V69 V75 8363.97798977232
L69_75 V69 V75 1.7290526617456124e-12
C69_75 V69 V75 1.1153467512048698e-19

R69_76 V69 V76 29760.710681655517
L69_76 V69 V76 2.688889683762151e-12
C69_76 V69 V76 -2.265550521672878e-20

R69_77 V69 V77 -68885.48062707804
L69_77 V69 V77 4.463674847033361e-12
C69_77 V69 V77 4.322576041876262e-20

R69_78 V69 V78 34433.52274192852
L69_78 V69 V78 3.3431979473414247e-12
C69_78 V69 V78 -3.9547475285514924e-20

R69_79 V69 V79 -4854.175026197657
L69_79 V69 V79 -3.9588943374682775e-12
C69_79 V69 V79 -8.168833598088707e-20

R69_80 V69 V80 9879.65762564745
L69_80 V69 V80 5.413934181260793e-12
C69_80 V69 V80 1.5641901043755332e-19

R69_81 V69 V81 976791.8073072876
L69_81 V69 V81 -2.6041484054656955e-12
C69_81 V69 V81 -1.1107020728592806e-19

R69_82 V69 V82 -11609.627205617542
L69_82 V69 V82 -3.349795230919063e-12
C69_82 V69 V82 -2.0223240374460689e-19

R69_83 V69 V83 15412.142050847662
L69_83 V69 V83 -1.548242057317195e-10
C69_83 V69 V83 -7.056332703640274e-20

R69_84 V69 V84 -6642.448912000469
L69_84 V69 V84 -2.1129975229659085e-12
C69_84 V69 V84 -7.60601541005875e-20

R69_85 V69 V85 -8357.023276907492
L69_85 V69 V85 -2.4508801029809863e-12
C69_85 V69 V85 -9.154621609251293e-20

R69_86 V69 V86 -9592.679205363174
L69_86 V69 V86 1.401031584301918e-11
C69_86 V69 V86 1.2780438765809272e-19

R69_87 V69 V87 -23966.280096018047
L69_87 V69 V87 3.374845357775922e-12
C69_87 V69 V87 1.5489339114123831e-19

R69_88 V69 V88 63176.71203150346
L69_88 V69 V88 7.464619193987945e-12
C69_88 V69 V88 5.467219080766801e-20

R69_89 V69 V89 16425.623304933677
L69_89 V69 V89 3.803188029362425e-12
C69_89 V69 V89 5.576524794257133e-20

R69_90 V69 V90 8077.684730828411
L69_90 V69 V90 2.5016603815173135e-12
C69_90 V69 V90 1.9500307384167832e-19

R69_91 V69 V91 -15717.501724081114
L69_91 V69 V91 -2.1521418627891635e-12
C69_91 V69 V91 -2.9851105210203763e-19

R69_92 V69 V92 84102.24861512736
L69_92 V69 V92 7.504686957813922e-12
C69_92 V69 V92 3.048988549936184e-20

R69_93 V69 V93 -31508.92552652832
L69_93 V69 V93 1.12721676122617e-10
C69_93 V69 V93 4.3378696652761765e-20

R69_94 V69 V94 41788.38269270724
L69_94 V69 V94 -1.1851209519869205e-11
C69_94 V69 V94 4.287473101261702e-20

R69_95 V69 V95 -112768.9107859543
L69_95 V69 V95 -6.29586679527645e-12
C69_95 V69 V95 -1.09412791338298e-19

R69_96 V69 V96 13475.965239767853
L69_96 V69 V96 3.5984122598239955e-12
C69_96 V69 V96 8.998049364495416e-20

R69_97 V69 V97 88877.121203456
L69_97 V69 V97 4.083027736237561e-12
C69_97 V69 V97 1.2168450501485286e-19

R69_98 V69 V98 -16492.9567539878
L69_98 V69 V98 6.701809993351668e-12
C69_98 V69 V98 -1.3530568729143874e-20

R69_99 V69 V99 -32352.306419600533
L69_99 V69 V99 -1.4255622526474117e-11
C69_99 V69 V99 -7.322500202482569e-21

R69_100 V69 V100 46264.38534978183
L69_100 V69 V100 1.1276588801878537e-10
C69_100 V69 V100 1.1865405326243698e-20

R69_101 V69 V101 -194042.12648097787
L69_101 V69 V101 9.526734359435183e-12
C69_101 V69 V101 -7.633109709137978e-21

R69_102 V69 V102 10700.489485079794
L69_102 V69 V102 1.911086487058455e-12
C69_102 V69 V102 3.16078287654917e-19

R69_103 V69 V103 -7673.702857318334
L69_103 V69 V103 -3.868426973644365e-12
C69_103 V69 V103 -1.8206849221810282e-19

R69_104 V69 V104 12688.80374241658
L69_104 V69 V104 2.5720995129129877e-12
C69_104 V69 V104 2.3617645600291476e-19

R69_105 V69 V105 21361.1019444098
L69_105 V69 V105 -1.5546050042575288e-11
C69_105 V69 V105 -2.952219993804498e-20

R69_106 V69 V106 13166.004045286023
L69_106 V69 V106 -7.111598449204514e-12
C69_106 V69 V106 -9.466495917815681e-20

R69_107 V69 V107 17022.294782033438
L69_107 V69 V107 4.8114567399095265e-12
C69_107 V69 V107 1.4033278819912176e-19

R69_108 V69 V108 -10940.739396961531
L69_108 V69 V108 -3.905744846462889e-12
C69_108 V69 V108 -1.8137803759873445e-19

R69_109 V69 V109 -86266.28588312372
L69_109 V69 V109 1.0104267570130625e-11
C69_109 V69 V109 2.1101253870754676e-20

R69_110 V69 V110 38803.2109604049
L69_110 V69 V110 1.548794439092753e-11
C69_110 V69 V110 6.619574103125982e-20

R69_111 V69 V111 -24166.626269271463
L69_111 V69 V111 8.000259826709433e-11
C69_111 V69 V111 -1.8272803786403847e-20

R69_112 V69 V112 21444.916601373166
L69_112 V69 V112 3.769620301727703e-12
C69_112 V69 V112 4.8642351479173755e-20

R69_113 V69 V113 125193.95797653538
L69_113 V69 V113 8.618837925351652e-12
C69_113 V69 V113 3.7406742921579516e-20

R69_114 V69 V114 46383.50189865114
L69_114 V69 V114 -1.3057063161284554e-11
C69_114 V69 V114 -1.0268630245819704e-19

R69_115 V69 V115 20786.20874605168
L69_115 V69 V115 8.82153267266381e-12
C69_115 V69 V115 8.977574691674588e-20

R69_116 V69 V116 -26223.904121775893
L69_116 V69 V116 -4.454154881368733e-12
C69_116 V69 V116 -1.2158329762349821e-19

R69_117 V69 V117 -22269.213214487707
L69_117 V69 V117 -8.018846016990218e-12
C69_117 V69 V117 -1.0762084279964788e-19

R69_118 V69 V118 17070.756318305823
L69_118 V69 V118 1.2551309037684913e-11
C69_118 V69 V118 8.991395327802573e-20

R69_119 V69 V119 -127463.43028680267
L69_119 V69 V119 8.564269519744848e-12
C69_119 V69 V119 1.0397215910832343e-19

R69_120 V69 V120 -46803.3563700734
L69_120 V69 V120 -2.35420298732746e-11
C69_120 V69 V120 -9.84297590514178e-21

R69_121 V69 V121 -18786.744738447
L69_121 V69 V121 7.666631590880156e-12
C69_121 V69 V121 -9.787302730651446e-21

R69_122 V69 V122 56016.70354604121
L69_122 V69 V122 2.754767639775908e-12
C69_122 V69 V122 1.1487720624947415e-20

R69_123 V69 V123 143471.96890057655
L69_123 V69 V123 1.8398508375641826e-11
C69_123 V69 V123 -9.686351901693112e-21

R69_124 V69 V124 -88752.05013083038
L69_124 V69 V124 -6.993897284499379e-11
C69_124 V69 V124 -2.0220873287938387e-20

R69_125 V69 V125 23409.14489755382
L69_125 V69 V125 -6.447570889476673e-12
C69_125 V69 V125 1.3628688521592395e-20

R69_126 V69 V126 -39751.72587901999
L69_126 V69 V126 -4.6958994374782484e-12
C69_126 V69 V126 4.0312446215315537e-20

R69_127 V69 V127 -146445.94146923153
L69_127 V69 V127 7.492913641932128e-12
C69_127 V69 V127 -7.7267577256817e-21

R69_128 V69 V128 -21374.73963527699
L69_128 V69 V128 -1.0137725999388688e-11
C69_128 V69 V128 -5.810758411553552e-20

R69_129 V69 V129 -74119.94714149335
L69_129 V69 V129 -2.6424633120375462e-11
C69_129 V69 V129 -7.404261589013761e-20

R69_130 V69 V130 -12153.362289581253
L69_130 V69 V130 -4.605063876324373e-12
C69_130 V69 V130 -8.069548733599512e-20

R69_131 V69 V131 -59307.34613150856
L69_131 V69 V131 -3.143950268540998e-11
C69_131 V69 V131 7.289824775317474e-20

R69_132 V69 V132 -73203.31162027057
L69_132 V69 V132 -3.970127190374912e-12
C69_132 V69 V132 -1.173565908267205e-19

R69_133 V69 V133 75610.29274061165
L69_133 V69 V133 -7.488275625509243e-12
C69_133 V69 V133 -6.990848952529895e-20

R69_134 V69 V134 22649.502820595266
L69_134 V69 V134 -6.147089680539864e-11
C69_134 V69 V134 4.633730633735874e-20

R69_135 V69 V135 166853.1539203174
L69_135 V69 V135 8.971558031352572e-12
C69_135 V69 V135 -1.0173451119913704e-20

R69_136 V69 V136 -52547.30307345716
L69_136 V69 V136 1.0535286329333949e-11
C69_136 V69 V136 1.0168861753775204e-19

R69_137 V69 V137 -37915.60180074188
L69_137 V69 V137 -1.2651952288070151e-11
C69_137 V69 V137 4.3951761489242114e-20

R69_138 V69 V138 -13511.44501871808
L69_138 V69 V138 -2.700530850828126e-12
C69_138 V69 V138 -6.891179602523943e-20

R69_139 V69 V139 49767.31180338056
L69_139 V69 V139 4.925167054549154e-12
C69_139 V69 V139 -6.633642158627374e-21

R69_140 V69 V140 24979.084125860383
L69_140 V69 V140 -1.3030648070285073e-11
C69_140 V69 V140 1.7635003620437902e-20

R69_141 V69 V141 -112026.82186094175
L69_141 V69 V141 -3.218271528966004e-10
C69_141 V69 V141 2.721551289088473e-20

R69_142 V69 V142 44654.52601294482
L69_142 V69 V142 -6.605462870184371e-12
C69_142 V69 V142 -5.751046945920253e-20

R69_143 V69 V143 -42767.637392231074
L69_143 V69 V143 -1.3098500565905424e-11
C69_143 V69 V143 -2.2256596851152284e-20

R69_144 V69 V144 290851.8475144214
L69_144 V69 V144 1.2667934253126447e-11
C69_144 V69 V144 -2.6851841285934505e-20

R70_70 V70 0 -136.50603543397628
L70_70 V70 0 -1.0089335830663487e-12
C70_70 V70 0 6.503489572595892e-19

R70_71 V70 V71 -1746.9285508029488
L70_71 V70 V71 -7.057911773699576e-13
C70_71 V70 V71 -1.9706503826210422e-19

R70_72 V70 V72 -3431.9323675659043
L70_72 V70 V72 -1.571058376729111e-12
C70_72 V70 V72 -9.867562577646852e-20

R70_73 V70 V73 10124.726644218314
L70_73 V70 V73 -5.345009674871845e-12
C70_73 V70 V73 -6.542803560897876e-20

R70_74 V70 V74 32756.762256520735
L70_74 V70 V74 -3.908130320680077e-12
C70_74 V70 V74 2.5619942046683762e-20

R70_75 V70 V75 3265.5865384933527
L70_75 V70 V75 1.4349724267154596e-12
C70_75 V70 V75 2.937493654375911e-19

R70_76 V70 V76 7568.455482006235
L70_76 V70 V76 -6.724907219702383e-12
C70_76 V70 V76 -3.6111095542254965e-19

R70_77 V70 V77 9352.256636967519
L70_77 V70 V77 3.989731450308445e-12
C70_77 V70 V77 1.8281043421541436e-20

R70_78 V70 V78 -9461.933609215113
L70_78 V70 V78 -2.4021002669313477e-12
C70_78 V70 V78 -3.2357896059181003e-19

R70_79 V70 V79 -9886.41671208698
L70_79 V70 V79 -1.5394209881153954e-12
C70_79 V70 V79 -3.689257050156508e-19

R70_80 V70 V80 10640.529823461091
L70_80 V70 V80 2.127983315055848e-12
C70_80 V70 V80 4.4296290125738015e-19

R70_81 V70 V81 -8696.432217122006
L70_81 V70 V81 -1.4590327706411252e-12
C70_81 V70 V81 -2.1347856072494888e-19

R70_82 V70 V82 3191.818789416221
L70_82 V70 V82 6.189247961113721e-13
C70_82 V70 V82 8.193221428456185e-19

R70_83 V70 V83 8955.030733505302
L70_83 V70 V83 1.1421140672631556e-12
C70_83 V70 V83 7.305955985212609e-19

R70_84 V70 V84 39760.67054077793
L70_84 V70 V84 -3.3040920457585247e-12
C70_84 V70 V84 -1.0895615494278207e-19

R70_85 V70 V85 -4786.451090254258
L70_85 V70 V85 -1.1057922342981464e-12
C70_85 V70 V85 -4.333732446398919e-19

R70_86 V70 V86 -25088.824709119657
L70_86 V70 V86 -1.9292266205793258e-12
C70_86 V70 V86 -3.044079391732945e-19

R70_87 V70 V87 -5756.042674259881
L70_87 V70 V87 -1.021298624856146e-12
C70_87 V70 V87 -6.121676205611401e-19

R70_88 V70 V88 -21703.710052774994
L70_88 V70 V88 -4.248060894402567e-12
C70_88 V70 V88 -1.77683244206488e-19

R70_89 V70 V89 5276.781368494158
L70_89 V70 V89 1.6205014295243777e-12
C70_89 V70 V89 2.929463462819054e-19

R70_90 V70 V90 20030.382965391644
L70_90 V70 V90 2.3020548341438627e-12
C70_90 V70 V90 3.0332466722910425e-19

R70_91 V70 V91 5045.077642586724
L70_91 V70 V91 8.487986353137035e-13
C70_91 V70 V91 7.30541088430657e-19

R70_92 V70 V92 5045.149333177141
L70_92 V70 V92 1.0677512786037023e-12
C70_92 V70 V92 5.428421793189224e-19

R70_93 V70 V93 -6515.948046164074
L70_93 V70 V93 -3.5569475259607225e-12
C70_93 V70 V93 -1.2264200628615564e-19

R70_94 V70 V94 -10095.1200494942
L70_94 V70 V94 -2.054460722066632e-12
C70_94 V70 V94 -2.037237609099059e-19

R70_95 V70 V95 6753.777927965271
L70_95 V70 V95 1.5185045948162868e-12
C70_95 V70 V95 4.3174236961083086e-19

R70_96 V70 V96 5719.310239731234
L70_96 V70 V96 1.5506261465191687e-12
C70_96 V70 V96 3.9378863313579065e-19

R70_97 V70 V97 -5858.792480276625
L70_97 V70 V97 -5.133756389934377e-12
C70_97 V70 V97 -1.0207071025824069e-19

R70_98 V70 V98 -11640.538687729328
L70_98 V70 V98 1.19014634872412e-12
C70_98 V70 V98 4.792268596701843e-19

R70_99 V70 V99 -16856.4125094694
L70_99 V70 V99 -3.4048528001492087e-12
C70_99 V70 V99 -1.0233766772624246e-19

R70_100 V70 V100 4268220.870352597
L70_100 V70 V100 -4.143502616265871e-12
C70_100 V70 V100 -1.173171812897734e-19

R70_101 V70 V101 11321.298111476493
L70_101 V70 V101 1.21827248705813e-12
C70_101 V70 V101 4.933364783941216e-19

R70_102 V70 V102 3872.3450924645435
L70_102 V70 V102 7.041305093417172e-13
C70_102 V70 V102 9.065505283445376e-19

R70_103 V70 V103 -4823.919345161936
L70_103 V70 V103 -1.8867643169881887e-12
C70_103 V70 V103 -4.484282032678171e-19

R70_104 V70 V104 10803.532005483125
L70_104 V70 V104 9.66394519495569e-12
C70_104 V70 V104 8.583917092044248e-20

R70_105 V70 V105 -9219.41173437997
L70_105 V70 V105 -8.78060016604642e-13
C70_105 V70 V105 -6.771882739601089e-19

R70_106 V70 V106 1687.0385149199071
L70_106 V70 V106 5.441258680372294e-13
C70_106 V70 V106 1.2143569619042212e-18

R70_107 V70 V107 4088.666360863932
L70_107 V70 V107 9.018358502626171e-13
C70_107 V70 V107 7.81957543464468e-19

R70_108 V70 V108 -2756.1247509772866
L70_108 V70 V108 -9.029855147859756e-13
C70_108 V70 V108 -7.279105621444102e-19

R70_109 V70 V109 -6797.6587919577005
L70_109 V70 V109 -4.2921824315857796e-12
C70_109 V70 V109 -1.6856715488429463e-19

R70_110 V70 V110 -2859.0449750235107
L70_110 V70 V110 -7.51448956812362e-13
C70_110 V70 V110 -9.445853428095724e-19

R70_111 V70 V111 -6466.758890874116
L70_111 V70 V111 -1.1831920935283866e-12
C70_111 V70 V111 -5.151775663136423e-19

R70_112 V70 V112 7946.105508128882
L70_112 V70 V112 8.145383244340918e-13
C70_112 V70 V112 7.085168707961185e-19

R70_113 V70 V113 12825.179280856377
L70_113 V70 V113 1.9825621424293587e-12
C70_113 V70 V113 2.6332830342937776e-19

R70_114 V70 V114 5946.181982895699
L70_114 V70 V114 1.121620426014528e-12
C70_114 V70 V114 5.911579448113397e-19

R70_115 V70 V115 9381.938724693138
L70_115 V70 V115 1.5915777379899255e-12
C70_115 V70 V115 4.1718123543475564e-19

R70_116 V70 V116 -5675.239233164708
L70_116 V70 V116 -1.2952149278454527e-12
C70_116 V70 V116 -4.324726263870661e-19

R70_117 V70 V117 -4009.2660700634115
L70_117 V70 V117 -2.3115811310437887e-12
C70_117 V70 V117 -3.2368204072853434e-19

R70_118 V70 V118 -27152.95135192854
L70_118 V70 V118 -1.345696590607022e-12
C70_118 V70 V118 -4.581120633830168e-19

R70_119 V70 V119 -6446.658803996025
L70_119 V70 V119 -9.45172793623488e-13
C70_119 V70 V119 -6.625608954212958e-19

R70_120 V70 V120 -4210.403130816789
L70_120 V70 V120 1.0213049205805818e-11
C70_120 V70 V120 -2.191055555075049e-19

R70_121 V70 V121 -9445.980464179213
L70_121 V70 V121 3.1678549577699277e-12
C70_121 V70 V121 1.2510581677321972e-19

R70_122 V70 V122 -3102.449725651565
L70_122 V70 V122 1.5923210678581873e-12
C70_122 V70 V122 9.497650777441803e-21

R70_123 V70 V123 -8781.576651992335
L70_123 V70 V123 -4.1053925112179023e-11
C70_123 V70 V123 -7.684803088007047e-20

R70_124 V70 V124 -19901.737788983603
L70_124 V70 V124 -3.291901582108498e-12
C70_124 V70 V124 -1.7078653649703288e-19

R70_125 V70 V125 81859.25748724655
L70_125 V70 V125 -6.542698361094907e-12
C70_125 V70 V125 -9.867533389603716e-20

R70_126 V70 V126 2929.7032447264755
L70_126 V70 V126 -1.6572615781352002e-12
C70_126 V70 V126 1.2326542548480647e-19

R70_127 V70 V127 -3842.7566835216567
L70_127 V70 V127 1.6154450834605854e-12
C70_127 V70 V127 -1.4895845312930225e-20

R70_128 V70 V128 -10419.178472935084
L70_128 V70 V128 1.103765909592844e-11
C70_128 V70 V128 -2.812950371984918e-20

R70_129 V70 V129 -7055.914934209397
L70_129 V70 V129 1.32399234145811e-11
C70_129 V70 V129 -7.407793067966506e-20

R70_130 V70 V130 -10550.962480549451
L70_130 V70 V130 -2.5377051512270854e-12
C70_130 V70 V130 -2.3570659741639595e-19

R70_131 V70 V131 8286.183034530624
L70_131 V70 V131 5.197180413772634e-12
C70_131 V70 V131 2.2265801331462313e-19

R70_132 V70 V132 12906.966485418843
L70_132 V70 V132 -5.359072918673542e-12
C70_132 V70 V132 -5.484395850523385e-21

R70_133 V70 V133 4725.239972002709
L70_133 V70 V133 1.7863839078158003e-12
C70_133 V70 V133 3.6591621131544977e-19

R70_134 V70 V134 4577.739304500045
L70_134 V70 V134 -2.1698404027271172e-11
C70_134 V70 V134 -9.561143134132407e-21

R70_135 V70 V135 -5552.657027583278
L70_135 V70 V135 2.8442544737772064e-12
C70_135 V70 V135 -6.523030561865966e-20

R70_136 V70 V136 -43317.68442995506
L70_136 V70 V136 7.596234914636138e-10
C70_136 V70 V136 -3.2507832684109454e-20

R70_137 V70 V137 -15400.390556073258
L70_137 V70 V137 -3.437827724979547e-12
C70_137 V70 V137 -1.9609156268504765e-19

R70_138 V70 V138 3789.962851717165
L70_138 V70 V138 -1.4856413589279654e-12
C70_138 V70 V138 -9.670138400711091e-20

R70_139 V70 V139 -2940.540313220949
L70_139 V70 V139 1.1157198289986609e-12
C70_139 V70 V139 1.497500411617574e-19

R70_140 V70 V140 5959.171502801462
L70_140 V70 V140 -2.8831247065360834e-12
C70_140 V70 V140 -6.98191133561539e-20

R70_141 V70 V141 37672.67279075651
L70_141 V70 V141 -4.308547674588366e-12
C70_141 V70 V141 -3.618831278053486e-20

R70_142 V70 V142 9780.396449712376
L70_142 V70 V142 -2.6554906691898737e-12
C70_142 V70 V142 -1.1588802711811667e-19

R70_143 V70 V143 13458.999463451431
L70_143 V70 V143 -5.331667755410171e-12
C70_143 V70 V143 1.1128092091127756e-20

R70_144 V70 V144 46595.78337062649
L70_144 V70 V144 3.111421961851698e-12
C70_144 V70 V144 5.666707080861736e-20

R71_71 V71 0 -907.7125972505695
L71_71 V71 0 -1.9165597644907517e-13
C71_71 V71 0 -1.9638817471114922e-19

R71_72 V71 V72 2317.8647334416974
L71_72 V71 V72 1.7902536861860683e-12
C71_72 V71 V72 5.890147872448001e-20

R71_73 V71 V73 1992.1386943197672
L71_73 V71 V73 1.2068047084923452e-12
C71_73 V71 V73 4.0511674366294826e-20

R71_74 V71 V74 2187.925614567915
L71_74 V71 V74 3.678846312612973e-12
C71_74 V71 V74 -2.5036139668504066e-20

R71_75 V71 V75 -9251.893657102106
L71_75 V71 V75 1.6688022013418182e-12
C71_75 V71 V75 2.7297239775265216e-19

R71_76 V71 V76 10714.388552768347
L71_76 V71 V76 -3.370131376165265e-12
C71_76 V71 V76 -2.5751355222368174e-19

R71_77 V71 V77 9908.306123756358
L71_77 V71 V77 -1.5698292335348285e-11
C71_77 V71 V77 -6.268946782424867e-20

R71_78 V71 V78 6697.761455244363
L71_78 V71 V78 -1.1886958481244047e-11
C71_78 V71 V78 -2.203967284259718e-19

R71_79 V71 V79 5631.868494736699
L71_79 V71 V79 -1.5094175353124864e-12
C71_79 V71 V79 -4.206869029400213e-19

R71_80 V71 V80 -22552.96852298855
L71_80 V71 V80 2.1896400358948802e-12
C71_80 V71 V80 3.475816301041025e-19

R71_81 V71 V81 -9725.922085370708
L71_81 V71 V81 -4.778597823835869e-12
C71_81 V71 V81 3.3952628638066994e-20

R71_82 V71 V82 8923.049912274493
L71_82 V71 V82 1.1423599470769283e-12
C71_82 V71 V82 2.732173032837443e-19

R71_83 V71 V83 -4061.4633626740087
L71_83 V71 V83 -3.322574581485278e-12
C71_83 V71 V83 2.918553112849934e-19

R71_84 V71 V84 6561.736467194276
L71_84 V71 V84 -3.026421221668441e-11
C71_84 V71 V84 -1.0102584381225762e-19

R71_85 V71 V85 -51596.62047694124
L71_85 V71 V85 -1.865630254553053e-12
C71_85 V71 V85 -2.7067653867637444e-19

R71_86 V71 V86 4317.502865581442
L71_86 V71 V86 2.9746345303581262e-12
C71_86 V71 V86 -4.7819937884204327e-20

R71_87 V71 V87 -12646.739789322899
L71_87 V71 V87 -1.9610872776186383e-12
C71_87 V71 V87 -2.0771525096628872e-19

R71_88 V71 V88 785170.4294214272
L71_88 V71 V88 -1.3808961681140929e-11
C71_88 V71 V88 -2.314727254400169e-20

R71_89 V71 V89 18183.948862004523
L71_89 V71 V89 2.7061301174587054e-12
C71_89 V71 V89 7.333020506361505e-20

R71_90 V71 V90 93531.28023364197
L71_90 V71 V90 1.674769744191976e-12
C71_90 V71 V90 3.960592500285233e-19

R71_91 V71 V91 23968.56584814248
L71_91 V71 V91 3.010738789470459e-12
C71_91 V71 V91 2.138965022830599e-19

R71_92 V71 V92 12906.716775661898
L71_92 V71 V92 2.9741790943128357e-12
C71_92 V71 V92 1.6621881973754592e-19

R71_93 V71 V93 -43720.370833048066
L71_93 V71 V93 -5.1636703793535515e-12
C71_93 V71 V93 -8.081359653152018e-20

R71_94 V71 V94 -9071.010905467963
L71_94 V71 V94 -9.66022345338369e-12
C71_94 V71 V94 4.178863334003796e-20

R71_95 V71 V95 26923.687495096503
L71_95 V71 V95 5.392036857910805e-12
C71_95 V71 V95 1.3150684989549152e-19

R71_96 V71 V96 11112.145195467183
L71_96 V71 V96 3.858334414014908e-12
C71_96 V71 V96 1.1246015048110582e-19

R71_97 V71 V97 20842.340010990058
L71_97 V71 V97 2.4186659054692648e-12
C71_97 V71 V97 1.276190568369931e-19

R71_98 V71 V98 -20304.222050648514
L71_98 V71 V98 2.2309026760366658e-12
C71_98 V71 V98 1.9369968910100518e-19

R71_99 V71 V99 -5595.83953583397
L71_99 V71 V99 -2.5804319208910458e-12
C71_99 V71 V99 -5.354768837297726e-20

R71_100 V71 V100 164460.51840044121
L71_100 V71 V100 3.993995820611731e-11
C71_100 V71 V100 3.4782166474740464e-20

R71_101 V71 V101 308407.84142001544
L71_101 V71 V101 3.7415773485101564e-12
C71_101 V71 V101 1.06844298816411e-19

R71_102 V71 V102 4373.776685143219
L71_102 V71 V102 6.285237001357028e-13
C71_102 V71 V102 8.21547147514707e-19

R71_103 V71 V103 -9398.976856464164
L71_103 V71 V103 -1.2890716949597668e-12
C71_103 V71 V103 -4.996675220931588e-19

R71_104 V71 V104 35395.80703383609
L71_104 V71 V104 8.807709908855507e-12
C71_104 V71 V104 8.418472846530216e-20

R71_105 V71 V105 -8256.11154388126
L71_105 V71 V105 -1.4224078114377748e-12
C71_105 V71 V105 -3.2918594587324884e-19

R71_106 V71 V106 3494.365715479615
L71_106 V71 V106 9.163920804995768e-13
C71_106 V71 V106 5.830040585880726e-19

R71_107 V71 V107 4686.44660955551
L71_107 V71 V107 7.288924696774335e-13
C71_107 V71 V107 7.059216761889933e-19

R71_108 V71 V108 -3445.8403836236253
L71_108 V71 V108 -9.118785159917595e-13
C71_108 V71 V108 -5.166152498554011e-19

R71_109 V71 V109 -6459.54019675659
L71_109 V71 V109 -2.065578905745895e-12
C71_109 V71 V109 -2.2819525631475776e-19

R71_110 V71 V110 -16197.671929068565
L71_110 V71 V110 -1.793007037417139e-12
C71_110 V71 V110 -4.2308709672286496e-19

R71_111 V71 V111 -4465.361382437694
L71_111 V71 V111 -1.2805411953915936e-12
C71_111 V71 V111 -3.1598193746718163e-19

R71_112 V71 V112 8462.817475225678
L71_112 V71 V112 9.39016932368166e-13
C71_112 V71 V112 4.043570401443103e-19

R71_113 V71 V113 14727.524774032778
L71_113 V71 V113 1.8615214493249446e-12
C71_113 V71 V113 2.0470306815124444e-19

R71_114 V71 V114 6860.208088238452
L71_114 V71 V114 1.938755887072569e-12
C71_114 V71 V114 1.9085428225755043e-19

R71_115 V71 V115 8604.834309761338
L71_115 V71 V115 1.2362090521922282e-12
C71_115 V71 V115 4.054009410576387e-19

R71_116 V71 V116 -5463.176171077807
L71_116 V71 V116 -1.3581807181585301e-12
C71_116 V71 V116 -3.246384451301153e-19

R71_117 V71 V117 -25927.35854609516
L71_117 V71 V117 -2.2884871370462386e-12
C71_117 V71 V117 -2.9825565711296006e-19

R71_118 V71 V118 -11303.72552603524
L71_118 V71 V118 -2.009990941819366e-12
C71_118 V71 V118 -2.1617718115530113e-19

R71_119 V71 V119 -5186.891107253534
L71_119 V71 V119 -1.596982548005483e-12
C71_119 V71 V119 -2.453547718391151e-19

R71_120 V71 V120 3185.082195907427
L71_120 V71 V120 1.8745344774424303e-12
C71_120 V71 V120 -9.494023912215443e-20

R71_121 V71 V121 -8210.580379083633
L71_121 V71 V121 4.059065126104606e-12
C71_121 V71 V121 7.909687853700543e-20

R71_122 V71 V122 5436.383804065859
L71_122 V71 V122 9.84767846923438e-13
C71_122 V71 V122 -5.436432181420691e-21

R71_123 V71 V123 14009.417164278226
L71_123 V71 V123 5.335317407485604e-12
C71_123 V71 V123 -5.178927676456076e-20

R71_124 V71 V124 -24996.16599058695
L71_124 V71 V124 -4.688753796510489e-12
C71_124 V71 V124 -7.452413564266281e-20

R71_125 V71 V125 5093.349149630496
L71_125 V71 V125 -2.234515712636436e-09
C71_125 V71 V125 -5.372064761533281e-20

R71_126 V71 V126 -2498.097435055343
L71_126 V71 V126 -8.50464243340806e-13
C71_126 V71 V126 9.579508511891222e-20

R71_127 V71 V127 2875.5009955907353
L71_127 V71 V127 1.0028273095338633e-12
C71_127 V71 V127 9.001139491267874e-21

R71_128 V71 V128 -59176.12596746523
L71_128 V71 V128 7.74306431807785e-11
C71_128 V71 V128 -4.5482517939051226e-20

R71_129 V71 V129 7223.9585387678435
L71_129 V71 V129 3.2807045757251342e-12
C71_129 V71 V129 -4.679959638608159e-20

R71_130 V71 V130 -4023.493639125091
L71_130 V71 V130 -1.283350669293758e-12
C71_130 V71 V130 -1.8945185187294556e-19

R71_131 V71 V131 -14161.902589140904
L71_131 V71 V131 -4.270592569944046e-11
C71_131 V71 V131 1.755966496687687e-19

R71_132 V71 V132 -14106.086185030295
L71_132 V71 V132 -3.2092992448100738e-12
C71_132 V71 V132 -4.721376207612374e-20

R71_133 V71 V133 9135.530314808704
L71_133 V71 V133 4.43767101239498e-12
C71_133 V71 V133 1.3612733897203934e-19

R71_134 V71 V134 26188.448363706197
L71_134 V71 V134 -9.241234855403351e-12
C71_134 V71 V134 2.8124113390238123e-20

R71_135 V71 V135 4016.4556152143705
L71_135 V71 V135 1.6409398472189245e-12
C71_135 V71 V135 -6.167219309987149e-20

R71_136 V71 V136 1151586.9973628279
L71_136 V71 V136 1.5441617091276198e-11
C71_136 V71 V136 4.379380778942979e-20

R71_137 V71 V137 14179.651633836698
L71_137 V71 V137 -5.9458634562843805e-12
C71_137 V71 V137 -4.651537502339139e-20

R71_138 V71 V138 -3044.413816531194
L71_138 V71 V138 -8.044236886096888e-13
C71_138 V71 V138 -7.273830900413192e-20

R71_139 V71 V139 2386.3477643201713
L71_139 V71 V139 7.17717889210453e-13
C71_139 V71 V139 7.75354867979454e-20

R71_140 V71 V140 -7800.840355705225
L71_140 V71 V140 -2.220515983596261e-12
C71_140 V71 V140 -2.2609337741549748e-20

R71_141 V71 V141 -15789.271994030985
L71_141 V71 V141 -3.351627775432005e-12
C71_141 V71 V141 -1.5146720373623448e-20

R71_142 V71 V142 -5697.822378122313
L71_142 V71 V142 -1.788389090342175e-12
C71_142 V71 V142 -7.205516585910971e-20

R71_143 V71 V143 -4910.818755040203
L71_143 V71 V143 -2.000059486892809e-12
C71_143 V71 V143 -4.911152894374716e-20

R71_144 V71 V144 7282.381168919682
L71_144 V71 V144 2.650751720377296e-12
C71_144 V71 V144 4.185622190119523e-20

R72_72 V72 0 -84.83255555757259
L72_72 V72 0 -1.574628290693109e-13
C72_72 V72 0 -2.50152011293116e-20

R72_73 V72 V73 -4537.520993777357
L72_73 V72 V73 -1.1658543771423437e-12
C72_73 V72 V73 3.607784883488254e-21

R72_74 V72 V74 -2557.8812868739433
L72_74 V72 V74 -1.2646972483233415e-12
C72_74 V72 V74 2.9345746590651836e-20

R72_75 V72 V75 2701.400647135944
L72_75 V72 V75 1.752092361876595e-12
C72_75 V72 V75 6.727776214212829e-21

R72_76 V72 V76 4546.943095190125
L72_76 V72 V76 1.187919115325462e-12
C72_76 V72 V76 5.236545402011483e-20

R72_77 V72 V77 67055.5262674001
L72_77 V72 V77 3.1545462404508206e-12
C72_77 V72 V77 3.2012639375284096e-21

R72_78 V72 V78 -7142.519369504539
L72_78 V72 V78 6.122044918902432e-11
C72_78 V72 V78 -4.4256211718413136e-20

R72_79 V72 V79 -6515.424307316106
L72_79 V72 V79 -6.03027378003874e-12
C72_79 V72 V79 8.305577013690172e-20

R72_80 V72 V80 -38398.52761175339
L72_80 V72 V80 -2.6896538219226673e-12
C72_80 V72 V80 -1.2426993448612102e-19

R72_81 V72 V81 24548.809304244733
L72_81 V72 V81 -5.88136921326332e-12
C72_81 V72 V81 6.424528092661353e-20

R72_82 V72 V82 9343.853814156355
L72_82 V72 V82 1.0835521384612624e-12
C72_82 V72 V82 3.043730864328563e-19

R72_83 V72 V83 6853.627055253396
L72_83 V72 V83 2.3402140901784905e-12
C72_83 V72 V83 1.779055231851324e-19

R72_84 V72 V84 -13794.916517503098
L72_84 V72 V84 -2.24558883148639e-12
C72_84 V72 V84 3.7211618430952654e-20

R72_85 V72 V85 -7157.970829005309
L72_85 V72 V85 -1.980156724578708e-12
C72_85 V72 V85 -1.8604203520153445e-21

R72_86 V72 V86 -5739.20129935475
L72_86 V72 V86 -1.5617241625212923e-12
C72_86 V72 V86 -1.2725758330808156e-19

R72_87 V72 V87 -30877.95753724556
L72_87 V72 V87 -3.9926788192691805e-12
C72_87 V72 V87 -1.3149171162843842e-19

R72_88 V72 V88 -2284647.419902593
L72_88 V72 V88 1.7584639700053707e-11
C72_88 V72 V88 -3.43296144234285e-20

R72_89 V72 V89 12996.604377223213
L72_89 V72 V89 2.63566504908716e-12
C72_89 V72 V89 4.5175577665490065e-20

R72_90 V72 V90 -279958.9109324073
L72_90 V72 V90 -1.0368786809531308e-11
C72_90 V72 V90 -1.0331081825175178e-19

R72_91 V72 V91 10550.464426956412
L72_91 V72 V91 1.3870782230958072e-12
C72_91 V72 V91 3.245524481542636e-19

R72_92 V72 V92 43246.324145839186
L72_92 V72 V92 6.123438914495733e-12
C72_92 V72 V92 4.359229028859454e-20

R72_93 V72 V93 -8282.387906350072
L72_93 V72 V93 -3.001299389811363e-11
C72_93 V72 V93 -6.3245807129488724e-21

R72_94 V72 V94 -98875.59816647711
L72_94 V72 V94 -4.1882197535486876e-12
C72_94 V72 V94 -8.65024124530781e-20

R72_95 V72 V95 10413.196590678683
L72_95 V72 V95 2.699516467319779e-12
C72_95 V72 V95 1.6944950752374102e-19

R72_96 V72 V96 29295.178586080245
L72_96 V72 V96 -9.15185423552156e-12
C72_96 V72 V96 -5.35545160142587e-20

R72_97 V72 V97 -4239.678845768272
L72_97 V72 V97 -2.864390419383995e-12
C72_97 V72 V97 -1.2416239385871098e-19

R72_98 V72 V98 -3752.1858693765253
L72_98 V72 V98 4.699676634325677e-12
C72_98 V72 V98 8.049100114112506e-20

R72_99 V72 V99 -517484.0821311001
L72_99 V72 V99 1.3901031890255523e-11
C72_99 V72 V99 1.4890054634475593e-21

R72_100 V72 V100 30201.377697254746
L72_100 V72 V100 -1.8925087089596424e-11
C72_100 V72 V100 -7.486498047766419e-21

R72_101 V72 V101 -13629.970879870265
L72_101 V72 V101 2.8744039082564817e-12
C72_101 V72 V101 8.706111953597451e-20

R72_102 V72 V102 -12075.910702991669
L72_102 V72 V102 -2.2112982574532758e-11
C72_102 V72 V102 -8.232829289733505e-20

R72_103 V72 V103 -16783.419657768256
L72_103 V72 V103 3.5043264381600447e-12
C72_103 V72 V103 1.3147088907095944e-19

R72_104 V72 V104 41987.928931873816
L72_104 V72 V104 -3.3377857014880026e-12
C72_104 V72 V104 -1.6805449703852845e-19

R72_105 V72 V105 8833.362834787442
L72_105 V72 V105 -5.188131511501046e-12
C72_105 V72 V105 -8.322462159290443e-20

R72_106 V72 V106 3455.030774892808
L72_106 V72 V106 2.0057913498552047e-12
C72_106 V72 V106 2.2093165221959337e-19

R72_107 V72 V107 -11107.624285416287
L72_107 V72 V107 -5.753461203366266e-12
C72_107 V72 V107 -5.086533804738386e-20

R72_108 V72 V108 -33889.73430630583
L72_108 V72 V108 8.04798940065555e-12
C72_108 V72 V108 1.0109168411944585e-19

R72_109 V72 V109 -14059.982666800728
L72_109 V72 V109 -1.0315101674016246e-11
C72_109 V72 V109 -7.090914610604796e-20

R72_110 V72 V110 -16759.022910968808
L72_110 V72 V110 -2.021507626655749e-12
C72_110 V72 V110 -2.096981213409748e-19

R72_111 V72 V111 -43966.40611896274
L72_111 V72 V111 2.660066350742858e-11
C72_111 V72 V111 -2.4174283737195202e-20

R72_112 V72 V112 -6745.736499152384
L72_112 V72 V112 9.606422310232627e-12
C72_112 V72 V112 2.4527343568992312e-20

R72_113 V72 V113 -44880.57338709549
L72_113 V72 V113 1.0515465384388598e-11
C72_113 V72 V113 6.30778738701969e-20

R72_114 V72 V114 17488.24371604215
L72_114 V72 V114 3.896491833505691e-12
C72_114 V72 V114 1.6297401655642562e-19

R72_115 V72 V115 -42713.76712495045
L72_115 V72 V115 -9.950057055704775e-12
C72_115 V72 V115 -4.576908014511159e-20

R72_116 V72 V116 48956.11286339464
L72_116 V72 V116 1.2413087633951668e-11
C72_116 V72 V116 8.14421513204672e-20

R72_117 V72 V117 -9010.978945978064
L72_117 V72 V117 -1.2875327062239353e-11
C72_117 V72 V117 2.2621052519046273e-21

R72_118 V72 V118 8785.600914821316
L72_118 V72 V118 -4.836138667384985e-12
C72_118 V72 V118 -1.327093443450507e-19

R72_119 V72 V119 -58809.72292666111
L72_119 V72 V119 -4.5573722529223355e-12
C72_119 V72 V119 -1.3247278966676974e-19

R72_120 V72 V120 -8813.484432825495
L72_120 V72 V120 -4.4648971674626354e-12
C72_120 V72 V120 9.494178503412689e-22

R72_121 V72 V121 -5238.537453662253
L72_121 V72 V121 9.189005363627105e-12
C72_121 V72 V121 2.817083849040358e-20

R72_122 V72 V122 -3297.130388482014
L72_122 V72 V122 -5.582179678976814e-12
C72_122 V72 V122 -1.3196713737497953e-21

R72_123 V72 V123 -16329.317294146445
L72_123 V72 V123 -6.8132273526093175e-12
C72_123 V72 V123 -3.8010613875100614e-20

R72_124 V72 V124 -3515727.789299826
L72_124 V72 V124 2.2744374220744577e-11
C72_124 V72 V124 -1.0528524066734974e-20

R72_125 V72 V125 6781.460770340906
L72_125 V72 V125 -8.981905884595631e-12
C72_125 V72 V125 4.089999105565295e-21

R72_126 V72 V126 4056.721016316098
L72_126 V72 V126 3.3484536868658688e-12
C72_126 V72 V126 3.8603048584127386e-21

R72_127 V72 V127 -4375.539919755004
L72_127 V72 V127 -5.116945868960596e-12
C72_127 V72 V127 -2.9214597890606666e-21

R72_128 V72 V128 -14445.591109871053
L72_128 V72 V128 -8.470530292878867e-11
C72_128 V72 V128 -5.934835397524636e-21

R72_129 V72 V129 -13274.720539550613
L72_129 V72 V129 -1.0496916098335641e-11
C72_129 V72 V129 -1.0732651651784439e-20

R72_130 V72 V130 -26723.481559231004
L72_130 V72 V130 4.727722751443536e-12
C72_130 V72 V130 2.776972656875314e-20

R72_131 V72 V131 -131666.05398101397
L72_131 V72 V131 1.2102692465035469e-11
C72_131 V72 V131 3.510841261504464e-21

R72_132 V72 V132 10653.164759982054
L72_132 V72 V132 8.795405027595219e-12
C72_132 V72 V132 4.830586398074811e-20

R72_133 V72 V133 8378.147961565879
L72_133 V72 V133 5.175306124716788e-12
C72_133 V72 V133 8.622326713173054e-20

R72_134 V72 V134 4499.354826304519
L72_134 V72 V134 1.1592371659909164e-11
C72_134 V72 V134 -1.1784562680735938e-20

R72_135 V72 V135 -7710.164671340921
L72_135 V72 V135 -7.28527236725913e-12
C72_135 V72 V135 1.4772514017500343e-20

R72_136 V72 V136 -26058.743285783086
L72_136 V72 V136 -1.0216427348254449e-11
C72_136 V72 V136 -5.63919221305165e-20

R72_137 V72 V137 50455.86168645323
L72_137 V72 V137 -9.781871142187324e-12
C72_137 V72 V137 -5.3854486976832273e-20

R72_138 V72 V138 5044.616434583964
L72_138 V72 V138 3.575613056746301e-12
C72_138 V72 V138 -8.998182662057183e-21

R72_139 V72 V139 -3164.9297975372624
L72_139 V72 V139 -2.9965419499143658e-12
C72_139 V72 V139 2.955360108958916e-21

R72_140 V72 V140 4107.902665138844
L72_140 V72 V140 2.2758427224581043e-11
C72_140 V72 V140 -1.374046633629915e-20

R72_141 V72 V141 38730.09921604416
L72_141 V72 V141 2.0003745316973655e-11
C72_141 V72 V141 -1.7687533888230013e-20

R72_142 V72 V142 8842.492256938027
L72_142 V72 V142 3.809846421841964e-11
C72_142 V72 V142 -2.2071513985645033e-20

R72_143 V72 V143 18920.81975382104
L72_143 V72 V143 5.393256933741876e-12
C72_143 V72 V143 3.6599517776390126e-20

R72_144 V72 V144 -22092.64776181941
L72_144 V72 V144 3.898338263981872e-11
C72_144 V72 V144 2.745060562063496e-20

R73_73 V73 0 1908.850639001822
L73_73 V73 0 1.8019880451479343e-13
C73_73 V73 0 9.79410100399271e-19

R73_74 V73 V74 -4361.624599534928
L73_74 V73 V74 -3.0929008977316555e-12
C73_74 V73 V74 3.581199649618978e-20

R73_75 V73 V75 9854.524491314669
L73_75 V73 V75 3.4640665629575155e-12
C73_75 V73 V75 3.8931788443241746e-20

R73_76 V73 V76 -11539.59245324853
L73_76 V73 V76 2.2919886744238394e-11
C73_76 V73 V76 -4.841160229778962e-20

R73_77 V73 V77 148624.57057749017
L73_77 V73 V77 2.2518610703623475e-12
C73_77 V73 V77 1.64437068415412e-19

R73_78 V73 V78 -9782.41258123366
L73_78 V73 V78 -1.4464147577753224e-11
C73_78 V73 V78 -7.499932913063873e-20

R73_79 V73 V79 -8362.159765038296
L73_79 V73 V79 -5.818652446576878e-12
C73_79 V73 V79 5.862584071890273e-20

R73_80 V73 V80 6459.8202490665235
L73_80 V73 V80 3.664753517233905e-12
C73_80 V73 V80 1.5081650428776908e-19

R73_81 V73 V81 -9361.748661979716
L73_81 V73 V81 -1.1279586289015442e-12
C73_81 V73 V81 -4.473189641545328e-19

R73_82 V73 V82 21595.041232251893
L73_82 V73 V82 4.9851072842072884e-12
C73_82 V73 V82 9.328791774219542e-20

R73_83 V73 V83 5677.835998003847
L73_83 V73 V83 2.224769132031073e-12
C73_83 V73 V83 1.7169760046280498e-19

R73_84 V73 V84 -11424.180988193239
L73_84 V73 V84 -2.648041762075333e-12
C73_84 V73 V84 3.210738202509947e-20

R73_85 V73 V85 -11318.984411491754
L73_85 V73 V85 -2.039084392941955e-12
C73_85 V73 V85 -1.0162599853498209e-19

R73_86 V73 V86 -7294.7165127713515
L73_86 V73 V86 -3.1548709822931586e-12
C73_86 V73 V86 -4.641788607985292e-20

R73_87 V73 V87 -19525.60522588794
L73_87 V73 V87 -8.782143736510008e-12
C73_87 V73 V87 -6.667620632796364e-20

R73_88 V73 V88 -97669.15535345236
L73_88 V73 V88 -1.29239031580995e-11
C73_88 V73 V88 -9.812082981024193e-20

R73_89 V73 V89 12793.501154353187
L73_89 V73 V89 2.6830166353778472e-12
C73_89 V73 V89 1.3597946706730682e-19

R73_90 V73 V90 51435.92595841304
L73_90 V73 V90 1.41453406509696e-11
C73_90 V73 V90 -5.3802475141017853e-20

R73_91 V73 V91 163777.84678885108
L73_91 V73 V91 -1.995144357859909e-11
C73_91 V73 V91 -9.779113623084355e-21

R73_92 V73 V92 9201.909921825305
L73_92 V73 V92 1.839940715579517e-12
C73_92 V73 V92 3.1305810306542543e-19

R73_93 V73 V93 21276.204454687377
L73_93 V73 V93 -2.8035902108011855e-11
C73_93 V73 V93 -1.3268299653494058e-21

R73_94 V73 V94 57960.25271613009
L73_94 V73 V94 -3.0642159466648144e-12
C73_94 V73 V94 -2.1332419895309043e-19

R73_95 V73 V95 23272.346119148082
L73_95 V73 V95 2.5847143777015403e-11
C73_95 V73 V95 3.2571725987658753e-20

R73_96 V73 V96 7199.776536519425
L73_96 V73 V96 1.5072146626563122e-12
C73_96 V73 V96 3.9036449007013695e-19

R73_97 V73 V97 -7801.9697066418685
L73_97 V73 V97 -5.077044572373844e-12
C73_97 V73 V97 -1.368481970154296e-19

R73_98 V73 V98 -29833.873697584986
L73_98 V73 V98 3.078483963342843e-12
C73_98 V73 V98 1.3109994689973984e-19

R73_99 V73 V99 22045.383508393523
L73_99 V73 V99 -2.7969547690194584e-11
C73_99 V73 V99 -5.0381287745244535e-20

R73_100 V73 V100 -32211.274726116437
L73_100 V73 V100 -4.074604360838503e-12
C73_100 V73 V100 -1.7184544199173917e-19

R73_101 V73 V101 10525.648043243464
L73_101 V73 V101 2.210833080186348e-12
C73_101 V73 V101 2.0618711192505002e-19

R73_102 V73 V102 -27685.49376647471
L73_102 V73 V102 7.84886138807341e-12
C73_102 V73 V102 -5.1945194109836846e-20

R73_103 V73 V103 -19486.114308444485
L73_103 V73 V103 -4.715482005315124e-10
C73_103 V73 V103 4.97828435366194e-20

R73_104 V73 V104 8221.296576230428
L73_104 V73 V104 1.8256835552529907e-12
C73_104 V73 V104 3.4524769153335026e-19

R73_105 V73 V105 195652.19648211356
L73_105 V73 V105 -3.131264890778041e-12
C73_105 V73 V105 -2.0645041636913634e-19

R73_106 V73 V106 9228.705769226342
L73_106 V73 V106 3.5919856349940368e-12
C73_106 V73 V106 1.8230053608845117e-19

R73_107 V73 V107 -28353.04446830883
L73_107 V73 V107 -1.8259087620030027e-11
C73_107 V73 V107 -8.745893847551063e-20

R73_108 V73 V108 -12569.110006134906
L73_108 V73 V108 -3.1755113735334177e-12
C73_108 V73 V108 -1.518450297939356e-19

R73_109 V73 V109 25712.29829144257
L73_109 V73 V109 2.227671115204871e-12
C73_109 V73 V109 3.2507797262178303e-19

R73_110 V73 V110 -9685.510746935151
L73_110 V73 V110 -2.9101556600207734e-12
C73_110 V73 V110 -1.7060940738658078e-19

R73_111 V73 V111 -42013.33008652629
L73_111 V73 V111 -2.5473448620982946e-11
C73_111 V73 V111 -5.853818107782868e-20

R73_112 V73 V112 -14238.496329214091
L73_112 V73 V112 3.969448729758969e-12
C73_112 V73 V112 8.212456446256105e-20

R73_113 V73 V113 -22243.04939760193
L73_113 V73 V113 -2.4378110123487324e-11
C73_113 V73 V113 -9.214711208468797e-20

R73_114 V73 V114 -26970.488391883442
L73_114 V73 V114 8.804841754160351e-12
C73_114 V73 V114 1.0246117896249943e-19

R73_115 V73 V115 -44126.44864438964
L73_115 V73 V115 -1.3251004263831884e-11
C73_115 V73 V115 -4.4068391709845614e-20

R73_116 V73 V116 -86883.61433488582
L73_116 V73 V116 -5.422223301722304e-12
C73_116 V73 V116 -9.041280260613037e-20

R73_117 V73 V117 -32452.978928507768
L73_117 V73 V117 -1.4730576779871342e-11
C73_117 V73 V117 4.112731048449361e-20

R73_118 V73 V118 17467.331480138648
L73_118 V73 V118 3.6159671817704533e-11
C73_118 V73 V118 3.642660429595058e-20

R73_119 V73 V119 -27857.020733998215
L73_119 V73 V119 -8.019867902739956e-12
C73_119 V73 V119 -1.4196736535065284e-19

R73_120 V73 V120 -8074.245922266813
L73_120 V73 V120 -2.8939791686556936e-12
C73_120 V73 V120 -8.51285640331829e-20

R73_121 V73 V121 -7007.002575863281
L73_121 V73 V121 8.525366584418888e-12
C73_121 V73 V121 7.184393842040528e-21

R73_122 V73 V122 -3061.6176785921225
L73_122 V73 V122 -1.3026063986620629e-09
C73_122 V73 V122 3.677013465523956e-20

R73_123 V73 V123 -7595.76456612182
L73_123 V73 V123 -3.6019216030541035e-11
C73_123 V73 V123 1.8935635559471306e-20

R73_124 V73 V124 -17013.668230144856
L73_124 V73 V124 -8.971282759750213e-12
C73_124 V73 V124 -8.65748134099438e-20

R73_125 V73 V125 11915.27364312534
L73_125 V73 V125 -4.231010429030987e-12
C73_125 V73 V125 -8.57132317688652e-21

R73_126 V73 V126 3098.2546013633855
L73_126 V73 V126 4.543646335027183e-12
C73_126 V73 V126 -2.218725542467591e-21

R73_127 V73 V127 -4844.339673026617
L73_127 V73 V127 -6.114814283739548e-12
C73_127 V73 V127 -1.4348078613484223e-20

R73_128 V73 V128 -19938.79176488628
L73_128 V73 V128 5.565295134425065e-11
C73_128 V73 V128 -2.572899797633737e-20

R73_129 V73 V129 -5931.959973203691
L73_129 V73 V129 -6.791224148600727e-12
C73_129 V73 V129 -3.9416368998354966e-20

R73_130 V73 V130 8043.979615976163
L73_130 V73 V130 2.6171776687894845e-11
C73_130 V73 V130 -5.2330283632259973e-20

R73_131 V73 V131 7009.706009936145
L73_131 V73 V131 1.8042552425955444e-11
C73_131 V73 V131 -2.3782612773943656e-20

R73_132 V73 V132 30060.512529550037
L73_132 V73 V132 -8.609841386165435e-12
C73_132 V73 V132 -8.408881462092119e-20

R73_133 V73 V133 12888.305684355193
L73_133 V73 V133 8.998551146353759e-12
C73_133 V73 V133 7.978766955037473e-20

R73_134 V73 V134 13305.905032002674
L73_134 V73 V134 1.1578501670603721e-10
C73_134 V73 V134 -4.5481279482419554e-21

R73_135 V73 V135 -6427.229639108199
L73_135 V73 V135 -7.714421296910115e-12
C73_135 V73 V135 -9.298099254870793e-21

R73_136 V73 V136 35149.88414219878
L73_136 V73 V136 6.96850287139613e-12
C73_136 V73 V136 7.73348767071996e-20

R73_137 V73 V137 34551.13191966652
L73_137 V73 V137 -7.008901451272827e-12
C73_137 V73 V137 -6.666152501887392e-20

R73_138 V73 V138 3070.232243785903
L73_138 V73 V138 3.9524492706212025e-12
C73_138 V73 V138 1.6145452756578144e-20

R73_139 V73 V139 -4120.407239511703
L73_139 V73 V139 -5.083925605332095e-12
C73_139 V73 V139 3.609653098872739e-20

R73_140 V73 V140 9530.176668162445
L73_140 V73 V140 2.2689587687234046e-11
C73_140 V73 V140 1.0775214458456887e-20

R73_141 V73 V141 16181.272299665532
L73_141 V73 V141 2.973940033475246e-11
C73_141 V73 V141 3.6243504453056183e-20

R73_142 V73 V142 6023.70063168231
L73_142 V73 V142 1.3562290944509625e-11
C73_142 V73 V142 -1.9024188949319073e-20

R73_143 V73 V143 9991.38364612063
L73_143 V73 V143 6.343611825646327e-12
C73_143 V73 V143 1.1416374166201262e-20

R73_144 V73 V144 -14235.296146889075
L73_144 V73 V144 -3.1481031698107316e-11
C73_144 V73 V144 -5.54549668025379e-20

R74_74 V74 0 -153.2817995021561
L74_74 V74 0 -1.3831885958561567e-13
C74_74 V74 0 -8.594764254598136e-19

R74_75 V74 V75 5279.991009393942
L74_75 V74 V75 2.7196106665232946e-12
C74_75 V74 V75 -3.4800825391772517e-20

R74_76 V74 V76 22227.705830692026
L74_76 V74 V76 3.5503418690968727e-12
C74_76 V74 V76 -5.885493259251898e-20

R74_77 V74 V77 -166211.43385146727
L74_77 V74 V77 9.0175971023236e-12
C74_77 V74 V77 -4.31628496101126e-20

R74_78 V74 V78 -52367.19799631725
L74_78 V74 V78 1.9720772567951763e-12
C74_78 V74 V78 1.8320794310421204e-19

R74_79 V74 V79 -4528.7947132015815
L74_79 V74 V79 -2.2986649717106794e-12
C74_79 V74 V79 -1.7562431789776546e-19

R74_80 V74 V80 11960.465712131061
L74_80 V74 V80 1.121264887340397e-11
C74_80 V74 V80 1.1618940267133303e-19

R74_81 V74 V81 37612.57566384333
L74_81 V74 V81 -6.0756916270447065e-12
C74_81 V74 V81 -2.3200458622403964e-20

R74_82 V74 V82 -7261.033155161901
L74_82 V74 V82 -1.7129160469852e-12
C74_82 V74 V82 -3.257409673515683e-19

R74_83 V74 V83 13760.33149591857
L74_83 V74 V83 -3.61158989461874e-12
C74_83 V74 V83 -1.551371143778289e-19

R74_84 V74 V84 -9236.948317440361
L74_84 V74 V84 -2.2295975543682648e-12
C74_84 V74 V84 -3.452488488687907e-20

R74_85 V74 V85 -10397.2759272297
L74_85 V74 V85 -4.404608647787235e-12
C74_85 V74 V85 3.529806363108072e-20

R74_86 V74 V86 -11499.972807839085
L74_86 V74 V86 4.708720461990298e-12
C74_86 V74 V86 1.7741462824080823e-19

R74_87 V74 V87 195667.64719033914
L74_87 V74 V87 4.914993101127463e-12
C74_87 V74 V87 7.01235591008883e-20

R74_88 V74 V88 30245.118682725664
L74_88 V74 V88 5.565901034666484e-12
C74_88 V74 V88 4.357326375583837e-20

R74_89 V74 V89 -38002.02823228657
L74_89 V74 V89 -1.855454661255694e-11
C74_89 V74 V89 -1.3251721291550527e-19

R74_90 V74 V90 9277.518920892353
L74_90 V74 V90 3.0702292322656252e-12
C74_90 V74 V90 9.395083957655371e-20

R74_91 V74 V91 -10324.968943633807
L74_91 V74 V91 -1.4931189166208718e-12
C74_91 V74 V91 -3.6964266906233217e-19

R74_92 V74 V92 -594965.649165164
L74_92 V74 V92 -1.1064963151389905e-11
C74_92 V74 V92 -2.759401367522693e-20

R74_93 V74 V93 -22475.47101241549
L74_93 V74 V93 -1.5178667918053225e-10
C74_93 V74 V93 -4.464168499407856e-21

R74_94 V74 V94 11279.938342421661
L74_94 V74 V94 4.049842407905773e-12
C74_94 V74 V94 1.9599417002641308e-19

R74_95 V74 V95 -71704.97501243066
L74_95 V74 V95 -3.224832661641369e-12
C74_95 V74 V95 -1.7215134600316918e-19

R74_96 V74 V96 21858.979902162668
L74_96 V74 V96 7.365360940116163e-12
C74_96 V74 V96 7.035873640078939e-20

R74_97 V74 V97 -21500.53733870741
L74_97 V74 V97 2.7804486611390984e-12
C74_97 V74 V97 1.301537889367323e-19

R74_98 V74 V98 -5171.975629095217
L74_98 V74 V98 -2.804645440694729e-11
C74_98 V74 V98 -4.891239415490942e-20

R74_99 V74 V99 -42770.43919626162
L74_99 V74 V99 -7.696392184771367e-12
C74_99 V74 V99 -2.1660956814475463e-20

R74_100 V74 V100 15575.723123734448
L74_100 V74 V100 1.4418666916325036e-11
C74_100 V74 V100 2.2695000671975686e-21

R74_101 V74 V101 -8435.661057279174
L74_101 V74 V101 -5.5838431913215025e-12
C74_101 V74 V101 -1.4092783688976707e-19

R74_102 V74 V102 11925.781430288796
L74_102 V74 V102 2.2312199878057602e-12
C74_102 V74 V102 1.7203156716235123e-19

R74_103 V74 V103 -6510.316612853315
L74_103 V74 V103 -2.768834606865102e-12
C74_103 V74 V103 -2.0723533181166561e-19

R74_104 V74 V104 10482.227048648732
L74_104 V74 V104 9.405780572855993e-12
C74_104 V74 V104 5.99496606871616e-20

R74_105 V74 V105 11336.9413205358
L74_105 V74 V105 5.3821888039156576e-12
C74_105 V74 V105 1.0240916418817743e-19

R74_106 V74 V106 9996.907777078675
L74_106 V74 V106 -2.6970257487090544e-12
C74_106 V74 V106 -2.0151181493061017e-19

R74_107 V74 V107 20071.101301797746
L74_107 V74 V107 2.612988913512784e-12
C74_107 V74 V107 2.1424235167981944e-19

R74_108 V74 V108 -10220.507564414691
L74_108 V74 V108 -3.49219451669114e-12
C74_108 V74 V108 -1.5736743224083056e-19

R74_109 V74 V109 -15782.245351357158
L74_109 V74 V109 -9.074571406204993e-12
C74_109 V74 V109 -2.76817036506061e-20

R74_110 V74 V110 10865.464843233327
L74_110 V74 V110 1.659466529313817e-12
C74_110 V74 V110 3.048011187879583e-19

R74_111 V74 V111 -12319.034807855382
L74_111 V74 V111 -8.457885503563203e-12
C74_111 V74 V111 -7.184707876506385e-20

R74_112 V74 V112 -15055.868564889468
L74_112 V74 V112 3.3251994929459206e-12
C74_112 V74 V112 1.1434305312474818e-19

R74_113 V74 V113 -12373.348349521288
L74_113 V74 V113 1.1388961880914906e-10
C74_113 V74 V113 -4.37904984887321e-20

R74_114 V74 V114 17708.052572931352
L74_114 V74 V114 -1.1110170186700752e-11
C74_114 V74 V114 -1.217701527929381e-19

R74_115 V74 V115 13316.591570022892
L74_115 V74 V115 4.700203631020648e-12
C74_115 V74 V115 1.236880134730451e-19

R74_116 V74 V116 -48829.04250101945
L74_116 V74 V116 -1.1843805871875752e-11
C74_116 V74 V116 -2.993323015184984e-20

R74_117 V74 V117 -25082.093511624473
L74_117 V74 V117 1.2588268367866682e-11
C74_117 V74 V117 4.2638883030535305e-20

R74_118 V74 V118 8887.475086283259
L74_118 V74 V118 4.673545123965055e-12
C74_118 V74 V118 1.641273329810499e-19

R74_119 V74 V119 -23822.410517889057
L74_119 V74 V119 7.227731187002962e-12
C74_119 V74 V119 1.1019134442508634e-19

R74_120 V74 V120 61968.53203588588
L74_120 V74 V120 7.082113903617961e-12
C74_120 V74 V120 -4.140962996332709e-20

R74_121 V74 V121 -5365.751908640232
L74_121 V74 V121 -2.4091545405652908e-11
C74_121 V74 V121 -4.303764984268095e-20

R74_122 V74 V122 -5450.329287220175
L74_122 V74 V122 3.0045546530150338e-12
C74_122 V74 V122 -3.098641273099779e-20

R74_123 V74 V123 31720.06773792627
L74_123 V74 V123 4.110701525045189e-12
C74_123 V74 V123 4.044817982682787e-20

R74_124 V74 V124 10668.583410552506
L74_124 V74 V124 1.784205105390161e-11
C74_124 V74 V124 -1.9003312392031405e-20

R74_125 V74 V125 4968.45843507949
L74_125 V74 V125 1.2095293899917356e-11
C74_125 V74 V125 3.3760726536291934e-20

R74_126 V74 V126 10634.833956132392
L74_126 V74 V126 -2.485887371892556e-12
C74_126 V74 V126 9.971547358133605e-21

R74_127 V74 V127 -14675.69578553429
L74_127 V74 V127 3.462879295517224e-12
C74_127 V74 V127 -5.6634831471189156e-21

R74_128 V74 V128 -7416.753447659573
L74_128 V74 V128 1.1289487654697713e-11
C74_128 V74 V128 7.169811668243886e-20

R74_129 V74 V129 14734.801002465822
L74_129 V74 V129 3.724861031943088e-12
C74_129 V74 V129 4.2246411242483524e-20

R74_130 V74 V130 -7132.399467103981
L74_130 V74 V130 -3.4776997674032846e-12
C74_130 V74 V130 -1.5894148918048858e-20

R74_131 V74 V131 -17081.198106126434
L74_131 V74 V131 -8.921568371396008e-12
C74_131 V74 V131 6.37142113833067e-20

R74_132 V74 V132 37923.235545965406
L74_132 V74 V132 -1.2392621837215494e-11
C74_132 V74 V132 1.4560753713016525e-20

R74_133 V74 V133 36334.251342840485
L74_133 V74 V133 -9.353339793328738e-12
C74_133 V74 V133 -4.4958632676867826e-20

R74_134 V74 V134 7696.3536756726435
L74_134 V74 V134 -6.285920934616383e-11
C74_134 V74 V134 3.569186859490676e-20

R74_135 V74 V135 -25481.72852139356
L74_135 V74 V135 5.255113199092344e-12
C74_135 V74 V135 -4.241249179369793e-20

R74_136 V74 V136 -18502.749885145993
L74_136 V74 V136 -9.766237742512847e-12
C74_136 V74 V136 -5.973567542840439e-20

R74_137 V74 V137 8438.656457108455
L74_137 V74 V137 -3.778560543872226e-11
C74_137 V74 V137 -3.071040147073269e-20

R74_138 V74 V138 -80613.13221401429
L74_138 V74 V138 -2.017889253697498e-12
C74_138 V74 V138 -3.367037411255956e-20

R74_139 V74 V139 -8625.844860805018
L74_139 V74 V139 2.526012326199096e-12
C74_139 V74 V139 2.0686118938582693e-20

R74_140 V74 V140 22112.538272420727
L74_140 V74 V140 -4.232711877555549e-12
C74_140 V74 V140 -5.887571795128966e-20

R74_141 V74 V141 10671.71766431524
L74_141 V74 V141 -1.6126908246565162e-11
C74_141 V74 V141 -1.3847989519932786e-20

R74_142 V74 V142 108582.1455691046
L74_142 V74 V142 -4.871113261837982e-12
C74_142 V74 V142 -3.854296447650672e-21

R74_143 V74 V143 -22551.432490315467
L74_143 V74 V143 -1.270402317884734e-11
C74_143 V74 V143 5.2571028620203965e-20

R74_144 V74 V144 4817228.152606465
L74_144 V74 V144 6.188498151148797e-12
C74_144 V74 V144 1.5797455672242725e-20

R75_75 V75 0 129.69073593046815
L75_75 V75 0 1.6098149181818187e-13
C75_75 V75 0 7.910449075010147e-19

R75_76 V75 V76 -22253.255349666702
L75_76 V75 V76 -3.920891105025347e-11
C75_76 V75 V76 2.4772956633431192e-19

R75_77 V75 V77 -27548.198489842496
L75_77 V75 V77 -3.945090751702436e-12
C75_77 V75 V77 -5.894586681410689e-20

R75_78 V75 V78 6836.153737266667
L75_78 V75 V78 2.2880629272603913e-12
C75_78 V75 V78 3.331538818839655e-19

R75_79 V75 V79 4384.054742246432
L75_79 V75 V79 1.596058993358735e-12
C75_79 V75 V79 3.7484510888414707e-19

R75_80 V75 V80 -10930.27450978483
L75_80 V75 V80 -3.2614046161253247e-12
C75_80 V75 V80 -3.2316854922414184e-19

R75_81 V75 V81 21435.31428600105
L75_81 V75 V81 2.578823108106239e-12
C75_81 V75 V81 1.7332210070185972e-19

R75_82 V75 V82 -7436.905718837035
L75_82 V75 V82 -1.0273147684893035e-12
C75_82 V75 V82 -5.394988013580604e-19

R75_83 V75 V83 -3651.20661793598
L75_83 V75 V83 -1.1870046730266976e-12
C75_83 V75 V83 -5.799184461500151e-19

R75_84 V75 V84 22656.148028852156
L75_84 V75 V84 4.842832612814769e-12
C75_84 V75 V84 1.1786239336338968e-20

R75_85 V75 V85 5528.1972018518545
L75_85 V75 V85 1.4505678229902394e-12
C75_85 V75 V85 3.464735663935669e-19

R75_86 V75 V86 8127.630488965314
L75_86 V75 V86 2.547257675106567e-12
C75_86 V75 V86 1.7164336064790327e-19

R75_87 V75 V87 8922.326304717259
L75_87 V75 V87 1.9039283231207355e-12
C75_87 V75 V87 3.13511024478726e-19

R75_88 V75 V88 24822.0503479395
L75_88 V75 V88 1.1974303019363294e-11
C75_88 V75 V88 1.1126607017701143e-19

R75_89 V75 V89 -298209.5076693391
L75_89 V75 V89 -5.127146577567753e-12
C75_89 V75 V89 -8.892020097747423e-20

R75_90 V75 V90 -5503.35947039935
L75_90 V75 V90 -1.7442849493729635e-12
C75_90 V75 V90 -3.4668683248347292e-19

R75_91 V75 V91 -6583.931579092527
L75_91 V75 V91 -1.1907856577496253e-12
C75_91 V75 V91 -4.823832599388357e-19

R75_92 V75 V92 -7884.687115960344
L75_92 V75 V92 -1.7558434613560505e-12
C75_92 V75 V92 -3.6369422146289985e-19

R75_93 V75 V93 5636.237953627117
L75_93 V75 V93 4.874298185833016e-12
C75_93 V75 V93 1.440581402292641e-19

R75_94 V75 V94 9294.285803156117
L75_94 V75 V94 3.6032328496456305e-12
C75_94 V75 V94 1.2269981862381685e-19

R75_95 V75 V95 -7489.902317280193
L75_95 V75 V95 -2.0394417666050513e-12
C75_95 V75 V95 -2.8446714559330105e-19

R75_96 V75 V96 -6351.596314899133
L75_96 V75 V96 -2.350983597688082e-12
C75_96 V75 V96 -2.9015682268593725e-19

R75_97 V75 V97 10481.559171877201
L75_97 V75 V97 1.0155328756766082e-11
C75_97 V75 V97 3.1690345304001685e-20

R75_98 V75 V98 59066.54056018511
L75_98 V75 V98 -2.41798725291299e-12
C75_98 V75 V98 -3.0347590819306396e-19

R75_99 V75 V99 6184.311858358554
L75_99 V75 V99 3.975362256668222e-12
C75_99 V75 V99 7.318499614673508e-20

R75_100 V75 V100 70530.73692457062
L75_100 V75 V100 9.264819417819e-12
C75_100 V75 V100 6.330537538690147e-20

R75_101 V75 V101 29745.02769637434
L75_101 V75 V101 -3.1352872491909536e-12
C75_101 V75 V101 -2.095884235662616e-19

R75_102 V75 V102 -3770.850109181348
L75_102 V75 V102 -7.922640469818773e-13
C75_102 V75 V102 -8.223121064132966e-19

R75_103 V75 V103 3822.722450391086
L75_103 V75 V103 1.515468535229585e-12
C75_103 V75 V103 4.682472124460867e-19

R75_104 V75 V104 -49390.960982111086
L75_104 V75 V104 -5.0934167249623036e-12
C75_104 V75 V104 -1.8276993928132823e-19

R75_105 V75 V105 10330.299183677333
L75_105 V75 V105 1.0946926754380335e-12
C75_105 V75 V105 5.857846069607496e-19

R75_106 V75 V106 -2491.661642561667
L75_106 V75 V106 -6.780525521587272e-13
C75_106 V75 V106 -9.235917855750765e-19

R75_107 V75 V107 -4318.543875176572
L75_107 V75 V107 -9.988105069557993e-13
C75_107 V75 V107 -7.119054191061209e-19

R75_108 V75 V108 5825.382629448563
L75_108 V75 V108 1.259538904704532e-12
C75_108 V75 V108 5.094122691755438e-19

R75_109 V75 V109 8624.232862364715
L75_109 V75 V109 4.380165846897113e-12
C75_109 V75 V109 9.048094641999274e-20

R75_110 V75 V110 13637.716814455247
L75_110 V75 V110 1.0762921625301686e-12
C75_110 V75 V110 7.077578975498457e-19

R75_111 V75 V111 3467.093917562383
L75_111 V75 V111 1.2915568497929764e-12
C75_111 V75 V111 4.0306999705596677e-19

R75_112 V75 V112 -5151.925398258753
L75_112 V75 V112 -1.5137138071336583e-12
C75_112 V75 V112 -4.396797377509693e-19

R75_113 V75 V113 -5370.788266187093
L75_113 V75 V113 -2.5046750315927867e-12
C75_113 V75 V113 -2.184484601038077e-19

R75_114 V75 V114 -11913.448957118691
L75_114 V75 V114 -1.886681956206675e-12
C75_114 V75 V114 -3.5884194435504133e-19

R75_115 V75 V115 -5290.653571799255
L75_115 V75 V115 -1.695873300237058e-12
C75_115 V75 V115 -3.878156165929154e-19

R75_116 V75 V116 5486.545669447048
L75_116 V75 V116 1.801181183837697e-12
C75_116 V75 V116 3.153096822147493e-19

R75_117 V75 V117 11894.785785786262
L75_117 V75 V117 2.873385424605741e-12
C75_117 V75 V117 2.9369282329265696e-19

R75_118 V75 V118 16011.85074425876
L75_118 V75 V118 1.901896240077837e-12
C75_118 V75 V118 3.3432854386315413e-19

R75_119 V75 V119 5722.350681601923
L75_119 V75 V119 1.328757492498171e-12
C75_119 V75 V119 4.2122269623489013e-19

R75_120 V75 V120 -3235.434755077816
L75_120 V75 V120 -2.4128286394695626e-12
C75_120 V75 V120 1.1759079616383686e-19

R75_121 V75 V121 26197.299070609635
L75_121 V75 V121 -1.4098371150704839e-11
C75_121 V75 V121 -1.3999045004133576e-19

R75_122 V75 V122 -2598.058255064964
L75_122 V75 V122 -2.5053442901897037e-12
C75_122 V75 V122 -8.985864772373509e-21

R75_123 V75 V123 27865.42629624766
L75_123 V75 V123 1.1710056741018702e-11
C75_123 V75 V123 8.047707732452417e-20

R75_124 V75 V124 6165.251239879273
L75_124 V75 V124 3.5415357425141587e-12
C75_124 V75 V124 1.1812566549112113e-19

R75_125 V75 V125 -8615.817177180905
L75_125 V75 V125 -4.582604169247924e-12
C75_125 V75 V125 6.051319498449742e-20

R75_126 V75 V126 1733.7643936424251
L75_126 V75 V126 1.7421451169993987e-12
C75_126 V75 V126 -1.132728457508615e-19

R75_127 V75 V127 -2159.990421894232
L75_127 V75 V127 -1.5565664292572519e-12
C75_127 V75 V127 1.5356365586153235e-21

R75_128 V75 V128 -25343.744173060495
L75_128 V75 V128 2.3555042270599948e-11
C75_128 V75 V128 1.0338427966936913e-19

R75_129 V75 V129 -18657.396752769335
L75_129 V75 V129 -2.8342986003437463e-11
C75_129 V75 V129 8.11538025746507e-20

R75_130 V75 V130 8482.337874964698
L75_130 V75 V130 2.461645974157343e-12
C75_130 V75 V130 2.3346671017880596e-19

R75_131 V75 V131 428602.10026841244
L75_131 V75 V131 -4.887918827700585e-12
C75_131 V75 V131 -2.1311793650432838e-19

R75_132 V75 V132 9278.49361520241
L75_132 V75 V132 3.91660715203522e-12
C75_132 V75 V132 8.813313722064429e-20

R75_133 V75 V133 -7331.450559881789
L75_133 V75 V133 -2.1473214777103177e-12
C75_133 V75 V133 -2.6628617548446833e-19

R75_134 V75 V134 -38270.48327192907
L75_134 V75 V134 -3.2704901349415165e-11
C75_134 V75 V134 -1.024367954971495e-20

R75_135 V75 V135 -3417.092119443385
L75_135 V75 V135 -2.7590004050748703e-12
C75_135 V75 V135 5.404700481042496e-20

R75_136 V75 V136 -30426.30468625021
L75_136 V75 V136 -4.960404613981973e-12
C75_136 V75 V136 -1.0579944242952803e-19

R75_137 V75 V137 30497.027923671256
L75_137 V75 V137 6.146161027233385e-11
C75_137 V75 V137 9.908152127120699e-20

R75_138 V75 V138 2356.233624212824
L75_138 V75 V138 1.8111261070570875e-12
C75_138 V75 V138 6.335001727587254e-20

R75_139 V75 V139 -1640.9692880454966
L75_139 V75 V139 -1.0902887623216623e-12
C75_139 V75 V139 -1.0757755505663293e-19

R75_140 V75 V140 32801.54975823699
L75_140 V75 V140 5.520916912336889e-12
C75_140 V75 V140 3.70319645880116e-21

R75_141 V75 V141 5238.476607310911
L75_141 V75 V141 6.615264840058784e-12
C75_141 V75 V141 -6.946516048405707e-21

R75_142 V75 V142 29205.284082857546
L75_142 V75 V142 2.8882640915854733e-12
C75_142 V75 V142 1.2221032276554245e-19

R75_143 V75 V143 5369.155658017143
L75_143 V75 V143 3.497643285082201e-12
C75_143 V75 V143 2.7901671313250184e-20

R75_144 V75 V144 -10010.375556533601
L75_144 V75 V144 -6.792130243422067e-12
C75_144 V75 V144 -9.723269176816881e-21

R76_76 V76 0 139.36326060134965
L76_76 V76 0 7.790526901698648e-14
C76_76 V76 0 1.1293521954967006e-18

R76_77 V76 V77 -13711.250159397394
L76_77 V76 V77 -4.875663944732585e-12
C76_77 V76 V77 3.2610728168863854e-22

R76_78 V76 V78 -9492.825960849947
L76_78 V76 V78 -1.973017030738464e-12
C76_78 V76 V78 -2.4014195398684425e-19

R76_79 V76 V79 -5267.171758351939
L76_79 V76 V79 -1.727868310488952e-12
C76_79 V76 V79 -4.965162150068458e-19

R76_80 V76 V80 2836.1972895864965
L76_80 V76 V80 8.987283684053434e-13
C76_80 V76 V80 7.159874190084183e-19

R76_81 V76 V81 -20694.26554248547
L76_81 V76 V81 -3.000419106129829e-12
C76_81 V76 V81 -2.82341557954862e-19

R76_82 V76 V82 5786.918871984327
L76_82 V76 V82 1.7488521723072157e-12
C76_82 V76 V82 4.794327142721756e-19

R76_83 V76 V83 4703.50642939796
L76_83 V76 V83 1.1618788935898017e-12
C76_83 V76 V83 4.637647673799186e-19

R76_84 V76 V84 -4783.695907453084
L76_84 V76 V84 -3.704829219116397e-12
C76_84 V76 V84 -2.3854115381687035e-19

R76_85 V76 V85 -5009.449154397187
L76_85 V76 V85 -1.507135441886595e-12
C76_85 V76 V85 -5.035551959290309e-19

R76_86 V76 V86 -9995.160664889796
L76_86 V76 V86 -4.134270220705578e-12
C76_86 V76 V86 -1.6212071847081135e-19

R76_87 V76 V87 -4778.553450399863
L76_87 V76 V87 -1.1586543768762977e-12
C76_87 V76 V87 -5.435513617736386e-19

R76_88 V76 V88 -171910.12315021563
L76_88 V76 V88 -4.286584945136479e-12
C76_88 V76 V88 -1.1659576915076157e-19

R76_89 V76 V89 5706.854892286196
L76_89 V76 V89 2.163521003775056e-12
C76_89 V76 V89 3.734521308547483e-19

R76_90 V76 V90 3516.893256755167
L76_90 V76 V90 1.1837823767836698e-12
C76_90 V76 V90 4.707182009319335e-19

R76_91 V76 V91 6972.517058886026
L76_91 V76 V91 1.824321182888428e-12
C76_91 V76 V91 2.911433303688875e-19

R76_92 V76 V92 5735.6909984420445
L76_92 V76 V92 1.3553144511655342e-12
C76_92 V76 V92 5.000657174377954e-19

R76_93 V76 V93 8596.373750462719
L76_93 V76 V93 -3.8651597775419134e-12
C76_93 V76 V93 -5.166472505401666e-20

R76_94 V76 V94 -25609.005364638862
L76_94 V76 V94 -3.2769696831309085e-12
C76_94 V76 V94 -5.75538295242672e-20

R76_95 V76 V95 12015.066960486669
L76_95 V76 V95 3.2235595335914244e-12
C76_95 V76 V95 2.275467843215118e-19

R76_96 V76 V96 10468.954561282299
L76_96 V76 V96 1.4699885921567299e-12
C76_96 V76 V96 4.638312107104829e-19

R76_97 V76 V97 4609.7352639791725
L76_97 V76 V97 2.386766204196154e-12
C76_97 V76 V97 1.1419973334316387e-19

R76_98 V76 V98 2898.106771302654
L76_98 V76 V98 9.815325637148137e-13
C76_98 V76 V98 4.443983825200535e-19

R76_99 V76 V99 -14349.173030213438
L76_99 V76 V99 -2.385586118191006e-12
C76_99 V76 V99 -1.1912706264819794e-19

R76_100 V76 V100 -30291.953051808767
L76_100 V76 V100 -4.7057237964556846e-12
C76_100 V76 V100 -1.4194650400655546e-19

R76_101 V76 V101 3830.075639791621
L76_101 V76 V101 1.2608871024731226e-12
C76_101 V76 V101 5.291783876793899e-19

R76_102 V76 V102 1595.4229862031875
L76_102 V76 V102 4.89550829600408e-13
C76_102 V76 V102 1.2068159543021586e-18

R76_103 V76 V103 -5676.320016450721
L76_103 V76 V103 -1.051536671807325e-12
C76_103 V76 V103 -6.689924187828037e-19

R76_104 V76 V104 19689.294025928855
L76_104 V76 V104 4.433103255137651e-12
C76_104 V76 V104 2.7208747475785655e-19

R76_105 V76 V105 -3335.949965395316
L76_105 V76 V105 -9.12062493136061e-13
C76_105 V76 V105 -5.978661073799779e-19

R76_106 V76 V106 3787.567159898758
L76_106 V76 V106 6.94893707988393e-13
C76_106 V76 V106 1.0325087019464471e-18

R76_107 V76 V107 2570.800767122386
L76_107 V76 V107 6.326326869262486e-13
C76_107 V76 V107 9.57103499158693e-19

R76_108 V76 V108 -2540.1455510078276
L76_108 V76 V108 -6.470324880310264e-13
C76_108 V76 V108 -1.0666877544270016e-18

R76_109 V76 V109 -11201.38026402779
L76_109 V76 V109 -2.699552965847137e-12
C76_109 V76 V109 -2.1176303221537486e-19

R76_110 V76 V110 -4911.914894921631
L76_110 V76 V110 -1.062683297723279e-12
C76_110 V76 V110 -7.107644918212356e-19

R76_111 V76 V111 -4312.883405853723
L76_111 V76 V111 -1.139857928674069e-12
C76_111 V76 V111 -5.398721171061462e-19

R76_112 V76 V112 2183.1887501631813
L76_112 V76 V112 5.613187761579417e-13
C76_112 V76 V112 8.760652250457769e-19

R76_113 V76 V113 8037.819079731039
L76_113 V76 V113 1.3642539137039073e-12
C76_113 V76 V113 3.143524076552551e-19

R76_114 V76 V114 3820.348698419896
L76_114 V76 V114 1.27653524622653e-12
C76_114 V76 V114 4.425994379076518e-19

R76_115 V76 V115 3649.2245063841333
L76_115 V76 V115 1.2836085933324101e-12
C76_115 V76 V115 5.034233606035986e-19

R76_116 V76 V116 -3605.321034659774
L76_116 V76 V116 -1.0055768599758307e-12
C76_116 V76 V116 -5.552907677729462e-19

R76_117 V76 V117 -10513.095604914986
L76_117 V76 V117 -1.8030721344511146e-12
C76_117 V76 V117 -4.448125539850862e-19

R76_118 V76 V118 -4559.185863889529
L76_118 V76 V118 -1.3527359581888954e-12
C76_118 V76 V118 -3.4140406984385255e-19

R76_119 V76 V119 -3223.620588100219
L76_119 V76 V119 -1.2056242659189965e-12
C76_119 V76 V119 -5.079895745246291e-19

R76_120 V76 V120 6231.766575985359
L76_120 V76 V120 4.575864941771609e-12
C76_120 V76 V120 -2.2774916730537625e-19

R76_121 V76 V121 10973.021502954627
L76_121 V76 V121 1.780749706103688e-12
C76_121 V76 V121 7.158467061203958e-20

R76_122 V76 V122 2716.9518486862266
L76_122 V76 V122 7.823707256006659e-13
C76_122 V76 V122 8.490421177288167e-21

R76_123 V76 V123 6643.832699356797
L76_123 V76 V123 4.382310812021011e-12
C76_123 V76 V123 -3.008372014172277e-20

R76_124 V76 V124 36384.48662824123
L76_124 V76 V124 -6.075599859928032e-12
C76_124 V76 V124 -1.4223841710158916e-19

R76_125 V76 V125 72628.30404908914
L76_125 V76 V125 -2.1349752805331706e-12
C76_125 V76 V125 -1.1152545521436697e-19

R76_126 V76 V126 -2795.8175741849645
L76_126 V76 V126 -8.369818695046544e-13
C76_126 V76 V126 1.1567687503520442e-19

R76_127 V76 V127 3054.003596713552
L76_127 V76 V127 1.0308739870083321e-12
C76_127 V76 V127 -1.4455290842836867e-20

R76_128 V76 V128 54799.44525184469
L76_128 V76 V128 2.2737551145368823e-11
C76_128 V76 V128 -3.292374938625581e-20

R76_129 V76 V129 4692.085027858509
L76_129 V76 V129 3.393654302695333e-12
C76_129 V76 V129 -6.433807624051677e-20

R76_130 V76 V130 -3241.118490319256
L76_130 V76 V130 -1.1998550447895098e-12
C76_130 V76 V130 -3.4991615790768317e-19

R76_131 V76 V131 -10981.177564170204
L76_131 V76 V131 2.4904686269517154e-11
C76_131 V76 V131 2.5997194198792896e-19

R76_132 V76 V132 -7833.301709519967
L76_132 V76 V132 -2.6991082905859774e-12
C76_132 V76 V132 -5.607735873952418e-20

R76_133 V76 V133 48189.54173352096
L76_133 V76 V133 3.360586122971188e-12
C76_133 V76 V133 2.8911639770013537e-19

R76_134 V76 V134 -8164.538230261047
L76_134 V76 V134 -4.017756667177135e-12
C76_134 V76 V134 2.6750044390187835e-20

R76_135 V76 V135 5915.762945141542
L76_135 V76 V135 1.788954082076327e-12
C76_135 V76 V135 -1.186704851762295e-19

R76_136 V76 V136 -54734.53993404378
L76_136 V76 V136 3.16333906639543e-11
C76_136 V76 V136 1.8042100617109146e-20

R76_137 V76 V137 67186.50075867324
L76_137 V76 V137 -2.1495760771600925e-12
C76_137 V76 V137 -1.981465141937069e-19

R76_138 V76 V138 -2186.3192705780243
L76_138 V76 V138 -7.809225048034391e-13
C76_138 V76 V138 -9.005621429175762e-20

R76_139 V76 V139 2054.286227771546
L76_139 V76 V139 6.89870351703907e-13
C76_139 V76 V139 1.7574733370930495e-19

R76_140 V76 V140 -3794.6484352762536
L76_140 V76 V140 -1.4881752011901316e-12
C76_140 V76 V140 -9.333893868643403e-20

R76_141 V76 V141 -69872.88537641145
L76_141 V76 V141 -3.259032386387793e-12
C76_141 V76 V141 -3.3897427837904406e-20

R76_142 V76 V142 -3099.478695642132
L76_142 V76 V142 -1.6826307530283249e-12
C76_142 V76 V142 -1.1924475398218595e-19

R76_143 V76 V143 -5821.160594822836
L76_143 V76 V143 -2.929605652212735e-12
C76_143 V76 V143 1.6337062805436887e-20

R76_144 V76 V144 14713.45495686565
L76_144 V76 V144 2.4723501442383822e-12
C76_144 V76 V144 2.2248083009444704e-20

R77_77 V77 0 541.2894726065747
L77_77 V77 0 4.823725576255749e-13
C77_77 V77 0 7.03316705914713e-20

R77_78 V77 V78 303505.73419948743
L77_78 V77 V78 3.1666094439007046e-11
C77_78 V77 V78 5.605447593099094e-20

R77_79 V77 V79 -18630.869671791377
L77_79 V77 V79 -1.4807057429240915e-11
C77_79 V77 V79 -7.981767628694453e-20

R77_80 V77 V80 -26421.522212382777
L77_80 V77 V80 -5.46163198386255e-12
C77_80 V77 V80 -1.1972484414146643e-19

R77_81 V77 V81 5074.10779432302
L77_81 V77 V81 9.417964691839169e-13
C77_81 V77 V81 6.074703714984018e-19

R77_82 V77 V82 -71860.98253505064
L77_82 V77 V82 -7.085879331279903e-12
C77_82 V77 V82 1.3274019562763545e-20

R77_83 V77 V83 -57179.87780056095
L77_83 V77 V83 -3.7864407056688684e-12
C77_83 V77 V83 -1.761187100534662e-19

R77_84 V77 V84 -9318.976264717914
L77_84 V77 V84 -9.119639223773707e-12
C77_84 V77 V84 -1.1853016759706886e-19

R77_85 V77 V85 -56036.81856345449
L77_85 V77 V85 4.529003970300566e-12
C77_85 V77 V85 5.968841004341769e-20

R77_86 V77 V86 -32251.19794969344
L77_86 V77 V86 5.29128799713534e-12
C77_86 V77 V86 3.123645012593901e-20

R77_87 V77 V87 -776854.0608357509
L77_87 V77 V87 2.445120921551802e-11
C77_87 V77 V87 1.0995822626195209e-20

R77_88 V77 V88 33843.566675174734
L77_88 V77 V88 5.244609103213331e-12
C77_88 V77 V88 1.348958899941331e-19

R77_89 V77 V89 -62134.552426391034
L77_89 V77 V89 -5.012587253526052e-12
C77_89 V77 V89 -3.028388495252702e-20

R77_90 V77 V90 9205.926931134187
L77_90 V77 V90 4.148513979909686e-12
C77_90 V77 V90 1.0786116340959691e-19

R77_91 V77 V91 20289.409888712813
L77_91 V77 V91 1.1569407049605676e-11
C77_91 V77 V91 7.229409583394925e-20

R77_92 V77 V92 -7101.636827687016
L77_92 V77 V92 -1.5769280133933039e-12
C77_92 V77 V92 -3.898121246931411e-19

R77_93 V77 V93 -43848.17186278245
L77_93 V77 V93 2.5407397942914127e-11
C77_93 V77 V93 4.087455479888582e-20

R77_94 V77 V94 63590.27641932502
L77_94 V77 V94 2.7046086828349814e-12
C77_94 V77 V94 2.459054784967727e-19

R77_95 V77 V95 -200337.909931593
L77_95 V77 V95 -6.09012316039565e-11
C77_95 V77 V95 8.504713400828266e-21

R77_96 V77 V96 -5078.842500658037
L77_96 V77 V96 -1.1759314606415536e-12
C77_96 V77 V96 -5.158074395534924e-19

R77_97 V77 V97 5710.903606824074
L77_97 V77 V97 2.3198179284877765e-12
C77_97 V77 V97 2.0772731810368785e-19

R77_98 V77 V98 7651.553202488859
L77_98 V77 V98 -5.537082731168816e-12
C77_98 V77 V98 -9.759590984247022e-20

R77_99 V77 V99 -26315.194504841493
L77_99 V77 V99 -3.378278526176009e-11
C77_99 V77 V99 4.3811397860732545e-20

R77_100 V77 V100 17578.54192478508
L77_100 V77 V100 2.6191161986551256e-12
C77_100 V77 V100 2.580199387008911e-19

R77_101 V77 V101 -47239.47362330314
L77_101 V77 V101 -2.7552437794234526e-12
C77_101 V77 V101 -1.4339204836942775e-19

R77_102 V77 V102 5943.9721891401205
L77_102 V77 V102 2.5177456452453325e-12
C77_102 V77 V102 2.4299139396138143e-19

R77_103 V77 V103 -35389.26125926601
L77_103 V77 V103 -6.581403451444736e-12
C77_103 V77 V103 -7.8779450097494e-20

R77_104 V77 V104 -5912.944200625271
L77_104 V77 V104 -1.4183746402515802e-12
C77_104 V77 V104 -4.741943064534841e-19

R77_105 V77 V105 -260470.77682174538
L77_105 V77 V105 3.604480047757631e-12
C77_105 V77 V105 2.3423189306537836e-19

R77_106 V77 V106 -9004.026960021047
L77_106 V77 V106 -4.4553518391180265e-12
C77_106 V77 V106 -1.2756222292574933e-19

R77_107 V77 V107 10362.14184020732
L77_107 V77 V107 2.993693527727594e-12
C77_107 V77 V107 1.8840955189251366e-19

R77_108 V77 V108 13686.548195975567
L77_108 V77 V108 1.3805682412994008e-11
C77_108 V77 V108 4.847312010976448e-20

R77_109 V77 V109 -9692.516985498967
L77_109 V77 V109 -1.550882892796091e-12
C77_109 V77 V109 -4.778893357350323e-19

R77_110 V77 V110 11589.058391718563
L77_110 V77 V110 3.39413999222355e-12
C77_110 V77 V110 9.774172053843149e-20

R77_111 V77 V111 -113907.39075613768
L77_111 V77 V111 -1.010480548400577e-11
C77_111 V77 V111 -6.781008481167734e-21

R77_112 V77 V112 5085.516406762806
L77_112 V77 V112 1.0353709244121149e-11
C77_112 V77 V112 4.854551505231847e-20

R77_113 V77 V113 6628.982991369081
L77_113 V77 V113 7.2292504828815045e-12
C77_113 V77 V113 1.1230603487280532e-19

R77_114 V77 V114 1430392.7707075293
L77_114 V77 V114 9.201612078173734e-11
C77_114 V77 V114 -1.3336701336159315e-20

R77_115 V77 V115 14582.27007775176
L77_115 V77 V115 5.287288354372292e-12
C77_115 V77 V115 8.738102038021694e-20

R77_116 V77 V116 -50397.27586331597
L77_116 V77 V116 3.9389794650158064e-11
C77_116 V77 V116 2.1989813328986715e-20

R77_117 V77 V117 -64238.16575887786
L77_117 V77 V117 -5.588257585278612e-11
C77_117 V77 V117 -7.98663354221298e-20

R77_118 V77 V118 -8338.229815819388
L77_118 V77 V118 -8.907287586725588e-12
C77_118 V77 V118 -6.017566899620535e-20

R77_119 V77 V119 19285.520338325958
L77_119 V77 V119 1.657937004122315e-11
C77_119 V77 V119 7.16512594476541e-20

R77_120 V77 V120 5348.40468255963
L77_120 V77 V120 2.8692107858140125e-12
C77_120 V77 V120 4.10354679785293e-20

R77_121 V77 V121 4867.628638661856
L77_121 V77 V121 8.168176510639581e-11
C77_121 V77 V121 -1.2308654733995332e-20

R77_122 V77 V122 2016.448967384607
L77_122 V77 V122 3.207292512512511e-12
C77_122 V77 V122 -4.208454587080888e-20

R77_123 V77 V123 11983.917449500655
L77_123 V77 V123 1.788977462917674e-11
C77_123 V77 V123 -5.2479539697476944e-20

R77_124 V77 V124 65333.19153391431
L77_124 V77 V124 2.0750860511376575e-11
C77_124 V77 V124 6.870229246433657e-20

R77_125 V77 V125 -7126.769867053217
L77_125 V77 V125 9.29433331485008e-12
C77_125 V77 V125 -3.603193855963354e-21

R77_126 V77 V126 -2116.144894902997
L77_126 V77 V126 -1.9456947277393264e-12
C77_126 V77 V126 2.5369915540900108e-21

R77_127 V77 V127 2884.1499332886333
L77_127 V77 V127 2.7214052958855236e-12
C77_127 V77 V127 1.236754113886772e-20

R77_128 V77 V128 14624.048282280874
L77_128 V77 V128 8.299888225203781e-12
C77_128 V77 V128 6.760304466687367e-20

R77_129 V77 V129 7855.593783999966
L77_129 V77 V129 4.934081019346569e-12
C77_129 V77 V129 1.987990873638198e-20

R77_130 V77 V130 -14652.730970445753
L77_130 V77 V130 -7.492790134817974e-12
C77_130 V77 V130 3.6754306164420584e-20

R77_131 V77 V131 -10482.175006545307
L77_131 V77 V131 -1.583563126389887e-11
C77_131 V77 V131 6.045940981891271e-20

R77_132 V77 V132 -19194.200991154074
L77_132 V77 V132 8.096805500684299e-12
C77_132 V77 V132 1.3224444387271773e-19

R77_133 V77 V133 -11350.065467066299
L77_133 V77 V133 -6.537692104162369e-12
C77_133 V77 V133 -8.410869154649268e-20

R77_134 V77 V134 -8000.264407541313
L77_134 V77 V134 -1.4320659152293843e-11
C77_134 V77 V134 4.925130489873466e-21

R77_135 V77 V135 4420.577199628787
L77_135 V77 V135 4.0476435090761455e-12
C77_135 V77 V135 -7.372116395288672e-21

R77_136 V77 V136 95228.95855240371
L77_136 V77 V136 -5.685374283427814e-12
C77_136 V77 V136 -1.1852523292959357e-19

R77_137 V77 V137 -13545.000960699697
L77_137 V77 V137 1.5472745258689538e-11
C77_137 V77 V137 5.1762380386275995e-20

R77_138 V77 V138 -2358.8263647451868
L77_138 V77 V138 -1.737269320775072e-12
C77_138 V77 V138 -6.251546931681731e-20

R77_139 V77 V139 2280.73771762101
L77_139 V77 V139 2.232077145724786e-12
C77_139 V77 V139 -3.105824668757701e-20

R77_140 V77 V140 -6463.874742165929
L77_140 V77 V140 -6.082555204370345e-12
C77_140 V77 V140 -3.7868274841321955e-20

R77_141 V77 V141 -7330.319769560031
L77_141 V77 V141 -6.058162535738422e-12
C77_141 V77 V141 -5.667125236089786e-20

R77_142 V77 V142 -8739.418056361057
L77_142 V77 V142 -4.394573357950582e-12
C77_142 V77 V142 -7.233768724648238e-21

R77_143 V77 V143 -9085.958893092182
L77_143 V77 V143 -4.828729525644567e-12
C77_143 V77 V143 -4.5672215929934904e-21

R77_144 V77 V144 11759.098923672318
L77_144 V77 V144 1.2518652796712158e-11
C77_144 V77 V144 4.638990929506878e-20

R78_78 V78 0 4046.493832438698
L78_78 V78 0 1.7785317214142426e-13
C78_78 V78 0 1.0422458860643176e-18

R78_79 V78 V79 -10062.182168968859
L78_79 V78 V79 -1.8156706423367824e-11
C78_79 V78 V79 -7.948689267855017e-20

R78_80 V78 V80 9246.503991972777
L78_80 V78 V80 4.270901091098787e-12
C78_80 V78 V80 1.6968350964856562e-19

R78_81 V78 V81 -28093.9498555908
L78_81 V78 V81 -7.269626017274518e-12
C78_81 V78 V81 -1.3895285500664108e-19

R78_82 V78 V82 3328.0679300155857
L78_82 V78 V82 6.817463939371311e-13
C78_82 V78 V82 1.027028106061704e-18

R78_83 V78 V83 3475.1006659792924
L78_83 V78 V83 8.232115013997891e-13
C78_83 V78 V83 7.372119825764136e-19

R78_84 V78 V84 -12396.191031431026
L78_84 V78 V84 -2.3042037194346067e-11
C78_84 V78 V84 -2.615578022777724e-20

R78_85 V78 V85 -6192.847057835891
L78_85 V78 V85 -1.7324717211300201e-12
C78_85 V78 V85 -4.050238967671937e-19

R78_86 V78 V86 -6552.988832444134
L78_86 V78 V86 -2.2530287635994663e-12
C78_86 V78 V86 -2.745590609188307e-19

R78_87 V78 V87 -6415.940433927193
L78_87 V78 V87 -1.6797424559028579e-12
C78_87 V78 V87 -4.189097803899839e-19

R78_88 V78 V88 -22701.319194185086
L78_88 V78 V88 -3.791061867574618e-12
C78_88 V78 V88 -1.750366743216737e-19

R78_89 V78 V89 7555.7880535306695
L78_89 V78 V89 2.5226296827502893e-12
C78_89 V78 V89 3.2939376491926516e-19

R78_90 V78 V90 9723.697648846026
L78_90 V78 V90 3.569238857120129e-12
C78_90 V78 V90 1.4609847239191043e-19

R78_91 V78 V91 3691.041630106056
L78_91 V78 V91 8.675824711768682e-13
C78_91 V78 V91 7.3128937245856865e-19

R78_92 V78 V92 7096.797539749281
L78_92 V78 V92 1.7791043969762846e-12
C78_92 V78 V92 3.886334995989474e-19

R78_93 V78 V93 -22617.09239859873
L78_93 V78 V93 -6.616343392771939e-12
C78_93 V78 V93 -5.444436963122367e-20

R78_94 V78 V94 -7164.274128759226
L78_94 V78 V94 -1.683041694060893e-12
C78_94 V78 V94 -3.761490432956219e-19

R78_95 V78 V95 6235.299321242131
L78_95 V78 V95 1.4019901924817436e-12
C78_95 V78 V95 4.820130382027915e-19

R78_96 V78 V96 14208.286605204048
L78_96 V78 V96 3.7403647383807534e-12
C78_96 V78 V96 2.3966524293734693e-19

R78_97 V78 V97 -40502.06097320528
L78_97 V78 V97 -3.5145672149932723e-12
C78_97 V78 V97 -2.0801846112964156e-19

R78_98 V78 V98 4909.492197568006
L78_98 V78 V98 1.3466825843270904e-12
C78_98 V78 V98 4.467717482430918e-19

R78_99 V78 V99 -15902.565429316084
L78_99 V78 V99 -5.335966286172705e-12
C78_99 V78 V99 -9.577001276608852e-20

R78_100 V78 V100 -35759.81258120186
L78_100 V78 V100 -4.657689930790692e-12
C78_100 V78 V100 -1.2847177243117065e-19

R78_101 V78 V101 6391.844896747462
L78_101 V78 V101 1.4470642473841899e-12
C78_101 V78 V101 4.754391380591496e-19

R78_102 V78 V102 3726.759172585213
L78_102 V78 V102 9.495803870410043e-13
C78_102 V78 V102 6.413772165293978e-19

R78_103 V78 V103 -20942.443569052164
L78_103 V78 V103 -4.091199145595238e-12
C78_103 V78 V103 -1.6201480487232176e-19

R78_104 V78 V104 -75850.08730564729
L78_104 V78 V104 -2.4564263171440626e-11
C78_104 V78 V104 7.239182472441873e-20

R78_105 V78 V105 -5136.308939482963
L78_105 V78 V105 -9.57235355092177e-13
C78_105 V78 V105 -6.625204479542052e-19

R78_106 V78 V106 3242.2181530939342
L78_106 V78 V106 6.27474490999075e-13
C78_106 V78 V106 1.0814336341011077e-18

R78_107 V78 V107 5891.853641414096
L78_107 V78 V107 1.4273865016412502e-12
C78_107 V78 V107 4.404167412217507e-19

R78_108 V78 V108 -7103.322893129361
L78_108 V78 V108 -1.5303027306584154e-12
C78_108 V78 V108 -4.396133065490566e-19

R78_109 V78 V109 -18585.703305587984
L78_109 V78 V109 -3.737433692887221e-12
C78_109 V78 V109 -1.3622605663607488e-19

R78_110 V78 V110 -3803.6041934046993
L78_110 V78 V110 -6.499082863138982e-13
C78_110 V78 V110 -1.0987507356375982e-18

R78_111 V78 V111 -7170.527031715172
L78_111 V78 V111 -1.6452670080288269e-12
C78_111 V78 V111 -3.935982369400735e-19

R78_112 V78 V112 3874.794084375508
L78_112 V78 V112 1.2636270687299454e-12
C78_112 V78 V112 4.397045120723294e-19

R78_113 V78 V113 7544.013665136036
L78_113 V78 V113 1.9613697645072543e-12
C78_113 V78 V113 2.683031779516178e-19

R78_114 V78 V114 4231.060773410362
L78_114 V78 V114 1.270177442698625e-12
C78_114 V78 V114 5.904146710828191e-19

R78_115 V78 V115 8855.287580563941
L78_115 V78 V115 3.1989953477050683e-12
C78_115 V78 V115 1.9553503156785642e-19

R78_116 V78 V116 -7650.460578546295
L78_116 V78 V116 -1.8732372150839368e-12
C78_116 V78 V116 -3.114266699302496e-19

R78_117 V78 V117 -11542.609736948807
L78_117 V78 V117 -2.231803116941616e-12
C78_117 V78 V117 -3.0109332620141977e-19

R78_118 V78 V118 -5214.332022936348
L78_118 V78 V118 -1.4425863983552515e-12
C78_118 V78 V118 -4.282055167400531e-19

R78_119 V78 V119 -4534.954449132333
L78_119 V78 V119 -1.3514228990397867e-12
C78_119 V78 V119 -5.112240155827734e-19

R78_120 V78 V120 28752.578518661438
L78_120 V78 V120 1.7588749689893113e-11
C78_120 V78 V120 -1.0014397249725294e-19

R78_121 V78 V121 8505.541127699238
L78_121 V78 V121 2.640382351525997e-12
C78_121 V78 V121 1.6984761835314117e-19

R78_122 V78 V122 3985.8695185165725
L78_122 V78 V122 2.849158416935096e-12
C78_122 V78 V122 9.937089058672886e-21

R78_123 V78 V123 23666.304893099365
L78_123 V78 V123 -5.74863641652809e-12
C78_123 V78 V123 -1.432285418215855e-19

R78_124 V78 V124 -67794.06405086363
L78_124 V78 V124 -5.37195046735532e-12
C78_124 V78 V124 -1.0887724041125926e-19

R78_125 V78 V125 -14975.987301839796
L78_125 V78 V125 -4.499917859714499e-12
C78_125 V78 V125 -9.225128666420709e-20

R78_126 V78 V126 -4481.9483903683495
L78_126 V78 V126 -3.748245697188561e-12
C78_126 V78 V126 9.34380634955457e-20

R78_127 V78 V127 5985.735958739754
L78_127 V78 V127 2.8468648186219853e-12
C78_127 V78 V127 9.498838769255332e-21

R78_128 V78 V128 -89933.18976735325
L78_128 V78 V128 -2.0807743001040583e-11
C78_128 V78 V128 -1.237445781522335e-19

R78_129 V78 V129 12417.539795181001
L78_129 V78 V129 -1.1417674423975188e-11
C78_129 V78 V129 -1.2769509266326169e-19

R78_130 V78 V130 -7733.6284390024075
L78_130 V78 V130 -5.168700433963218e-12
C78_130 V78 V130 -1.5510552928639992e-19

R78_131 V78 V131 -16894.606210232465
L78_131 V78 V131 5.102755541491846e-12
C78_131 V78 V131 1.4927076207848804e-19

R78_132 V78 V132 -19357.87793471144
L78_132 V78 V132 -5.89541993855639e-12
C78_132 V78 V132 -7.990312101572616e-20

R78_133 V78 V133 12822.902456509146
L78_133 V78 V133 3.1106170961516148e-12
C78_133 V78 V133 2.115694129424506e-19

R78_134 V78 V134 -20466.810798225288
L78_134 V78 V134 1.6292609876281728e-10
C78_134 V78 V134 3.431520356557617e-20

R78_135 V78 V135 9158.30425429319
L78_135 V78 V135 6.967072039812625e-12
C78_135 V78 V135 -4.2661502418101236e-20

R78_136 V78 V136 832139.5685591869
L78_136 V78 V136 5.7914822440953234e-12
C78_136 V78 V136 1.0312750995641367e-19

R78_137 V78 V137 -17340.82816610742
L78_137 V78 V137 -6.457636736867677e-12
C78_137 V78 V137 -8.554579945336881e-20

R78_138 V78 V138 -3550.948775696157
L78_138 V78 V138 -3.1394990956343e-12
C78_138 V78 V138 -9.728924198399927e-20

R78_139 V78 V139 4537.974378703891
L78_139 V78 V139 2.0414643468920823e-12
C78_139 V78 V139 7.917537386813646e-20

R78_140 V78 V140 -11193.546381821943
L78_140 V78 V140 -9.818863541830035e-12
C78_140 V78 V140 1.3610426136758006e-20

R78_141 V78 V141 -22096.638285703528
L78_141 V78 V141 -6.151263686922772e-12
C78_141 V78 V141 -2.8490320183854556e-20

R78_142 V78 V142 -8327.447611409967
L78_142 V78 V142 -2.5843585044402664e-12
C78_142 V78 V142 -1.811280802407733e-19

R78_143 V78 V143 -11748.066992261896
L78_143 V78 V143 -7.680832127512493e-12
C78_143 V78 V143 -4.173117093842812e-20

R78_144 V78 V144 16992.52324424975
L78_144 V78 V144 4.0744311324784474e-11
C78_144 V78 V144 -4.0126616189926e-20

R79_79 V79 0 -300.2828602273704
L79_79 V79 0 -3.3755448456478966e-12
C79_79 V79 0 1.6019997710858458e-19

R79_80 V79 V80 3525.148553526308
L79_80 V79 V80 9.485915623522994e-13
C79_80 V79 V80 7.524811502676447e-19

R79_81 V79 V81 44420.54979375804
L79_81 V79 V81 -5.9089850186820246e-12
C79_81 V79 V81 -2.8928587404902176e-20

R79_82 V79 V82 290212.2431816863
L79_82 V79 V82 7.0510960326098155e-12
C79_82 V79 V82 1.244895988864152e-19

R79_83 V79 V83 3448.2179657299926
L79_83 V79 V83 1.4628359578513017e-12
C79_83 V79 V83 4.916292028543536e-19

R79_84 V79 V84 -7083.634806704034
L79_84 V79 V84 -1.8595261331522616e-12
C79_84 V79 V84 -1.4441613453170218e-19

R79_85 V79 V85 -4628.478918905285
L79_85 V79 V85 -1.2211643576723453e-12
C79_85 V79 V85 -4.118634477193363e-19

R79_86 V79 V86 -12142.179115238028
L79_86 V79 V86 -1.3499232019431044e-11
C79_86 V79 V86 4.814151171115303e-22

R79_87 V79 V87 -6365.677429920125
L79_87 V79 V87 -1.6233570920986815e-12
C79_87 V79 V87 -4.0090283300279724e-19

R79_88 V79 V88 56787.47191109015
L79_88 V79 V88 1.1462233610835498e-11
C79_88 V79 V88 -3.4889913899874124e-20

R79_89 V79 V89 -6640.970107463679
L79_89 V79 V89 -1.014778327790624e-11
C79_89 V79 V89 -1.6088612068011422e-19

R79_90 V79 V90 2334.9049503696288
L79_90 V79 V90 6.975559499525521e-13
C79_90 V79 V90 8.089140070115081e-19

R79_91 V79 V91 13675.488200105934
L79_91 V79 V91 4.451909847692106e-12
C79_91 V79 V91 1.3609154841043412e-19

R79_92 V79 V92 8592.806597551838
L79_92 V79 V92 1.8159117205889718e-12
C79_92 V79 V92 3.6196667810887157e-19

R79_93 V79 V93 -3698879.8158283993
L79_93 V79 V93 -2.8851228353933836e-12
C79_93 V79 V93 -2.778634520658623e-19

R79_94 V79 V94 16003.737773081104
L79_94 V79 V94 1.0952678429736704e-11
C79_94 V79 V94 2.3058512175890593e-19

R79_95 V79 V95 7259.459272930301
L79_95 V79 V95 6.601669584828772e-12
C79_95 V79 V95 8.695964511983496e-20

R79_96 V79 V96 5980.501872838298
L79_96 V79 V96 1.6101310286309805e-12
C79_96 V79 V96 3.7003498520223274e-19

R79_97 V79 V97 12812.389311545703
L79_97 V79 V97 1.529730470303258e-12
C79_97 V79 V97 3.1774322925879484e-19

R79_98 V79 V98 -21772.261138404425
L79_98 V79 V98 2.142141965568214e-12
C79_98 V79 V98 2.8376104190300684e-19

R79_99 V79 V99 -3846.477789552007
L79_99 V79 V99 -1.6726915537289984e-12
C79_99 V79 V99 -1.3087367967414603e-19

R79_100 V79 V100 59597.70952110502
L79_100 V79 V100 1.4384752140206808e-11
C79_100 V79 V100 3.3373347162261386e-20

R79_101 V79 V101 -8062.373211110588
L79_101 V79 V101 -3.3320918359088566e-11
C79_101 V79 V101 -3.586954033959737e-20

R79_102 V79 V102 1466.9604668228858
L79_102 V79 V102 4.0595788097617197e-13
C79_102 V79 V102 1.524444056349606e-18

R79_103 V79 V103 -1890.3178389668292
L79_103 V79 V103 -6.102077100389281e-13
C79_103 V79 V103 -1.155562640768119e-18

R79_104 V79 V104 17289.0595120899
L79_104 V79 V104 4.049757207205148e-12
C79_104 V79 V104 1.9925995767525647e-19

R79_105 V79 V105 -5093.501671984453
L79_105 V79 V105 -1.136537086411247e-12
C79_105 V79 V105 -5.327915281539566e-19

R79_106 V79 V106 2097.7203045611564
L79_106 V79 V106 6.948972409176677e-13
C79_106 V79 V106 9.704143545045512e-19

R79_107 V79 V107 1934.8015124923843
L79_107 V79 V107 4.3519333538555217e-13
C79_107 V79 V107 1.5835937417538445e-18

R79_108 V79 V108 -2520.224803647717
L79_108 V79 V108 -5.935205505509491e-13
C79_108 V79 V108 -1.042464030651439e-18

R79_109 V79 V109 -3557.2488586792238
L79_109 V79 V109 -1.4366748793800154e-12
C79_109 V79 V109 -3.618523407540074e-19

R79_110 V79 V110 8062.7187479817285
L79_110 V79 V110 -2.758896843851071e-12
C79_110 V79 V110 -4.790558335413534e-19

R79_111 V79 V111 -1492.7929559511472
L79_111 V79 V111 -7.387579870441045e-13
C79_111 V79 V111 -6.845637882392015e-19

R79_112 V79 V112 4123.784195193346
L79_112 V79 V112 7.49860449218326e-13
C79_112 V79 V112 7.709733697996697e-19

R79_113 V79 V113 6014.575044970544
L79_113 V79 V113 1.6862043239046134e-12
C79_113 V79 V113 2.858969646343727e-19

R79_114 V79 V114 4910.141441207671
L79_114 V79 V114 1.7417961946938096e-12
C79_114 V79 V114 2.561503263354316e-19

R79_115 V79 V115 1918.0918869700324
L79_115 V79 V115 7.066373539912419e-13
C79_115 V79 V115 9.06512975614768e-19

R79_116 V79 V116 -3153.493401288435
L79_116 V79 V116 -8.671626262730774e-13
C79_116 V79 V116 -6.051210196228382e-19

R79_117 V79 V117 115843.38012867008
L79_117 V79 V117 -2.4571843713718404e-12
C79_117 V79 V117 -4.310830050852366e-19

R79_118 V79 V118 -9284.558775134716
L79_118 V79 V118 -1.6129410854093028e-12
C79_118 V79 V118 -3.284033730977004e-19

R79_119 V79 V119 -2090.999417645041
L79_119 V79 V119 -1.0157253206315718e-12
C79_119 V79 V119 -4.2914173283558764e-19

R79_120 V79 V120 1049.9424384106035
L79_120 V79 V120 9.77118620161149e-13
C79_120 V79 V120 -2.3870731866256485e-19

R79_121 V79 V121 -2747.1494210955593
L79_121 V79 V121 -4.853644630271425e-11
C79_121 V79 V121 1.0872365385700092e-19

R79_122 V79 V122 1705.6232351164845
L79_122 V79 V122 8.085133326900087e-13
C79_122 V79 V122 -4.3342397504901446e-20

R79_123 V79 V123 8275.80740629173
L79_123 V79 V123 2.9666851205125962e-12
C79_123 V79 V123 -1.6243674888250798e-20

R79_124 V79 V124 -6505.265395084685
L79_124 V79 V124 -3.0792227394351016e-12
C79_124 V79 V124 -1.7054072205086078e-19

R79_125 V79 V125 1442.2561310072415
L79_125 V79 V125 2.4007000592913067e-12
C79_125 V79 V125 -1.0354010529429454e-19

R79_126 V79 V126 -871.4121183543456
L79_126 V79 V126 -5.476493615295309e-13
C79_126 V79 V126 1.3394363098458425e-19

R79_127 V79 V127 941.7064109899943
L79_127 V79 V127 6.112226901973759e-13
C79_127 V79 V127 2.1113128874897747e-20

R79_128 V79 V128 17262.34352065561
L79_128 V79 V128 8.741277174626961e-12
C79_128 V79 V128 2.2981169803854812e-21

R79_129 V79 V129 2453.8288100298473
L79_129 V79 V129 1.5134448100342176e-12
C79_129 V79 V129 3.664176184331676e-20

R79_130 V79 V130 -2449.4506569172
L79_130 V79 V130 -9.491401686241119e-13
C79_130 V79 V130 -3.4298701009304225e-19

R79_131 V79 V131 -8936.510891482621
L79_131 V79 V131 -2.0630866163843e-11
C79_131 V79 V131 3.4263552443633613e-19

R79_132 V79 V132 -4321.355138480793
L79_132 V79 V132 -2.201140527223772e-12
C79_132 V79 V132 -3.9389542865201995e-20

R79_133 V79 V133 6214.399747573187
L79_133 V79 V133 2.652207386002846e-12
C79_133 V79 V133 2.585833767945196e-19

R79_134 V79 V134 -15954.904749474746
L79_134 V79 V134 -8.80092260510836e-12
C79_134 V79 V134 3.111979147657185e-20

R79_135 V79 V135 1605.806789565832
L79_135 V79 V135 1.0968936039011064e-12
C79_135 V79 V135 -1.7315937905317888e-19

R79_136 V79 V136 25398.707092742232
L79_136 V79 V136 1.1794460426050973e-10
C79_136 V79 V136 -2.5008030892460193e-20

R79_137 V79 V137 3109.6331420132124
L79_137 V79 V137 1.1770220744573265e-11
C79_137 V79 V137 -1.13462509561375e-19

R79_138 V79 V138 -1008.1950890919749
L79_138 V79 V138 -5.901191831736537e-13
C79_138 V79 V138 -6.579656616093383e-20

R79_139 V79 V139 698.4233034245401
L79_139 V79 V139 4.4361062586859995e-13
C79_139 V79 V139 2.0376222300936127e-19

R79_140 V79 V140 -3780.2688485641875
L79_140 V79 V140 -1.4100164298119514e-12
C79_140 V79 V140 -8.46359912152347e-20

R79_141 V79 V141 -5202.5986478556515
L79_141 V79 V141 -2.8292434889114474e-12
C79_141 V79 V141 -2.490581185228598e-20

R79_142 V79 V142 -2923.5749315652497
L79_142 V79 V142 -1.4503833615612674e-12
C79_142 V79 V142 -5.416948670243548e-20

R79_143 V79 V143 -1934.2389536851413
L79_143 V79 V143 -1.1615679898487035e-12
C79_143 V79 V143 -7.359692909866827e-20

R79_144 V79 V144 9571.108200817398
L79_144 V79 V144 1.7157164800389883e-12
C79_144 V79 V144 1.2383761554934006e-19

R80_80 V80 0 -408.21258966223166
L80_80 V80 0 -1.7244610175540924e-13
C80_80 V80 0 -3.068284830106572e-19

R80_81 V80 V81 3500.5426539728683
L80_81 V80 V81 6.86690500628371e-13
C80_81 V80 V81 8.894666844633835e-19

R80_82 V80 V82 -5958.339900153439
L80_82 V80 V82 -1.9601156077865167e-12
C80_82 V80 V82 -4.474466959088128e-19

R80_83 V80 V83 -3674.8425368901885
L80_83 V80 V83 -8.462376890309933e-13
C80_83 V80 V83 -7.092981692730818e-19

R80_84 V80 V84 3463.397912102008
L80_84 V80 V84 1.9363017527432002e-12
C80_84 V80 V84 3.862686751295787e-19

R80_85 V80 V85 2883.4597793345115
L80_85 V80 V85 9.628063060610002e-13
C80_85 V80 V85 7.300734360786707e-19

R80_86 V80 V86 8018.459300379459
L80_86 V80 V86 3.558585149817177e-12
C80_86 V80 V86 1.432467239354362e-19

R80_87 V80 V87 3559.6117204834386
L80_87 V80 V87 1.0198201431844668e-12
C80_87 V80 V87 7.020796411484835e-19

R80_88 V80 V88 9956.005525281138
L80_88 V80 V88 3.6534892687157615e-12
C80_88 V80 V88 1.5642909111759956e-19

R80_89 V80 V89 -2556.0123671029187
L80_89 V80 V89 -9.113200883051414e-13
C80_89 V80 V89 -7.888684238575092e-19

R80_90 V80 V90 -2446.3098050533595
L80_90 V80 V90 -8.011701671245022e-13
C80_90 V80 V90 -7.873449929055091e-19

R80_91 V80 V91 -13912.32319251536
L80_91 V80 V91 -3.401217841191706e-12
C80_91 V80 V91 -1.6735951300841773e-19

R80_92 V80 V92 -2691.7089629181874
L80_92 V80 V92 -5.634612993999422e-13
C80_92 V80 V92 -1.1902775750308053e-18

R80_93 V80 V93 7751.474352198237
L80_93 V80 V93 3.2747309030156067e-12
C80_93 V80 V93 2.2983636028832284e-21

R80_94 V80 V94 3399.8541538199993
L80_94 V80 V94 1.2356913265546867e-12
C80_94 V80 V94 3.181818150233062e-19

R80_95 V80 V95 -19755.307849568435
L80_95 V80 V95 -4.963832542298444e-12
C80_95 V80 V95 -1.9411042043583345e-19

R80_96 V80 V96 -3155.920344651295
L80_96 V80 V96 -5.629349564470222e-13
C80_96 V80 V96 -1.1393078197620991e-18

R80_97 V80 V97 -3323.8048620320205
L80_97 V80 V97 -2.0568257298787316e-12
C80_97 V80 V97 -1.6580002386073913e-19

R80_98 V80 V98 -1484.4463260599132
L80_98 V80 V98 -6.402030001234324e-13
C80_98 V80 V98 -7.357085568404446e-19

R80_99 V80 V99 4916.731433325655
L80_99 V80 V99 1.7111745355975085e-12
C80_99 V80 V99 2.2783220431948934e-19

R80_100 V80 V100 10070.166362289423
L80_100 V80 V100 2.4806909279219825e-12
C80_100 V80 V100 2.982819727766181e-19

R80_101 V80 V101 -2507.539582624493
L80_101 V80 V101 -7.83852766663195e-13
C80_101 V80 V101 -8.870931678419901e-19

R80_102 V80 V102 -1213.1804559895975
L80_102 V80 V102 -4.042836931787671e-13
C80_102 V80 V102 -1.6607225374054096e-18

R80_103 V80 V103 4005.826635560765
L80_103 V80 V103 9.473140703436992e-13
C80_103 V80 V103 8.394759043987958e-19

R80_104 V80 V104 -5450.401834477895
L80_104 V80 V104 -8.713615174321835e-13
C80_104 V80 V104 -8.81033337803431e-19

R80_105 V80 V105 2683.3620776346547
L80_105 V80 V105 7.355440683790388e-13
C80_105 V80 V105 8.582298850977638e-19

R80_106 V80 V106 -3759.9259949753227
L80_106 V80 V106 -6.416198567832533e-13
C80_106 V80 V106 -1.306290343050289e-18

R80_107 V80 V107 -1942.305312078789
L80_107 V80 V107 -5.328338772966668e-13
C80_107 V80 V107 -1.255855490942409e-18

R80_108 V80 V108 2189.308748319954
L80_108 V80 V108 4.3340627572333975e-13
C80_108 V80 V108 1.8006541504581417e-18

R80_109 V80 V109 -12061.571901134359
L80_109 V80 V109 -4.837284908631026e-12
C80_109 V80 V109 -9.70845711661316e-20

R80_110 V80 V110 4666.695392221863
L80_110 V80 V110 8.212596776426294e-13
C80_110 V80 V110 9.437820156509243e-19

R80_111 V80 V111 5429.153736369988
L80_111 V80 V111 1.136615224606518e-12
C80_111 V80 V111 6.57669417846452e-19

R80_112 V80 V112 -965.6422060267467
L80_112 V80 V112 -4.3237079706945915e-13
C80_112 V80 V112 -1.2608071643239683e-18

R80_113 V80 V113 -2918.100573751354
L80_113 V80 V113 -1.3198415608743302e-12
C80_113 V80 V113 -2.659933703806626e-19

R80_114 V80 V114 -3993.327594810087
L80_114 V80 V114 -1.290812845165937e-12
C80_114 V80 V114 -5.141440743434241e-19

R80_115 V80 V115 -3165.992724394504
L80_115 V80 V115 -9.376070882693985e-13
C80_115 V80 V115 -7.704760960604611e-19

R80_116 V80 V116 2005.1379917968352
L80_116 V80 V116 6.006963609822869e-13
C80_116 V80 V116 1.0638473937216157e-18

R80_117 V80 V117 5206.45151444254
L80_117 V80 V117 1.3517089347353226e-12
C80_117 V80 V117 5.955646865922842e-19

R80_118 V80 V118 3791.4991556886534
L80_118 V80 V118 1.311911731136137e-12
C80_118 V80 V118 3.410695497940729e-19

R80_119 V80 V119 4700.897216906521
L80_119 V80 V119 8.838915894647456e-13
C80_119 V80 V119 8.363835296262985e-19

R80_120 V80 V120 -39032.81101046536
L80_120 V80 V120 3.7048598358244386e-12
C80_120 V80 V120 4.932081123629834e-19

R80_121 V80 V121 -1571.6251279908302
L80_121 V80 V121 -1.4657899918972123e-12
C80_121 V80 V121 1.3682013114838926e-20

R80_122 V80 V122 -791.6501741133203
L80_122 V80 V122 -5.962117486695643e-13
C80_122 V80 V122 -5.8830613780697e-20

R80_123 V80 V123 -5049.884257333238
L80_123 V80 V123 -4.5440475121750145e-12
C80_123 V80 V123 1.8900304215428736e-20

R80_124 V80 V124 44446.33558395926
L80_124 V80 V124 1.70502416703621e-12
C80_124 V80 V124 4.001451827693791e-19

R80_125 V80 V125 1672.2908069253251
L80_125 V80 V125 1.1046242549715385e-12
C80_125 V80 V125 1.6495717634053318e-19

R80_126 V80 V126 966.9653160329532
L80_126 V80 V126 7.365543934503252e-13
C80_126 V80 V126 -1.335205860477987e-19

R80_127 V80 V127 -1489.8835720178683
L80_127 V80 V127 -9.918577766233677e-13
C80_127 V80 V127 3.614101892801348e-20

R80_128 V80 V128 186920.15477327828
L80_128 V80 V128 -8.379528528686722e-12
C80_128 V80 V128 7.066947991961285e-21

R80_129 V80 V129 -5056.939825699728
L80_129 V80 V129 -5.926182986528187e-12
C80_129 V80 V129 1.2074232239399963e-19

R80_130 V80 V130 2455.3605773721542
L80_130 V80 V130 1.1332459308696014e-12
C80_130 V80 V130 4.842131310443069e-19

R80_131 V80 V131 4809.658417527299
L80_131 V80 V131 5.493037367053876e-11
C80_131 V80 V131 -2.7018013208898826e-19

R80_132 V80 V132 3167.0196167547842
L80_132 V80 V132 1.4991921763940201e-12
C80_132 V80 V132 1.9688233581358266e-19

R80_133 V80 V133 11674.783042172394
L80_133 V80 V133 -2.552122918477948e-12
C80_133 V80 V133 -4.256560207880128e-19

R80_134 V80 V134 4646.499546670265
L80_134 V80 V134 2.894481633007987e-12
C80_134 V80 V134 -5.0882345369991705e-20

R80_135 V80 V135 -2325.972483357248
L80_135 V80 V135 -1.8451631513309328e-12
C80_135 V80 V135 1.7519954077143755e-19

R80_136 V80 V136 23174.86348706437
L80_136 V80 V136 -2.684327446678749e-11
C80_136 V80 V136 -6.755629054586145e-21

R80_137 V80 V137 2342.6449356213298
L80_137 V80 V137 1.3194577583291054e-12
C80_137 V80 V137 3.013607667362125e-19

R80_138 V80 V138 940.0739391695785
L80_138 V80 V138 7.072629266926976e-13
C80_138 V80 V138 1.1748849505429501e-19

R80_139 V80 V139 -1069.0027341152222
L80_139 V80 V139 -6.784328355433408e-13
C80_139 V80 V139 -1.6712658337558205e-19

R80_140 V80 V140 2109.1519099069733
L80_140 V80 V140 1.257080053338672e-12
C80_140 V80 V140 1.6651464035619054e-19

R80_141 V80 V141 4631.868489868631
L80_141 V80 V141 2.9796290797230003e-12
C80_141 V80 V141 -1.0813302314541381e-20

R80_142 V80 V142 2871.917769689747
L80_142 V80 V142 2.193310094050079e-12
C80_142 V80 V142 1.3038870247708308e-19

R80_143 V80 V143 4204.877228345898
L80_143 V80 V143 2.1391975813781787e-12
C80_143 V80 V143 9.15337815186192e-20

R80_144 V80 V144 -3475.6193503159416
L80_144 V80 V144 -1.3993450002207767e-12
C80_144 V80 V144 -1.493127227040204e-19

R81_81 V81 0 16370.316796358906
L81_81 V81 0 2.551492367326404e-13
C81_81 V81 0 7.639955244611038e-19

R81_82 V81 V82 14742.874639176844
L81_82 V81 V82 2.1359484534395074e-12
C81_82 V81 V82 1.621320069704913e-19

R81_83 V81 V83 5037.9726141451
L81_83 V81 V83 7.955080884182941e-13
C81_83 V81 V83 7.633918785752671e-19

R81_84 V81 V84 10015.654989173388
L81_84 V81 V84 3.8392437774492974e-12
C81_84 V81 V84 1.645733917781373e-19

R81_85 V81 V85 -13961.670921064871
L81_85 V81 V85 -1.3376822456629756e-12
C81_85 V81 V85 -3.219611206616135e-19

R81_86 V81 V86 18146.084145138157
L81_86 V81 V86 -4.292567582741456e-12
C81_86 V81 V86 3.3034840371621283e-20

R81_87 V81 V87 -12017.018576608709
L81_87 V81 V87 -1.6546456228366892e-12
C81_87 V81 V87 -3.455951285291712e-19

R81_88 V81 V88 -7590.956154060823
L81_88 V81 V88 -1.457006211028012e-12
C81_88 V81 V88 -4.682207790594815e-19

R81_89 V81 V89 6720.211082024471
L81_89 V81 V89 1.340559684575888e-12
C81_89 V81 V89 3.7676237841312305e-19

R81_90 V81 V90 -9491.259002985065
L81_90 V81 V90 -4.750679521502712e-12
C81_90 V81 V90 -7.989728703575156e-20

R81_91 V81 V91 -7243.004035651628
L81_91 V81 V91 -2.2946846517156384e-12
C81_91 V81 V91 -2.9822363975937135e-19

R81_92 V81 V92 1919.9696422261093
L81_92 V81 V92 3.720396611347993e-13
C81_92 V81 V92 1.6745483902342882e-18

R81_93 V81 V93 -86320.20002396996
L81_93 V81 V93 -3.4476602283945873e-12
C81_93 V81 V93 -1.5150119411094498e-19

R81_94 V81 V94 -5209.869309760534
L81_94 V81 V94 -8.452777301083319e-13
C81_94 V81 V94 -7.87948187929538e-19

R81_95 V81 V95 -109802.24248336011
L81_95 V81 V95 1.994062965611764e-11
C81_95 V81 V95 9.341281377201629e-21

R81_96 V81 V96 1595.5441108373384
L81_96 V81 V96 3.0548078744457676e-13
C81_96 V81 V96 1.947011550769601e-18

R81_97 V81 V97 -3602.8560577123935
L81_97 V81 V97 -9.871911145118975e-13
C81_97 V81 V97 -5.549230067945039e-19

R81_98 V81 V98 14630.925274580219
L81_98 V81 V98 9.619076444737282e-13
C81_98 V81 V98 5.671336162798039e-19

R81_99 V81 V99 52279.7085681554
L81_99 V81 V99 -4.558978918506288e-12
C81_99 V81 V99 -2.169392093827807e-19

R81_100 V81 V100 -4349.184009840387
L81_100 V81 V100 -8.615962249885248e-13
C81_100 V81 V100 -8.129349125203857e-19

R81_101 V81 V101 3954.8026166353893
L81_101 V81 V101 7.942718593728254e-13
C81_101 V81 V101 6.725045239334066e-19

R81_102 V81 V102 -5808.199021765206
L81_102 V81 V102 -2.1854353908065254e-11
C81_102 V81 V102 -1.2743182544372022e-19

R81_103 V81 V103 -426458.8640650249
L81_103 V81 V103 -1.1550212773072906e-11
C81_103 V81 V103 1.2789735799213466e-20

R81_104 V81 V104 1962.8956958740343
L81_104 V81 V104 4.233884576419596e-13
C81_104 V81 V104 1.5553081420900494e-18

R81_105 V81 V105 -5516.873639212901
L81_105 V81 V105 -8.291305468756043e-13
C81_105 V81 V105 -8.310123235435943e-19

R81_106 V81 V106 4684.779795635159
L81_106 V81 V106 8.977611650362201e-13
C81_106 V81 V106 6.424141783329887e-19

R81_107 V81 V107 -18594.798752126033
L81_107 V81 V107 7.767214448050681e-11
C81_107 V81 V107 -9.831961738846206e-20

R81_108 V81 V108 -3249.768290987148
L81_108 V81 V108 -7.914747050448722e-13
C81_108 V81 V108 -7.804322187285903e-19

R81_109 V81 V109 2451.9541767963
L81_109 V81 V109 5.368717976412016e-13
C81_109 V81 V109 1.4025322629100455e-18

R81_110 V81 V110 -3398.803882074534
L81_110 V81 V110 -8.72631129077382e-13
C81_110 V81 V110 -5.211332435605294e-19

R81_111 V81 V111 -49520.06760940659
L81_111 V81 V111 -2.1670368531931282e-12
C81_111 V81 V111 -3.1438723266349234e-19

R81_112 V81 V112 -33026.47289564814
L81_112 V81 V112 1.685480513224684e-12
C81_112 V81 V112 3.4901158388104915e-19

R81_113 V81 V113 -4491.253559916435
L81_113 V81 V113 -3.5838910517059734e-12
C81_113 V81 V113 -3.615458126834153e-19

R81_114 V81 V114 -29930.01044012467
L81_114 V81 V114 2.3744007389045645e-12
C81_114 V81 V114 3.255323165246186e-19

R81_115 V81 V115 -10497.349980015984
L81_115 V81 V115 -1.3760104840312636e-11
C81_115 V81 V115 -2.6609104287147678e-21

R81_116 V81 V116 -7532.649854922835
L81_116 V81 V116 -1.1751150188892369e-12
C81_116 V81 V116 -5.127873580561119e-19

R81_117 V81 V117 34085.67025412585
L81_117 V81 V117 3.526125607515303e-11
C81_117 V81 V117 1.9912769244306746e-19

R81_118 V81 V118 6410.700504223322
L81_118 V81 V118 5.305969086374615e-12
C81_118 V81 V118 1.8552742685294103e-19

R81_119 V81 V119 -7384.753555119759
L81_119 V81 V119 -1.0916988887831642e-12
C81_119 V81 V119 -6.620304262729669e-19

R81_120 V81 V120 -2163.7864085169645
L81_120 V81 V120 -9.44466439047703e-13
C81_120 V81 V120 -4.338354652119944e-19

R81_121 V81 V121 -7602.928036622476
L81_121 V81 V121 -4.061009249694259e-11
C81_121 V81 V121 -1.8916799317773258e-20

R81_122 V81 V122 -1697.3476064469933
L81_122 V81 V122 -2.4818450069591637e-12
C81_122 V81 V122 7.5347639281084e-20

R81_123 V81 V123 -4423.029004519738
L81_123 V81 V123 -5.0846503391050825e-12
C81_123 V81 V123 6.777513784718036e-20

R81_124 V81 V124 -6174.14520034424
L81_124 V81 V124 -1.297100661145622e-12
C81_124 V81 V124 -5.127375483532453e-19

R81_125 V81 V125 -24127.929598755625
L81_125 V81 V125 -2.4006072820513155e-12
C81_125 V81 V125 -5.3732405977574234e-20

R81_126 V81 V126 1494.7953322635854
L81_126 V81 V126 1.318132939714419e-12
C81_126 V81 V126 2.0942226082140765e-21

R81_127 V81 V127 -1976.7251670301418
L81_127 V81 V127 -1.7557941045041187e-12
C81_127 V81 V127 -1.085164728619414e-19

R81_128 V81 V128 -8819.75738196577
L81_128 V81 V128 7.839830666232394e-11
C81_128 V81 V128 -2.870363375941052e-20

R81_129 V81 V129 -2858.62981491598
L81_129 V81 V129 -1.8154267218374448e-12
C81_129 V81 V129 -1.2402588272145493e-19

R81_130 V81 V130 4431.46106635286
L81_130 V81 V130 6.1618531958602824e-12
C81_130 V81 V130 -1.2581463907520419e-19

R81_131 V81 V131 3560.0648918907987
L81_131 V81 V131 2.5971509191408223e-12
C81_131 V81 V131 6.12458611230722e-21

R81_132 V81 V132 -92925.0078309007
L81_132 V81 V132 -1.908837259036468e-12
C81_132 V81 V132 -3.571229455635395e-19

R81_133 V81 V133 7339.257696778247
L81_133 V81 V133 1.973231562410785e-12
C81_133 V81 V133 2.454394190884003e-19

R81_134 V81 V134 8377.835639610581
L81_134 V81 V134 1.1209886627099918e-10
C81_134 V81 V134 -3.460119019413892e-20

R81_135 V81 V135 -2904.161191334023
L81_135 V81 V135 -2.6141080761600753e-12
C81_135 V81 V135 -4.080670123716025e-20

R81_136 V81 V136 61075.23306079238
L81_136 V81 V136 3.694593644657097e-12
C81_136 V81 V136 1.2245896650210382e-19

R81_137 V81 V137 -14243.024175515638
L81_137 V81 V137 -3.1534106233680994e-12
C81_137 V81 V137 -2.148036768665108e-19

R81_138 V81 V138 1524.5640666427137
L81_138 V81 V138 1.2883587326901532e-12
C81_138 V81 V138 -5.038546646237955e-20

R81_139 V81 V139 -1627.998525709003
L81_139 V81 V139 -1.7286555939092865e-12
C81_139 V81 V139 6.267592687852686e-20

R81_140 V81 V140 7783.2227271578195
L81_140 V81 V140 2.834833014343401e-10
C81_140 V81 V140 -5.688155597503885e-20

R81_141 V81 V141 5695.89719366189
L81_141 V81 V141 5.835067978128039e-12
C81_141 V81 V141 1.1191771785191027e-19

R81_142 V81 V142 3797.0558230533475
L81_142 V81 V142 3.0685298754487067e-12
C81_142 V81 V142 -1.1169988234874018e-19

R81_143 V81 V143 4826.149729240948
L81_143 V81 V143 3.0124918626653373e-12
C81_143 V81 V143 -2.741878192205578e-20

R81_144 V81 V144 -13131.60700157424
L81_144 V81 V144 -1.3092866497119287e-10
C81_144 V81 V144 -8.018499867475425e-20

R82_82 V82 0 5131.682810352171
L82_82 V82 0 -1.8129644363512508e-13
C82_82 V82 0 -6.580317303595476e-19

R82_83 V82 V83 -1784.8497771528328
L82_83 V82 V83 -3.5381798336585187e-13
C82_83 V82 V83 -1.8403617929497373e-18

R82_84 V82 V84 13163.689232036608
L82_84 V82 V84 4.361075496879167e-12
C82_84 V82 V84 4.3893000779229004e-20

R82_85 V82 V85 3409.807276703422
L82_85 V82 V85 7.068115540310511e-13
C82_85 V82 V85 7.822302510634115e-19

R82_86 V82 V86 2961.324896723506
L82_86 V82 V86 6.609894737127903e-13
C82_86 V82 V86 8.97673056755841e-19

R82_87 V82 V87 2263.479270525013
L82_87 V82 V87 5.137543163738221e-13
C82_87 V82 V87 1.3007587211102101e-18

R82_88 V82 V88 7987.114363070909
L82_88 V82 V88 1.7628418493210835e-12
C82_88 V82 V88 3.7381783928434936e-19

R82_89 V82 V89 -2509.9236493183234
L82_89 V82 V89 -6.167865853270334e-13
C82_89 V82 V89 -9.6769217633215e-19

R82_90 V82 V90 -9039.091422918613
L82_90 V82 V90 -4.699646281914688e-12
C82_90 V82 V90 -1.3056772931958485e-19

R82_91 V82 V91 -1292.2307071623304
L82_91 V82 V91 -2.6696266606887366e-13
C82_91 V82 V91 -2.3224456537405227e-18

R82_92 V82 V92 -3098.5463701060544
L82_92 V82 V92 -5.781009409786508e-13
C82_92 V82 V92 -1.0579552016835426e-18

R82_93 V82 V93 14531.671334489876
L82_93 V82 V93 2.392841812454547e-12
C82_93 V82 V93 1.3810338687712436e-19

R82_94 V82 V94 2335.081994900191
L82_94 V82 V94 5.918974607799171e-13
C82_94 V82 V94 9.681080367225024e-19

R82_95 V82 V95 -2305.692816672646
L82_95 V82 V95 -4.972284647071706e-13
C82_95 V82 V95 -1.3084482934350384e-18

R82_96 V82 V96 -7002.253326865742
L82_96 V82 V96 -2.0335904530400663e-12
C82_96 V82 V96 -4.500376231419788e-19

R82_97 V82 V97 10655.998233702196
L82_97 V82 V97 1.0316509920836252e-12
C82_97 V82 V97 5.7186653444431075e-19

R82_98 V82 V98 -1921.510178336883
L82_98 V82 V98 -4.877200503100609e-13
C82_98 V82 V98 -1.1273066355649464e-18

R82_99 V82 V99 5602.688399441171
L82_99 V82 V99 3.106159553696744e-12
C82_99 V82 V99 2.1331596547503876e-19

R82_100 V82 V100 8955.60089939243
L82_100 V82 V100 1.8781104796012045e-12
C82_100 V82 V100 2.5632217447091727e-19

R82_101 V82 V101 -2159.900310730733
L82_101 V82 V101 -4.74712851385582e-13
C82_101 V82 V101 -1.2460907055218344e-18

R82_102 V82 V102 -2147.5331508103277
L82_102 V82 V102 -5.216037329183608e-13
C82_102 V82 V102 -1.1301534728777161e-18

R82_103 V82 V103 -55070.259235314974
L82_103 V82 V103 -3.826071104883725e-12
C82_103 V82 V103 -5.3020192822801973e-20

R82_104 V82 V104 7563.159890160812
L82_104 V82 V104 1.7727897727470418e-12
C82_104 V82 V104 2.1855098451882523e-19

R82_105 V82 V105 2202.948895159045
L82_105 V82 V105 4.167993597689547e-13
C82_105 V82 V105 1.444909576649929e-18

R82_106 V82 V106 -1332.45510859837
L82_106 V82 V106 -2.522383751018754e-13
C82_106 V82 V106 -2.6508173437822198e-18

R82_107 V82 V107 -3564.3165035656057
L82_107 V82 V107 -7.900746268628099e-13
C82_107 V82 V107 -8.601976255967204e-19

R82_108 V82 V108 3731.2308523352385
L82_108 V82 V108 6.544895878740158e-13
C82_108 V82 V108 9.768035826289621e-19

R82_109 V82 V109 7770.160160992989
L82_109 V82 V109 1.6569682966916087e-12
C82_109 V82 V109 4.114067029070506e-19

R82_110 V82 V110 1497.7203096619812
L82_110 V82 V110 2.511660433304108e-13
C82_110 V82 V110 2.5961395979961985e-18

R82_111 V82 V111 3384.9017108573735
L82_111 V82 V111 8.49870472338979e-13
C82_111 V82 V111 8.389171674266828e-19

R82_112 V82 V112 -1652.3642154927325
L82_112 V82 V112 -4.784624849363379e-13
C82_112 V82 V112 -1.094968052603848e-18

R82_113 V82 V113 -2377.158436404826
L82_113 V82 V113 -8.518457906612147e-13
C82_113 V82 V113 -6.120662971614386e-19

R82_114 V82 V114 -1983.0417100590532
L82_114 V82 V114 -4.984574532031345e-13
C82_114 V82 V114 -1.512363917205544e-18

R82_115 V82 V115 -6070.509512492495
L82_115 V82 V115 -2.042116492736023e-12
C82_115 V82 V115 -3.5904607853126283e-19

R82_116 V82 V116 3400.573033450228
L82_116 V82 V116 7.96007795323665e-13
C82_116 V82 V116 6.518803126209407e-19

R82_117 V82 V117 5117.516052348246
L82_117 V82 V117 9.36458515791339e-13
C82_117 V82 V117 6.061255606400761e-19

R82_118 V82 V118 1937.5938009600627
L82_118 V82 V118 4.937663894880868e-13
C82_118 V82 V118 1.2445538139114863e-18

R82_119 V82 V119 2090.5153167312783
L82_119 V82 V119 4.603102967737631e-13
C82_119 V82 V119 1.523030937965164e-18

R82_120 V82 V120 -5209.310431318969
L82_120 V82 V120 2.1005919180374337e-12
C82_120 V82 V120 3.1753831250433635e-19

R82_121 V82 V121 -3248.8953270811585
L82_121 V82 V121 -9.458340322081091e-13
C82_121 V82 V121 -3.183744629143533e-19

R82_122 V82 V122 -1312.5775259325212
L82_122 V82 V122 -1.7886017212678575e-12
C82_122 V82 V122 1.4695013735530515e-20

R82_123 V82 V123 -21796.861085825327
L82_123 V82 V123 1.4256893288780002e-12
C82_123 V82 V123 3.819484691029007e-19

R82_124 V82 V124 4656.070719101511
L82_124 V82 V124 1.630342280871997e-12
C82_124 V82 V124 3.4659984751404473e-19

R82_125 V82 V125 5180.30412911581
L82_125 V82 V125 9.594708082255717e-13
C82_125 V82 V125 2.6813925939595733e-19

R82_126 V82 V126 1361.384966366581
L82_126 V82 V126 3.020443902917865e-12
C82_126 V82 V126 -1.0577435180947707e-19

R82_127 V82 V127 -1851.3815667440267
L82_127 V82 V127 -2.532428863614107e-12
C82_127 V82 V127 -2.013152541108288e-21

R82_128 V82 V128 -7023.516636074306
L82_128 V82 V128 -1.3849258628548699e-11
C82_128 V82 V128 1.4487971504729686e-19

R82_129 V82 V129 -13317.49327584979
L82_129 V82 V129 3.037010396588488e-12
C82_129 V82 V129 1.8086716208533719e-19

R82_130 V82 V130 5128.56333409892
L82_130 V82 V130 2.12552976760704e-11
C82_130 V82 V130 3.091415239042914e-19

R82_131 V82 V131 10419.385127254576
L82_131 V82 V131 -2.2502090114196417e-12
C82_131 V82 V131 -1.9889609374806842e-19

R82_132 V82 V132 8260.29518833439
L82_132 V82 V132 3.931065845149748e-11
C82_132 V82 V132 -4.5755649367615807e-20

R82_133 V82 V133 -4313.577897789478
L82_133 V82 V133 -8.877152886072569e-13
C82_133 V82 V133 -7.542670767468435e-19

R82_134 V82 V134 6869.760784264677
L82_134 V82 V134 9.680549132851179e-12
C82_134 V82 V134 4.074876754471194e-20

R82_135 V82 V135 -2671.824852501578
L82_135 V82 V135 -2.7450469439502184e-11
C82_135 V82 V135 1.1136407729745325e-19

R82_136 V82 V136 -16495.749730923046
L82_136 V82 V136 -2.6052117050116858e-11
C82_136 V82 V136 3.627321583043079e-20

R82_137 V82 V137 4076.0238155231423
L82_137 V82 V137 1.3125120537581455e-12
C82_137 V82 V137 3.649158851371038e-19

R82_138 V82 V138 1429.7988832802841
L82_138 V82 V138 4.785805312382336e-12
C82_138 V82 V138 1.2018069910386416e-19

R82_139 V82 V139 -1343.3108436196972
L82_139 V82 V139 -2.077103472476409e-12
C82_139 V82 V139 -1.6059518781935696e-19

R82_140 V82 V140 5594.630274534326
L82_140 V82 V140 3.284936152326056e-12
C82_140 V82 V140 7.34726701620551e-20

R82_141 V82 V141 3438.8869582464536
L82_141 V82 V141 2.6779180034742955e-12
C82_141 V82 V141 9.331112158359969e-20

R82_142 V82 V142 4596.567516441503
L82_142 V82 V142 1.8413505600166377e-12
C82_142 V82 V142 3.3737928652802015e-19

R82_143 V82 V143 5201.874218736439
L82_143 V82 V143 2.407994532748827e-11
C82_143 V82 V143 5.747076239125728e-20

R82_144 V82 V144 -6562.084583614807
L82_144 V82 V144 -4.145194896486845e-12
C82_144 V82 V144 -7.175769730990156e-20

R83_83 V83 0 -3443.7579549551915
L83_83 V83 0 -1.9508890117327866e-13
C83_83 V83 0 -3.963265203616048e-19

R83_84 V83 V84 -55004.65913361562
L83_84 V83 V84 -7.337803835470577e-12
C83_84 V83 V84 -1.5710742722459222e-19

R83_85 V83 V85 4468.854599462544
L83_85 V83 V85 9.325328052545159e-13
C83_85 V83 V85 6.167454927320272e-19

R83_86 V83 V86 4251.8099688514285
L83_86 V83 V86 9.229836754580933e-13
C83_86 V83 V86 5.373779466350373e-19

R83_87 V83 V87 3030.9001081029737
L83_87 V83 V87 6.476653977267954e-13
C83_87 V83 V87 1.033646311991993e-18

R83_88 V83 V88 7916.445970768413
L83_88 V83 V88 1.7535486611711626e-12
C83_88 V83 V88 4.402216700119877e-19

R83_89 V83 V89 -20939.983796090193
L83_89 V83 V89 -1.569609226781073e-12
C83_89 V83 V89 -4.266659420380951e-19

R83_90 V83 V90 -7934.306604219353
L83_90 V83 V90 -1.687048362399237e-12
C83_90 V83 V90 -3.03796608648284e-19

R83_91 V83 V91 -2028.311684160281
L83_91 V83 V91 -3.8777376925727303e-13
C83_91 V83 V91 -1.5977383025543938e-18

R83_92 V83 V92 -2499.2224824245814
L83_92 V83 V92 -4.4007406817403086e-13
C83_92 V83 V92 -1.4201958061278928e-18

R83_93 V83 V93 13769.154343534017
L83_93 V83 V93 1.9037403197949938e-12
C83_93 V83 V93 3.442283326302666e-19

R83_94 V83 V94 8808.625965401072
L83_94 V83 V94 7.762531980845652e-13
C83_94 V83 V94 8.096903896003401e-19

R83_95 V83 V95 -3266.5838701527787
L83_95 V83 V95 -6.54164011278712e-13
C83_95 V83 V95 -9.36905572182057e-19

R83_96 V83 V96 -2870.5326655045733
L83_96 V83 V96 -5.879013213393215e-13
C83_96 V83 V96 -1.106528459931105e-18

R83_97 V83 V97 3938.541095354844
L83_97 V83 V97 9.497429725849111e-13
C83_97 V83 V97 5.603080051892229e-19

R83_98 V83 V98 -4953.689075315443
L83_98 V83 V98 -6.634876568789388e-13
C83_98 V83 V98 -9.832181953809952e-19

R83_99 V83 V99 158355.7379250744
L83_99 V83 V99 2.0591059922987e-12
C83_99 V83 V99 2.5959275285283104e-19

R83_100 V83 V100 7276.139091134828
L83_100 V83 V100 1.4772381878096752e-12
C83_100 V83 V100 4.216477581390462e-19

R83_101 V83 V101 -4126.70612564614
L83_101 V83 V101 -7.710813786182646e-13
C83_101 V83 V101 -7.924437443138061e-19

R83_102 V83 V102 -2901.2695369106204
L83_102 V83 V102 -5.262020134158461e-13
C83_102 V83 V102 -1.0861716536389964e-18

R83_103 V83 V103 3768.395439645545
L83_103 V83 V103 1.7640323943421315e-12
C83_103 V83 V103 3.4346944757376044e-19

R83_104 V83 V104 -8155.207756898924
L83_104 V83 V104 -1.947719182784569e-12
C83_104 V83 V104 -4.2005817065960355e-19

R83_105 V83 V105 2374.116533238595
L83_105 V83 V105 4.314824390502104e-13
C83_105 V83 V105 1.455852072560929e-18

R83_106 V83 V106 -1286.1624488335751
L83_106 V83 V106 -2.750145849413744e-13
C83_106 V83 V106 -2.3026560516962645e-18

R83_107 V83 V107 -2362.861893932742
L83_107 V83 V107 -5.813418527622855e-13
C83_107 V83 V107 -1.125169275803572e-18

R83_108 V83 V108 2602.0369892471103
L83_108 V83 V108 5.795237176314481e-13
C83_108 V83 V108 9.867107151502575e-19

R83_109 V83 V109 43089.693514392085
L83_109 V83 V109 9.355684900963532e-11
C83_109 V83 V109 -1.6584619896152972e-19

R83_110 V83 V110 1469.731811549525
L83_110 V83 V110 3.332097699559135e-13
C83_110 V83 V110 2.0123431943269314e-18

R83_111 V83 V111 2994.2960042190034
L83_111 V83 V111 6.085378098867436e-13
C83_111 V83 V111 9.092048920414273e-19

R83_112 V83 V112 -7474.573291993714
L83_112 V83 V112 -6.803493267011445e-13
C83_112 V83 V112 -9.346584806710843e-19

R83_113 V83 V113 -10933.8219519703
L83_113 V83 V113 -1.490056701428894e-12
C83_113 V83 V113 -3.0563512214091095e-19

R83_114 V83 V114 -3920.8932082127258
L83_114 V83 V114 -6.270858320882104e-13
C83_114 V83 V114 -1.182337307992821e-18

R83_115 V83 V115 -4945.487992668579
L83_115 V83 V115 -1.0237217762670477e-12
C83_115 V83 V115 -5.967792764664509e-19

R83_116 V83 V116 5959.051216483244
L83_116 V83 V116 7.78603379325068e-13
C83_116 V83 V116 6.615533118559393e-19

R83_117 V83 V117 6637.198607757302
L83_117 V83 V117 1.715689560808376e-12
C83_117 V83 V117 3.3164688956131287e-19

R83_118 V83 V118 4116.982289900465
L83_118 V83 V118 7.242393474200337e-13
C83_118 V83 V118 8.65496284951472e-19

R83_119 V83 V119 2410.973222223328
L83_119 V83 V119 4.4676186824373086e-13
C83_119 V83 V119 1.3771719274622544e-18

R83_120 V83 V120 4219.267327082468
L83_120 V83 V120 -3.1726254095165164e-11
C83_120 V83 V120 4.3396179666656e-19

R83_121 V83 V121 10360.119364041235
L83_121 V83 V121 -4.9598788267757324e-12
C83_121 V83 V121 -2.84817273898133e-19

R83_122 V83 V122 2146.8427218032784
L83_122 V83 V122 -6.811161153287156e-12
C83_122 V83 V122 1.8543338657004072e-20

R83_123 V83 V123 4279.725403249211
L83_123 V83 V123 1.766432568112139e-12
C83_123 V83 V123 2.7018286418996187e-19

R83_124 V83 V124 3743.8817692209655
L83_124 V83 V124 1.050163038387099e-12
C83_124 V83 V124 5.091531960209969e-19

R83_125 V83 V125 -13793.344969171305
L83_125 V83 V125 -1.0186224488966418e-11
C83_125 V83 V125 1.558762106738472e-19

R83_126 V83 V126 -2027.8957077573978
L83_126 V83 V126 2.5200430165079558e-12
C83_126 V83 V126 -1.4840996199164996e-19

R83_127 V83 V127 3829.8194747164057
L83_127 V83 V127 -1.4617955044692646e-12
C83_127 V83 V127 3.4715056405912974e-20

R83_128 V83 V128 -27288.690377895156
L83_128 V83 V128 -9.946224568895705e-12
C83_128 V83 V128 1.0632044890545329e-19

R83_129 V83 V129 4129.8313980473495
L83_129 V83 V129 4.4885351053387785e-12
C83_129 V83 V129 1.6339066019439608e-19

R83_130 V83 V130 -6552.930903963296
L83_130 V83 V130 4.503137548044665e-12
C83_130 V83 V130 2.9987369997822383e-19

R83_131 V83 V131 -2850.5716521708828
L83_131 V83 V131 -1.741801499089325e-12
C83_131 V83 V131 -2.6908623219094636e-19

R83_132 V83 V132 -16760.909802979466
L83_132 V83 V132 3.3201138069080158e-12
C83_132 V83 V132 9.671615025030273e-20

R83_133 V83 V133 -3043.844908390935
L83_133 V83 V133 -7.642777379166034e-13
C83_133 V83 V133 -7.292838525144775e-19

R83_134 V83 V134 -33413.12949128102
L83_134 V83 V134 -2.0719629623529372e-11
C83_134 V83 V134 2.7296540335274025e-20

R83_135 V83 V135 4084.1602133169476
L83_135 V83 V135 -4.7321484884973424e-12
C83_135 V83 V135 1.3787556424388634e-19

R83_136 V83 V136 -13091.641585015728
L83_136 V83 V136 -7.305471433694362e-12
C83_136 V83 V136 1.3324854373024702e-20

R83_137 V83 V137 36723.768250925685
L83_137 V83 V137 4.110680423415803e-12
C83_137 V83 V137 3.6010603034511935e-19

R83_138 V83 V138 -2309.0061841981837
L83_138 V83 V138 3.223528573277537e-12
C83_138 V83 V138 1.5268119802966568e-19

R83_139 V83 V139 4273.562086491712
L83_139 V83 V139 -9.877394067765783e-13
C83_139 V83 V139 -2.092579558762934e-19

R83_140 V83 V140 -6510.172664095177
L83_140 V83 V140 3.4285083078346203e-12
C83_140 V83 V140 8.254033053596569e-20

R83_141 V83 V141 -100888.69820710862
L83_141 V83 V141 4.237087641504375e-12
C83_141 V83 V141 2.0539436652832153e-20

R83_142 V83 V142 -6930.064316806765
L83_142 V83 V142 2.092795637190805e-12
C83_142 V83 V142 2.9955067481692295e-19

R83_143 V83 V143 -8394.014216207746
L83_143 V83 V143 4.522788345147524e-12
C83_143 V83 V143 3.565567340615123e-20

R83_144 V83 V144 10387.689163637107
L83_144 V83 V144 -2.898327172557247e-12
C83_144 V83 V144 -1.251160009300773e-19

R84_84 V84 0 826.6432713761857
L84_84 V84 0 3.668852995573702e-13
C84_84 V84 0 2.7345651263798675e-19

R84_85 V84 V85 -5259.639001315754
L84_85 V84 V85 -1.2872385231132061e-12
C84_85 V84 V85 -3.048296648938626e-19

R84_86 V84 V86 -10893.705413207017
L84_86 V84 V86 -4.086403219722527e-12
C84_86 V84 V86 -2.9389810866450804e-20

R84_87 V84 V87 -8044.812101838321
L84_87 V84 V87 -2.2507147196094103e-12
C84_87 V84 V87 -2.034623201627342e-19

R84_88 V84 V88 25348.906659160733
L84_88 V84 V88 1.0140328409873934e-11
C84_88 V84 V88 7.454437741145611e-20

R84_89 V84 V89 2900.351456109585
L84_89 V84 V89 1.130543727272954e-12
C84_89 V84 V89 4.757556643994141e-19

R84_90 V84 V90 7038.594870647084
L84_90 V84 V90 1.2368927940277752e-12
C84_90 V84 V90 3.373295411022868e-19

R84_91 V84 V91 1314541.573459499
L84_91 V84 V91 1.0762810108973185e-11
C84_91 V84 V91 -6.53425820109537e-20

R84_92 V84 V92 44169.57873700492
L84_92 V84 V92 -1.1164772132241257e-11
C84_92 V84 V92 -3.2292083762074824e-20

R84_93 V84 V93 12640.90271173487
L84_93 V84 V93 -2.460734388532904e-11
C84_93 V84 V93 1.773289960197548e-19

R84_94 V84 V94 10166.219095278248
L84_94 V84 V94 -1.4646073164275162e-11
C84_94 V84 V94 1.15956717143273e-19

R84_95 V84 V95 -37256.59973199834
L84_95 V84 V95 -2.942920015677309e-11
C84_95 V84 V95 8.829096265373182e-22

R84_96 V84 V96 -12106.944650253874
L84_96 V84 V96 -3.7112550709301406e-12
C84_96 V84 V96 -9.271760969228313e-20

R84_97 V84 V97 6464.550318646486
L84_97 V84 V97 1.1325538537568646e-12
C84_97 V84 V97 2.857454148203656e-19

R84_98 V84 V98 8610.328681000592
L84_98 V84 V98 1.2194353507045176e-12
C84_98 V84 V98 1.4193421950626194e-19

R84_99 V84 V99 7316.294770516825
L84_99 V84 V99 -5.662174792953644e-12
C84_99 V84 V99 1.1786295176358778e-22

R84_100 V84 V100 15845.257465601693
L84_100 V84 V100 6.496498638501731e-12
C84_100 V84 V100 7.733451176977559e-20

R84_101 V84 V101 3595.487937680338
L84_101 V84 V101 1.331589587447141e-12
C84_101 V84 V101 4.2084519819748736e-19

R84_102 V84 V102 2539.381126561273
L84_102 V84 V102 5.87584898820169e-13
C84_102 V84 V102 8.070094518732577e-19

R84_103 V84 V103 -11123.156050727406
L84_103 V84 V103 -1.9121724058525743e-12
C84_103 V84 V103 -3.39749719079005e-19

R84_104 V84 V104 21743.52365095203
L84_104 V84 V104 -3.5489964002799678e-12
C84_104 V84 V104 -5.3459485396687283e-20

R84_105 V84 V105 -29689.038661718267
L84_105 V84 V105 -3.827811759881377e-12
C84_105 V84 V105 2.4581044651847818e-21

R84_106 V84 V106 6225.291630947792
L84_106 V84 V106 4.404096361279871e-12
C84_106 V84 V106 2.0103928520874637e-19

R84_107 V84 V107 5026.0718735419205
L84_107 V84 V107 1.1250128639340356e-12
C84_107 V84 V107 3.6204767005272123e-19

R84_108 V84 V108 -2622.0837892972895
L84_108 V84 V108 -1.0569590356966168e-12
C84_108 V84 V108 -6.7207408262415275e-19

R84_109 V84 V109 -8150.52470363157
L84_109 V84 V109 -1.7237381469166013e-12
C84_109 V84 V109 -4.0857406709419936e-19

R84_110 V84 V110 -3292.5565351262326
L84_110 V84 V110 -3.3148541054158904e-12
C84_110 V84 V110 -1.722042758441444e-19

R84_111 V84 V111 5450.487927795252
L84_111 V84 V111 -1.337990534893677e-11
C84_111 V84 V111 -1.0758455083390223e-19

R84_112 V84 V112 3940.7099829692975
L84_112 V84 V112 6.031425468413404e-13
C84_112 V84 V112 5.382763559236374e-19

R84_113 V84 V113 55944.77540160184
L84_113 V84 V113 1.4438677269787314e-12
C84_113 V84 V113 2.306721472794326e-19

R84_114 V84 V114 11726.214433132414
L84_114 V84 V114 2.6615164496411083e-12
C84_114 V84 V114 1.1488954682264921e-19

R84_115 V84 V115 160992.0829870247
L84_115 V84 V115 2.288444792457525e-12
C84_115 V84 V115 2.1290830404371178e-19

R84_116 V84 V116 -7920.573502274748
L84_116 V84 V116 -1.3111760490859418e-12
C84_116 V84 V116 -3.879378329585019e-19

R84_117 V84 V117 -3049.73496034993
L84_117 V84 V117 -1.6445938491022424e-12
C84_117 V84 V117 -3.6634078297148622e-19

R84_118 V84 V118 -30488.899485538535
L84_118 V84 V118 -2.023406508390624e-12
C84_118 V84 V118 -1.0656447373134415e-19

R84_119 V84 V119 11576.28579359614
L84_119 V84 V119 -1.1369930016256931e-11
C84_119 V84 V119 -9.976118127183846e-20

R84_120 V84 V120 -1499.4630595253984
L84_120 V84 V120 -8.877400100855598e-12
C84_120 V84 V120 -8.330125897934476e-20

R84_121 V84 V121 8670.844570682637
L84_121 V84 V121 1.1113670002907956e-12
C84_121 V84 V121 -4.424950183064788e-20

R84_122 V84 V122 -2038.7727020430507
L84_122 V84 V122 6.279755471167109e-13
C84_122 V84 V122 3.015974952934627e-20

R84_123 V84 V123 -98726.51251157866
L84_123 V84 V123 3.0525281144658862e-12
C84_123 V84 V123 -2.1216517444573185e-21

R84_124 V84 V124 6080.650821506309
L84_124 V84 V124 4.201766992245749e-12
C84_124 V84 V124 4.233177443603296e-20

R84_125 V84 V125 -3050.4487808321887
L84_125 V84 V125 -9.677174503868067e-13
C84_125 V84 V125 -6.892090212986221e-20

R84_126 V84 V126 1137.497337447703
L84_126 V84 V126 -9.343067065542042e-13
C84_126 V84 V126 8.271368109218826e-20

R84_127 V84 V127 -1382.9744044342901
L84_127 V84 V127 1.4471243112085589e-12
C84_127 V84 V127 3.691265425939634e-21

R84_128 V84 V128 -9982.110672507777
L84_128 V84 V128 1.589369464317395e-11
C84_128 V84 V128 5.3260464977288e-20

R84_129 V84 V129 -5348.93799769926
L84_129 V84 V129 3.5454034083134864e-12
C84_129 V84 V129 -6.497647069029739e-20

R84_130 V84 V130 -11039.018977248013
L84_130 V84 V130 -1.562502501403491e-12
C84_130 V84 V130 -1.5149925586777352e-19

R84_131 V84 V131 10505.75893104268
L84_131 V84 V131 -4.319499781641433e-12
C84_131 V84 V131 1.1973177515255909e-19

R84_132 V84 V132 6093.533776380509
L84_132 V84 V132 -5.099670699980766e-12
C84_132 V84 V132 3.3582788726357753e-20

R84_133 V84 V133 -71157.84203659708
L84_133 V84 V133 -3.4989453207674807e-12
C84_133 V84 V133 -1.391198864692795e-20

R84_134 V84 V134 6108.46709083754
L84_134 V84 V134 -3.224411659791738e-12
C84_134 V84 V134 4.2367101074535384e-20

R84_135 V84 V135 -2004.0675794231886
L84_135 V84 V135 2.133694858334376e-12
C84_135 V84 V135 -1.944786555000949e-20

R84_136 V84 V136 -16566.594648542734
L84_136 V84 V136 -6.208158276855768e-12
C84_136 V84 V136 -5.001962575446115e-20

R84_137 V84 V137 -6447.151852002717
L84_137 V84 V137 -1.7126909482296158e-12
C84_137 V84 V137 -2.4045078779865487e-20

R84_138 V84 V138 1752.7995042397818
L84_138 V84 V138 -7.292894968525206e-13
C84_138 V84 V138 -1.0728556144477885e-19

R84_139 V84 V139 -1103.6576764920756
L84_139 V84 V139 1.0788677739205913e-12
C84_139 V84 V139 2.382569148273426e-20

R84_140 V84 V140 7873.510536419126
L84_140 V84 V140 -1.5341803704855102e-12
C84_140 V84 V140 -8.761825924330887e-20

R84_141 V84 V141 5711.286345160609
L84_141 V84 V141 -3.5236789542783647e-12
C84_141 V84 V141 -3.381804619366009e-20

R84_142 V84 V142 21914.63854817397
L84_142 V84 V142 -2.180258423347564e-12
C84_142 V84 V142 -1.384762241555706e-20

R84_143 V84 V143 3582.733514584639
L84_143 V84 V143 -3.84377144061544e-12
C84_143 V84 V143 -2.350599916863681e-20

R84_144 V84 V144 -17670.794088551374
L84_144 V84 V144 2.332792140823775e-12
C84_144 V84 V144 5.904953411596759e-20

R85_85 V85 0 -635.9304988527601
L85_85 V85 0 2.294545839610124e-13
C85_85 V85 0 8.84522743004181e-19

R85_86 V85 V86 -6673.021260968237
L85_86 V85 V86 -1.5421821099057009e-12
C85_86 V85 V86 -3.059335053787103e-19

R85_87 V85 V87 -3999.282432442999
L85_87 V85 V87 -9.409091303144306e-13
C85_87 V85 V87 -6.076841849915081e-19

R85_88 V85 V88 -39430.833029430585
L85_88 V85 V88 -4.5662540829193046e-12
C85_88 V85 V88 -1.3022726872752536e-19

R85_89 V85 V89 3081.062091144267
L85_89 V85 V89 9.76363540392797e-13
C85_89 V85 V89 5.800589433437407e-19

R85_90 V85 V90 4632.2339396366215
L85_90 V85 V90 1.0389602102333021e-12
C85_90 V85 V90 4.977506814698431e-19

R85_91 V85 V91 5274.136896148519
L85_91 V85 V91 1.0000197027615524e-12
C85_91 V85 V91 5.498300679063524e-19

R85_92 V85 V92 4737.788370552624
L85_92 V85 V92 9.805406014335778e-13
C85_92 V85 V92 5.771324107606526e-19

R85_93 V85 V93 -81181.65208467092
L85_93 V85 V93 -3.3500066009612718e-12
C85_93 V85 V93 -2.7733483256251446e-20

R85_94 V85 V94 -15078.40960536749
L85_94 V85 V94 -1.5354791614844809e-12
C85_94 V85 V94 -2.245434864025424e-19

R85_95 V85 V95 7749.113934679269
L85_95 V85 V95 1.7843452892894195e-12
C85_95 V85 V95 3.6774383640905363e-19

R85_96 V85 V96 6614.408401040237
L85_96 V85 V96 1.3206726067739672e-12
C85_96 V85 V96 4.493381817339998e-19

R85_97 V85 V97 36776.96025639666
L85_97 V85 V97 2.908892885691435e-12
C85_97 V85 V97 8.335911886256552e-20

R85_98 V85 V98 5268.525769691063
L85_98 V85 V98 7.388964160202685e-13
C85_98 V85 V98 5.571755276977791e-19

R85_99 V85 V99 -41282.64888160371
L85_99 V85 V99 -2.37479616779836e-12
C85_99 V85 V99 -1.2196060040320485e-19

R85_100 V85 V100 -72394.6036648883
L85_100 V85 V100 -4.040409793475221e-12
C85_100 V85 V100 -1.199988741219396e-19

R85_101 V85 V101 3210.097359713235
L85_101 V85 V101 8.277669551321713e-13
C85_101 V85 V101 6.902559904179644e-19

R85_102 V85 V102 1861.388549816985
L85_102 V85 V102 4.2281931719949575e-13
C85_102 V85 V102 1.323028602857449e-18

R85_103 V85 V103 -4113.253706230895
L85_103 V85 V103 -1.0979783359236385e-12
C85_103 V85 V103 -6.302766626647366e-19

R85_104 V85 V104 10840.725726792587
L85_104 V85 V104 3.277613899083189e-12
C85_104 V85 V104 2.85779727108708e-19

R85_105 V85 V105 -4936.952852081852
L85_105 V85 V105 -7.197092387738874e-13
C85_105 V85 V105 -7.371522749006439e-19

R85_106 V85 V106 2016.5178448077231
L85_106 V85 V106 5.127031005306017e-13
C85_106 V85 V106 1.2861036962073025e-18

R85_107 V85 V107 2689.486580439644
L85_107 V85 V107 6.3138664123981e-13
C85_107 V85 V107 9.176469890083478e-19

R85_108 V85 V108 -1977.5370863685198
L85_108 V85 V108 -5.56513334372216e-13
C85_108 V85 V108 -1.164922905216893e-18

R85_109 V85 V109 -6722.906262737339
L85_109 V85 V109 -2.9951759516611025e-12
C85_109 V85 V109 -2.412787380518113e-19

R85_110 V85 V110 -2362.9235294342407
L85_110 V85 V110 -6.273959093126735e-13
C85_110 V85 V110 -1.0490250094990325e-18

R85_111 V85 V111 -6988.71523424559
L85_111 V85 V111 -1.098813118522576e-12
C85_111 V85 V111 -5.575282583378568e-19

R85_112 V85 V112 2519.9536024845916
L85_112 V85 V112 4.81772261809999e-13
C85_112 V85 V112 9.280340248389796e-19

R85_113 V85 V113 6401.419274660092
L85_113 V85 V113 1.1020685927103426e-12
C85_113 V85 V113 3.7930139511979216e-19

R85_114 V85 V114 5248.89239658509
L85_114 V85 V114 1.0139928225789837e-12
C85_114 V85 V114 5.636715187347063e-19

R85_115 V85 V115 6068.209369594039
L85_115 V85 V115 1.269888873450053e-12
C85_115 V85 V115 4.850147115519334e-19

R85_116 V85 V116 -3522.533559879268
L85_116 V85 V116 -7.392755196838038e-13
C85_116 V85 V116 -7.124465923419492e-19

R85_117 V85 V117 -3428.119746197589
L85_117 V85 V117 -1.2088016585470355e-12
C85_117 V85 V117 -5.544884408588531e-19

R85_118 V85 V118 -7027.016976559887
L85_118 V85 V118 -9.814579515458551e-13
C85_118 V85 V118 -4.8116632017386475e-19

R85_119 V85 V119 -5250.686616305078
L85_119 V85 V119 -9.46160346188333e-13
C85_119 V85 V119 -6.530251451126813e-19

R85_120 V85 V120 -3608.2285095375373
L85_120 V85 V120 7.604812297967627e-11
C85_120 V85 V120 -2.380071797598129e-19

R85_121 V85 V121 25160.658116669903
L85_121 V85 V121 1.2385690359347169e-12
C85_121 V85 V121 9.140930365545502e-20

R85_122 V85 V122 -7635.525350739962
L85_122 V85 V122 6.833794549963968e-13
C85_122 V85 V122 2.76441599183749e-20

R85_123 V85 V123 -12909.65619638747
L85_123 V85 V123 7.383707509733597e-12
C85_123 V85 V123 -7.11217974774232e-20

R85_124 V85 V124 -26709.57137591659
L85_124 V85 V124 -4.073293277955628e-12
C85_124 V85 V124 -1.506010413719947e-19

R85_125 V85 V125 -7306.396715911241
L85_125 V85 V125 -1.141342472894865e-12
C85_125 V85 V125 -1.9438582963679974e-19

R85_126 V85 V126 3701.625540537961
L85_126 V85 V126 -8.423892621920141e-13
C85_126 V85 V126 1.352919469431953e-19

R85_127 V85 V127 -5227.24711260152
L85_127 V85 V127 1.0325343993278202e-12
C85_127 V85 V127 3.4310444627373596e-21

R85_128 V85 V128 -18567.20830136191
L85_128 V85 V128 1.6608270965596694e-11
C85_128 V85 V128 -7.37157415664819e-20

R85_129 V85 V129 -7079.8152792239325
L85_129 V85 V129 4.502098884555295e-12
C85_129 V85 V129 -7.593848798539631e-20

R85_130 V85 V130 -8660.619637707267
L85_130 V85 V130 -1.2516151434488753e-12
C85_130 V85 V130 -3.8036385832231116e-19

R85_131 V85 V131 7301.118006534425
L85_131 V85 V131 2.4563956555819724e-11
C85_131 V85 V131 2.3639267900546065e-19

R85_132 V85 V132 76858.36531742722
L85_132 V85 V132 -2.297695569490822e-12
C85_132 V85 V132 -9.176683459750528e-20

R85_133 V85 V133 7056.899143579869
L85_133 V85 V133 2.64802210777637e-12
C85_133 V85 V133 3.3860589330181066e-19

R85_134 V85 V134 10306.299424166991
L85_134 V85 V134 -3.617974326350932e-12
C85_134 V85 V134 2.347251103043838e-21

R85_135 V85 V135 -6175.247856509823
L85_135 V85 V135 1.8274429181794223e-12
C85_135 V85 V135 -9.374833830792032e-20

R85_136 V85 V136 -176569.59120423745
L85_136 V85 V136 8.252257398138826e-12
C85_136 V85 V136 7.838975558035646e-20

R85_137 V85 V137 -7881.976392799845
L85_137 V85 V137 -1.7162297106367194e-12
C85_137 V85 V137 -1.756912577868226e-19

R85_138 V85 V138 6755.744804059968
L85_138 V85 V138 -7.881157291371457e-13
C85_138 V85 V138 -9.308169785426839e-20

R85_139 V85 V139 -4848.026934552349
L85_139 V85 V139 7.298583065337749e-13
C85_139 V85 V139 1.5354501700703663e-19

R85_140 V85 V140 58923.463842683654
L85_140 V85 V140 -1.553584733273041e-12
C85_140 V85 V140 -7.457468530694118e-20

R85_141 V85 V141 65041.30420298284
L85_141 V85 V141 -2.5499259717289804e-12
C85_141 V85 V141 -3.50476386511447e-20

R85_142 V85 V142 35644.69683694257
L85_142 V85 V142 -1.7892557930108e-12
C85_142 V85 V142 -1.1302517388383452e-19

R85_143 V85 V143 14251.016872125889
L85_143 V85 V143 -2.496322906183583e-12
C85_143 V85 V143 -5.988459858988057e-20

R85_144 V85 V144 42430.933499689716
L85_144 V85 V144 2.8485547552089832e-12
C85_144 V85 V144 -2.6998066309236327e-20

R86_86 V86 0 5275.249474099035
L86_86 V86 0 3.925664271754976e-13
C86_86 V86 0 -4.061364646530079e-19

R86_87 V86 V87 -5409.969761094759
L86_87 V86 V87 -1.2720610544665727e-12
C86_87 V86 V87 -5.270755792300492e-19

R86_88 V86 V88 -69977.28580794376
L86_88 V86 V88 -4.775492680745597e-12
C86_88 V86 V88 -9.935863106650723e-20

R86_89 V86 V89 4549.8649206750015
L86_89 V86 V89 1.3663646591059514e-12
C86_89 V86 V89 4.2469561551201895e-19

R86_90 V86 V90 175345.19816894986
L86_90 V86 V90 9.823826539822097e-12
C86_90 V86 V90 1.8910385821750023e-20

R86_91 V86 V91 3180.4794310999655
L86_91 V86 V91 6.293478521560113e-13
C86_91 V86 V91 1.0686802651945464e-18

R86_92 V86 V92 12168.569243667056
L86_92 V86 V92 1.604840145157474e-12
C86_92 V86 V92 2.413192943318993e-19

R86_93 V86 V93 34536.65478250578
L86_93 V86 V93 -6.08600522248929e-12
C86_93 V86 V93 -1.2576309545643837e-20

R86_94 V86 V94 -128402.68534884036
L86_94 V86 V94 -1.654097119664919e-12
C86_94 V86 V94 -2.8055252508656965e-19

R86_95 V86 V95 6676.003543120022
L86_95 V86 V95 1.3243950479301904e-12
C86_95 V86 V95 4.990972485604667e-19

R86_96 V86 V96 -104516.28566720789
L86_96 V86 V96 1.2464700062088251e-11
C86_96 V86 V96 -3.1507877055844993e-20

R86_97 V86 V97 -10516.381224088735
L86_97 V86 V97 -3.274102003929836e-12
C86_97 V86 V97 -1.5358763966368226e-19

R86_98 V86 V98 15418.537746429101
L86_98 V86 V98 1.1709488410345558e-12
C86_98 V86 V98 3.676526422275772e-19

R86_99 V86 V99 9114.678788194675
L86_99 V86 V99 -2.5435196902777816e-11
C86_99 V86 V99 -3.2636895023636813e-20

R86_100 V86 V100 70507.06088504785
L86_100 V86 V100 -6.3279602429429144e-12
C86_100 V86 V100 1.9517032489249018e-20

R86_101 V86 V101 4174.89586692881
L86_101 V86 V101 1.0383511152104357e-12
C86_101 V86 V101 5.463647971552492e-19

R86_102 V86 V102 7059.784925419717
L86_102 V86 V102 1.5249757281636857e-12
C86_102 V86 V102 3.1595667275341346e-19

R86_103 V86 V103 -150544.433753364
L86_103 V86 V103 1.1199292848825009e-11
C86_103 V86 V103 3.34968959689981e-20

R86_104 V86 V104 -22491.421847894882
L86_104 V86 V104 -5.827368269382632e-12
C86_104 V86 V104 -1.7393827712134328e-19

R86_105 V86 V105 -9226.976547417631
L86_105 V86 V105 -1.0868997319472076e-12
C86_105 V86 V105 -4.934317174693713e-19

R86_106 V86 V106 2605.383108380804
L86_106 V86 V106 6.591291255860229e-13
C86_106 V86 V106 1.0340650217580334e-18

R86_107 V86 V107 10112.414671037826
L86_107 V86 V107 2.9116121564738777e-12
C86_107 V86 V107 2.0165679764250476e-19

R86_108 V86 V108 -4935.91888727288
L86_108 V86 V108 -1.8025604564066219e-12
C86_108 V86 V108 -3.057312465765899e-19

R86_109 V86 V109 -8173.931084304208
L86_109 V86 V109 -1.2042523634727175e-11
C86_109 V86 V109 -1.9998131278987084e-19

R86_110 V86 V110 -2161.632323482856
L86_110 V86 V110 -6.976568347857467e-13
C86_110 V86 V110 -8.914407764544137e-19

R86_111 V86 V111 19148.45105484391
L86_111 V86 V111 -4.211314559966622e-12
C86_111 V86 V111 -1.905897794777992e-19

R86_112 V86 V112 21793.21516153843
L86_112 V86 V112 1.097364964619821e-12
C86_112 V86 V112 3.955242860603183e-19

R86_113 V86 V113 31973.72781913343
L86_113 V86 V113 2.0466142171962807e-12
C86_113 V86 V113 2.819791535361556e-19

R86_114 V86 V114 7472.411728122027
L86_114 V86 V114 1.4654804280879734e-12
C86_114 V86 V114 4.6608640474099875e-19

R86_115 V86 V115 -29830.9622778061
L86_115 V86 V115 6.058317070051241e-12
C86_115 V86 V115 8.37935824751202e-20

R86_116 V86 V116 -24571.112998691457
L86_116 V86 V116 -2.1107220891344145e-12
C86_116 V86 V116 -1.9499288211913864e-19

R86_117 V86 V117 -4703.136216321007
L86_117 V86 V117 -1.8144503842646781e-12
C86_117 V86 V117 -3.248911790627761e-19

R86_118 V86 V118 -9607.078733774093
L86_118 V86 V118 -1.1808757939147456e-12
C86_118 V86 V118 -5.329708328464181e-19

R86_119 V86 V119 -11349.218231037374
L86_119 V86 V119 -1.352975007189139e-12
C86_119 V86 V119 -5.173796216551276e-19

R86_120 V86 V120 -2149.7629568604543
L86_120 V86 V120 -3.0700704099450595e-12
C86_120 V86 V120 -5.529184268234008e-20

R86_121 V86 V121 -31961.18704925315
L86_121 V86 V121 1.8832401466339133e-12
C86_121 V86 V121 9.60576644325889e-20

R86_122 V86 V122 -1710.789857344988
L86_122 V86 V122 2.5146242228413264e-12
C86_122 V86 V122 4.568486254089948e-20

R86_123 V86 V123 -6473.235781246769
L86_123 V86 V123 -1.6929784911032985e-11
C86_123 V86 V123 -4.485119204583829e-20

R86_124 V86 V124 25975.95397220143
L86_124 V86 V124 -8.143927757678055e-12
C86_124 V86 V124 -2.9849913061771674e-20

R86_125 V86 V125 -8209.65739615444
L86_125 V86 V125 -1.6862390967460924e-12
C86_125 V86 V125 -1.183521649106238e-19

R86_126 V86 V126 1269.5708555320284
L86_126 V86 V126 -3.288677604184866e-11
C86_126 V86 V126 5.865077463910034e-20

R86_127 V86 V127 -1715.347976978228
L86_127 V86 V127 1.53412399991306e-11
C86_127 V86 V127 2.0594616426274635e-20

R86_128 V86 V128 -11366.095242753194
L86_128 V86 V128 3.685032129147993e-11
C86_128 V86 V128 -1.0216645666405322e-19

R86_129 V86 V129 -4178.621303081297
L86_129 V86 V129 -1.20756550616935e-11
C86_129 V86 V129 -3.796192559049696e-20

R86_130 V86 V130 14164.477743105048
L86_130 V86 V130 -8.689251614420432e-12
C86_130 V86 V130 -2.0426575426406788e-19

R86_131 V86 V131 5439.909706535847
L86_131 V86 V131 2.959640487926184e-11
C86_131 V86 V131 -1.8139478136722367e-20

R86_132 V86 V132 6769.701662934915
L86_132 V86 V132 -1.0272571462811843e-10
C86_132 V86 V132 3.44805272426929e-20

R86_133 V86 V133 6771.910476963521
L86_133 V86 V133 1.798392577585334e-12
C86_133 V86 V133 4.2622894360826e-19

R86_134 V86 V134 7892.255759756766
L86_134 V86 V134 -1.0254977622950571e-11
C86_134 V86 V134 -6.457991172424894e-20

R86_135 V86 V135 -2431.613325792293
L86_135 V86 V135 -2.3650160769876e-10
C86_135 V86 V135 2.9140279808280108e-21

R86_136 V86 V136 -43251.02246916794
L86_136 V86 V136 1.0891639863132725e-11
C86_136 V86 V136 3.4526577663718144e-20

R86_137 V86 V137 -14393.449294737278
L86_137 V86 V137 -2.287742329970486e-12
C86_137 V86 V137 -1.7535599501408504e-19

R86_138 V86 V138 1559.212816734202
L86_138 V86 V138 3.1273843648982936e-11
C86_138 V86 V138 9.054660029522756e-20

R86_139 V86 V139 -1379.3341499593364
L86_139 V86 V139 8.76043016889724e-12
C86_139 V86 V139 1.054357124222195e-19

R86_140 V86 V140 5664.002891781249
L86_140 V86 V140 -1.6768881013919673e-11
C86_140 V86 V140 4.433259584830628e-21

R86_141 V86 V141 6959.365906696769
L86_141 V86 V141 -7.468586679668272e-12
C86_141 V86 V141 -1.4843721817190878e-20

R86_142 V86 V142 6837.064959600899
L86_142 V86 V142 -1.1894758343691164e-11
C86_142 V86 V142 -1.5232206948651838e-20

R86_143 V86 V143 4142.326447888088
L86_143 V86 V143 1.444038565685158e-11
C86_143 V86 V143 9.305025905342285e-21

R86_144 V86 V144 -11869.370132129166
L86_144 V86 V144 1.3816544340421663e-11
C86_144 V86 V144 7.976790359940855e-21

R87_87 V87 0 821.5006456673383
L87_87 V87 0 2.287269879634821e-13
C87_87 V87 0 1.6212796781014432e-19

R87_88 V87 V88 -11834.949546623355
L87_88 V87 V88 -2.364934277872578e-12
C87_88 V87 V88 -3.021851103499838e-19

R87_89 V87 V89 3313.150786468674
L87_89 V87 V89 1.05974654489966e-12
C87_89 V87 V89 6.191039286683654e-19

R87_90 V87 V90 6306.101472541677
L87_90 V87 V90 1.4641938583747744e-12
C87_90 V87 V90 3.324721423139353e-19

R87_91 V87 V91 2529.5428334440494
L87_91 V87 V91 5.680600646015836e-13
C87_91 V87 V91 1.2142050507145178e-18

R87_92 V87 V92 3363.7769743657477
L87_92 V87 V92 7.678251023681365e-13
C87_92 V87 V92 8.943716723782102e-19

R87_93 V87 V93 -18090.33107374888
L87_93 V87 V93 -2.540173550577432e-12
C87_93 V87 V93 -1.2611035812391915e-19

R87_94 V87 V94 -6694.568505127814
L87_94 V87 V94 -1.2393269845731626e-12
C87_94 V87 V94 -4.204438198019125e-19

R87_95 V87 V95 5414.0106750414325
L87_95 V87 V95 1.0814040951674279e-12
C87_95 V87 V95 6.803394004072063e-19

R87_96 V87 V96 7202.3645830058085
L87_96 V87 V96 1.2260619273965995e-12
C87_96 V87 V96 6.23530749578544e-19

R87_97 V87 V97 17512.81668138669
L87_97 V87 V97 -9.256289334563615e-12
C87_97 V87 V97 -2.180995733643591e-19

R87_98 V87 V98 2989.232930904286
L87_98 V87 V98 6.713388312249092e-13
C87_98 V87 V98 7.613109296009483e-19

R87_99 V87 V99 -214689.8788083321
L87_99 V87 V99 -2.6231512974859523e-12
C87_99 V87 V99 -1.4440367958141371e-19

R87_100 V87 V100 -34072.00320757417
L87_100 V87 V100 -2.8402070701664077e-12
C87_100 V87 V100 -2.2216424790295636e-19

R87_101 V87 V101 3110.219659335275
L87_101 V87 V101 7.029395354839113e-13
C87_101 V87 V101 9.279765786724805e-19

R87_102 V87 V102 1924.7774266609
L87_102 V87 V102 4.897894818169565e-13
C87_102 V87 V102 1.094972799141016e-18

R87_103 V87 V103 -10914.394328633538
L87_103 V87 V103 -1.5496097660620554e-12
C87_103 V87 V103 -4.494554193774145e-19

R87_104 V87 V104 13232.107865876924
L87_104 V87 V104 -2.3476108912640288e-11
C87_104 V87 V104 7.581727345566884e-20

R87_105 V87 V105 -2766.7063794930673
L87_105 V87 V105 -6.374997542571638e-13
C87_105 V87 V105 -9.471355149276609e-19

R87_106 V87 V106 1692.9512521041106
L87_106 V87 V106 4.136075487046949e-13
C87_106 V87 V106 1.774583634908848e-18

R87_107 V87 V107 2793.864331456523
L87_107 V87 V107 6.482748912200363e-13
C87_107 V87 V107 9.191706040126485e-19

R87_108 V87 V108 -2517.2196187648988
L87_108 V87 V108 -5.947689237089555e-13
C87_108 V87 V108 -1.0961032455145077e-18

R87_109 V87 V109 -23680.245788483586
L87_109 V87 V109 -2.469390268402691e-12
C87_109 V87 V109 -2.18307187429564e-19

R87_110 V87 V110 -1755.9569340595833
L87_110 V87 V110 -5.066477959577181e-13
C87_110 V87 V110 -1.4481684675228872e-18

R87_111 V87 V111 -12921.304390315096
L87_111 V87 V111 -1.009590760392503e-12
C87_111 V87 V111 -6.521716797684343e-19

R87_112 V87 V112 2201.8625297476
L87_112 V87 V112 4.789754612631273e-13
C87_112 V87 V112 1.0519553862503717e-18

R87_113 V87 V113 10102.679377808505
L87_113 V87 V113 1.1246670712107317e-12
C87_113 V87 V113 3.9638210762989467e-19

R87_114 V87 V114 2495.7443092881144
L87_114 V87 V114 7.836893226007938e-13
C87_114 V87 V114 8.892294718000466e-19

R87_115 V87 V115 6315.676546238121
L87_115 V87 V115 1.2428051609161808e-12
C87_115 V87 V115 4.972440093053264e-19

R87_116 V87 V116 -4241.349874669424
L87_116 V87 V116 -7.983474792600385e-13
C87_116 V87 V116 -6.742861065016527e-19

R87_117 V87 V117 -3892.1315533221427
L87_117 V87 V117 -1.2797594184587893e-12
C87_117 V87 V117 -4.918247849039476e-19

R87_118 V87 V118 -3851.6010139971054
L87_118 V87 V118 -8.085399021723341e-13
C87_118 V87 V118 -7.25209170422604e-19

R87_119 V87 V119 -3513.874720582382
L87_119 V87 V119 -6.751210414800216e-13
C87_119 V87 V119 -1.0492865663517705e-18

R87_120 V87 V120 -2570.8913166247735
L87_120 V87 V120 -8.954022970112835e-12
C87_120 V87 V120 -3.2538021844093393e-19

R87_121 V87 V121 4436.540064443913
L87_121 V87 V121 1.3227190999901584e-12
C87_121 V87 V121 1.4602014316955073e-19

R87_122 V87 V122 -164019.68492002942
L87_122 V87 V122 8.592522711617216e-13
C87_122 V87 V122 3.197642098042853e-20

R87_123 V87 V123 13337.400009457273
L87_123 V87 V123 1.458647814443683e-11
C87_123 V87 V123 -8.702707672962964e-20

R87_124 V87 V124 10070.053838230027
L87_124 V87 V124 -3.1857635391862024e-12
C87_124 V87 V124 -2.5427837939846975e-19

R87_125 V87 V125 -3485.3854852957475
L87_125 V87 V125 -1.3740866523617884e-12
C87_125 V87 V125 -1.7754326104698364e-19

R87_126 V87 V126 3623.483005639651
L87_126 V87 V126 -1.0969542099757722e-12
C87_126 V87 V126 1.411137680756668e-19

R87_127 V87 V127 -3821.7991811303473
L87_127 V87 V127 1.2768523741607803e-12
C87_127 V87 V127 -2.9623579070528955e-20

R87_128 V87 V128 -8068.939865172945
L87_128 V87 V128 5.9753565480794834e-12
C87_128 V87 V128 1.2044148384073988e-21

R87_129 V87 V129 22723.27145346281
L87_129 V87 V129 5.7297750604662785e-12
C87_129 V87 V129 -8.811156135351173e-20

R87_130 V87 V130 -3266.294601314348
L87_130 V87 V130 -1.7407669323654215e-12
C87_130 V87 V130 -3.08716404763312e-19

R87_131 V87 V131 -15237.34663076584
L87_131 V87 V131 6.835774186658605e-12
C87_131 V87 V131 2.3950536064757902e-19

R87_132 V87 V132 25793.163701596513
L87_132 V87 V132 -5.392499436996904e-12
C87_132 V87 V132 6.001141165230842e-20

R87_133 V87 V133 10417.500503828516
L87_133 V87 V133 1.5848353738557872e-12
C87_133 V87 V133 5.481399545155836e-19

R87_134 V87 V134 44445.4341570396
L87_134 V87 V134 -3.907739981002812e-12
C87_134 V87 V134 -4.2823267052225124e-20

R87_135 V87 V135 -5286.18282722241
L87_135 V87 V135 2.1893730257182805e-12
C87_135 V87 V135 -6.491250017839737e-20

R87_136 V87 V136 -11697.8562404127
L87_136 V87 V136 -9.602065046271656e-12
C87_136 V87 V136 -1.2363177851593403e-19

R87_137 V87 V137 -5510.278587697969
L87_137 V87 V137 -1.7439984739368649e-12
C87_137 V87 V137 -2.961692910542895e-19

R87_138 V87 V138 162466.30255826464
L87_138 V87 V138 -1.0163484239926288e-12
C87_138 V87 V138 -8.755075827976168e-20

R87_139 V87 V139 -3725.5002182580024
L87_139 V87 V139 8.953934387876455e-13
C87_139 V87 V139 1.5963674703265846e-19

R87_140 V87 V140 -17321.280359535325
L87_140 V87 V140 -1.5684950890867802e-12
C87_140 V87 V140 -1.3558882451417185e-19

R87_141 V87 V141 10233.297853327296
L87_141 V87 V141 -3.134341322628675e-12
C87_141 V87 V141 -4.0659764432966353e-20

R87_142 V87 V142 -4999.656314263014
L87_142 V87 V142 -1.8447777800638863e-12
C87_142 V87 V142 -1.2812765126609425e-19

R87_143 V87 V143 18197.665790941825
L87_143 V87 V143 -3.3759059236855344e-12
C87_143 V87 V143 -3.4711919684369127e-20

R87_144 V87 V144 21270.165737440006
L87_144 V87 V144 2.0608551445536976e-12
C87_144 V87 V144 1.3636268769355393e-19

R88_88 V88 0 -2285.2858568690117
L88_88 V88 0 6.65312336321291e-13
C88_88 V88 0 1.7134878832733449e-19

R88_89 V88 V89 204867.0378934015
L88_89 V88 V89 4.657617526909561e-12
C88_89 V88 V89 5.0753504388088884e-20

R88_90 V88 V90 -17795.639725667406
L88_90 V88 V90 -8.514581407591994e-12
C88_90 V88 V90 -5.122793998298826e-20

R88_91 V88 V91 11933.313686854173
L88_91 V88 V91 2.4576427576954644e-12
C88_91 V88 V91 2.913044703041602e-19

R88_92 V88 V92 5497.68390387644
L88_92 V88 V92 1.4040615254251265e-12
C88_92 V88 V92 5.175223191242667e-19

R88_93 V88 V93 5650.1316077222
L88_93 V88 V93 -7.2526450052572604e-12
C88_93 V88 V93 -1.1565157774523058e-19

R88_94 V88 V94 18351.0529171329
L88_94 V88 V94 -2.7071205304530733e-12
C88_94 V88 V94 -2.513495804181539e-19

R88_95 V88 V95 9845.66017855773
L88_95 V88 V95 3.867146395495081e-12
C88_95 V88 V95 1.8659049950587925e-19

R88_96 V88 V96 5732.335844347203
L88_96 V88 V96 1.414788409339962e-12
C88_96 V88 V96 5.358310953794077e-19

R88_97 V88 V97 -5089.170439027136
L88_97 V88 V97 -2.5646310705787414e-12
C88_97 V88 V97 -2.776737020991291e-19

R88_98 V88 V98 -4555.21115188142
L88_98 V88 V98 2.303076279534005e-12
C88_98 V88 V98 2.4592087168085454e-19

R88_99 V88 V99 24865.241599091278
L88_99 V88 V99 -7.147054713900774e-11
C88_99 V88 V99 -5.103287474829088e-20

R88_100 V88 V100 -21724.95738776451
L88_100 V88 V100 -3.066634483729967e-12
C88_100 V88 V100 -2.4701719334143787e-19

R88_101 V88 V101 15662.386334327015
L88_101 V88 V101 2.156599480671734e-12
C88_101 V88 V101 2.431869835845443e-19

R88_102 V88 V102 -32265.07900203751
L88_102 V88 V102 1.011275508887281e-11
C88_102 V88 V102 1.3236494210431204e-20

R88_103 V88 V103 -37417.163049662326
L88_103 V88 V103 -2.9097702764454915e-11
C88_103 V88 V103 -6.992798565857092e-20

R88_104 V88 V104 5354.991593884531
L88_104 V88 V104 3.0663082554548978e-12
C88_104 V88 V104 2.636131497042731e-19

R88_105 V88 V105 -10721.85865947863
L88_105 V88 V105 -2.01691923956006e-12
C88_105 V88 V105 -3.7768802765896807e-19

R88_106 V88 V106 2874.9775093004014
L88_106 V88 V106 1.3899061090931941e-12
C88_106 V88 V106 5.389059044188656e-19

R88_107 V88 V107 -23016.428294278197
L88_107 V88 V107 1.497954636599828e-11
C88_107 V88 V107 7.575878511348977e-20

R88_108 V88 V108 -3922.638091228625
L88_108 V88 V108 -3.4684259925060806e-12
C88_108 V88 V108 -1.7793536415311756e-19

R88_109 V88 V109 -54218.97370742918
L88_109 V88 V109 3.033801835303695e-12
C88_109 V88 V109 2.977103412766539e-19

R88_110 V88 V110 -5122.30929216536
L88_110 V88 V110 -1.4767527878386318e-12
C88_110 V88 V110 -4.408229267997534e-19

R88_111 V88 V111 -5639.689320740701
L88_111 V88 V111 -5.751492834676295e-12
C88_111 V88 V111 -1.9043560623995837e-19

R88_112 V88 V112 -3061.0587334516254
L88_112 V88 V112 2.8480836177849343e-12
C88_112 V88 V112 1.771291957906114e-19

R88_113 V88 V113 -4475.516765059369
L88_113 V88 V113 2.183887866972997e-11
C88_113 V88 V113 -3.0287794211537236e-20

R88_114 V88 V114 6849.216993771131
L88_114 V88 V114 2.695388071246446e-12
C88_114 V88 V114 2.839862216457662e-19

R88_115 V88 V115 26978.6548358152
L88_115 V88 V115 5.0973778197556776e-11
C88_115 V88 V115 6.057986129414452e-20

R88_116 V88 V116 -134080.36434072774
L88_116 V88 V116 -3.714847708489862e-12
C88_116 V88 V116 -1.396803744378694e-19

R88_117 V88 V117 140449.1364712359
L88_117 V88 V117 -1.1952045417944554e-11
C88_117 V88 V117 2.9594310185705636e-20

R88_118 V88 V118 15275.408291323307
L88_118 V88 V118 -5.38445052091152e-12
C88_118 V88 V118 -1.1373776458786498e-19

R88_119 V88 V119 -3397.8598835105704
L88_119 V88 V119 -2.1701947880484805e-12
C88_119 V88 V119 -3.78161053493717e-19

R88_120 V88 V120 23083.75163998646
L88_120 V88 V120 -3.727743826477699e-12
C88_120 V88 V120 -1.2571340767162416e-19

R88_121 V88 V121 -1766.790171619323
L88_121 V88 V121 5.902710628010975e-12
C88_121 V88 V121 6.598280002574004e-20

R88_122 V88 V122 -1218.9708112851433
L88_122 V88 V122 -8.400952674011916e-11
C88_122 V88 V122 2.35374320812935e-20

R88_123 V88 V123 -12969.86137740718
L88_123 V88 V123 -5.035227138941163e-11
C88_123 V88 V123 -3.719619267905908e-21

R88_124 V88 V124 -42902.53187722893
L88_124 V88 V124 -1.023788816198174e-11
C88_124 V88 V124 -1.441259083026916e-19

R88_125 V88 V125 1678.210328766492
L88_125 V88 V125 -5.6334880204301984e-12
C88_125 V88 V125 -3.032155941612408e-20

R88_126 V88 V126 1668.6157272414246
L88_126 V88 V126 4.860100068284862e-12
C88_126 V88 V126 5.062119232282123e-20

R88_127 V88 V127 -3202.698885497793
L88_127 V88 V127 -7.835049012224226e-12
C88_127 V88 V127 -3.0828580063611096e-20

R88_128 V88 V128 -11746.066514192466
L88_128 V88 V128 7.605924589930508e-11
C88_128 V88 V128 1.296788597908238e-20

R88_129 V88 V129 -31961.894212964904
L88_129 V88 V129 -9.792009421880198e-12
C88_129 V88 V129 -3.1863778921166997e-20

R88_130 V88 V130 -27525.843759089734
L88_130 V88 V130 4.671086501757662e-10
C88_130 V88 V130 -1.4922151316725067e-20

R88_131 V88 V131 9310.948792603194
L88_131 V88 V131 1.2274727229683197e-11
C88_131 V88 V131 5.203612626212666e-20

R88_132 V88 V132 8759.01951622249
L88_132 V88 V132 -2.922633131821653e-11
C88_132 V88 V132 -2.07181641379581e-20

R88_133 V88 V133 4931.439603610689
L88_133 V88 V133 4.6595331433268806e-12
C88_133 V88 V133 1.575343669254075e-19

R88_134 V88 V134 5753.592223348028
L88_134 V88 V134 4.785434500059381e-11
C88_134 V88 V134 -3.987787930468374e-20

R88_135 V88 V135 -4058.053493408202
L88_135 V88 V135 -3.394912231123887e-11
C88_135 V88 V135 2.0573914465050935e-20

R88_136 V88 V136 131545.92233433586
L88_136 V88 V136 -5.876588918177156e-11
C88_136 V88 V136 -2.753978705444615e-20

R88_137 V88 V137 2881.4441242869734
L88_137 V88 V137 -7.378466405400466e-12
C88_137 V88 V137 -9.564476112095817e-20

R88_138 V88 V138 1989.7972265025944
L88_138 V88 V138 1.0753385356679491e-11
C88_138 V88 V138 -5.143790698618197e-20

R88_139 V88 V139 -2732.229230660997
L88_139 V88 V139 -7.168055899503867e-12
C88_139 V88 V139 3.075769250815119e-20

R88_140 V88 V140 5682.259110729374
L88_140 V88 V140 -1.3007873251546106e-11
C88_140 V88 V140 -3.5050161890187583e-20

R88_141 V88 V141 4569.090715423446
L88_141 V88 V141 2.2655616736306772e-11
C88_141 V88 V141 1.705932714958594e-20

R88_142 V88 V142 362734.4032500153
L88_142 V88 V142 -2.185765459863147e-10
C88_142 V88 V142 -2.1191025963831112e-20

R88_143 V88 V143 42194.41697163169
L88_143 V88 V143 1.6806918992955177e-11
C88_143 V88 V143 -1.6969174276872074e-20

R88_144 V88 V144 -6057.435270021897
L88_144 V88 V144 3.483544585764591e-11
C88_144 V88 V144 1.0070582634984205e-20

R89_89 V89 0 632.8194912739057
L89_89 V89 0 -2.5295304617568916e-13
C89_89 V89 0 3.019074290179407e-19

R89_90 V89 V90 -8865.191146907759
L89_90 V89 V90 -2.723742378111055e-12
C89_90 V89 V90 -1.9173758659994733e-19

R89_91 V89 V91 -4301.289119351828
L89_91 V89 V91 -9.563906313442498e-13
C89_91 V89 V91 -6.534511182198876e-19

R89_92 V89 V92 -3938.072287284822
L89_92 V89 V92 -9.296822758151926e-13
C89_92 V89 V92 -6.752211354798482e-19

R89_93 V89 V93 -4944.460534228663
L89_93 V89 V93 -1.4957393821943176e-11
C89_93 V89 V93 -3.8690451945567454e-19

R89_94 V89 V94 2983.552645016419
L89_94 V89 V94 7.952143291010667e-13
C89_94 V89 V94 5.694870464903112e-19

R89_95 V89 V95 -5791.055744866486
L89_95 V89 V95 -2.095193967428191e-12
C89_95 V89 V95 -4.358168225264827e-19

R89_96 V89 V96 -8618.071502223558
L89_96 V89 V96 -2.1850699196024143e-12
C89_96 V89 V96 -3.7538330911410707e-19

R89_97 V89 V97 -11422.01165850367
L89_97 V89 V97 -2.481801146357026e-12
C89_97 V89 V97 3.353902041277108e-20

R89_98 V89 V98 -2457.853111645346
L89_98 V89 V98 -4.815533788110315e-13
C89_98 V89 V98 -6.75731908473106e-19

R89_99 V89 V99 9237.976701583792
L89_99 V89 V99 8.302032869123654e-12
C89_99 V89 V99 1.105465737443243e-19

R89_100 V89 V100 17922.288143179427
L89_100 V89 V100 3.6051506334783127e-12
C89_100 V89 V100 1.5556191097787998e-19

R89_101 V89 V101 -1374.9453366072912
L89_101 V89 V101 -4.4827218147519423e-13
C89_101 V89 V101 -1.3214304346670249e-18

R89_102 V89 V102 -2213.2027985296168
L89_102 V89 V102 -6.69250989508775e-13
C89_102 V89 V102 -8.231847290096658e-19

R89_103 V89 V103 -6183.622650247505
L89_103 V89 V103 -1.749992149501868e-12
C89_103 V89 V103 -2.0151731334640875e-19

R89_104 V89 V104 -11629.158115858512
L89_104 V89 V104 -4.1803334228484965e-12
C89_104 V89 V104 -2.7987004097661225e-19

R89_105 V89 V105 6108.6297068600215
L89_105 V89 V105 1.071205103880592e-12
C89_105 V89 V105 5.148298714407443e-19

R89_106 V89 V106 -3033.961836520827
L89_106 V89 V106 -1.1139928594514814e-12
C89_106 V89 V106 -9.596194802464414e-19

R89_107 V89 V107 18004.80345367939
L89_107 V89 V107 -2.9857431413703574e-12
C89_107 V89 V107 -7.537524291419724e-20

R89_108 V89 V108 1856.8551399983119
L89_108 V89 V108 7.903130578326326e-13
C89_108 V89 V108 1.1243899249555208e-18

R89_109 V89 V109 9841.883911779147
L89_109 V89 V109 -5.229691854763723e-12
C89_109 V89 V109 1.4091264942541976e-19

R89_110 V89 V110 2634.6987483635885
L89_110 V89 V110 5.590903889553208e-13
C89_110 V89 V110 1.077249461985575e-18

R89_111 V89 V111 -82732.41582279351
L89_111 V89 V111 -2.0023031293681658e-12
C89_111 V89 V111 1.4048072540739116e-19

R89_112 V89 V112 -1480.9732228737732
L89_112 V89 V112 -3.829090372478489e-13
C89_112 V89 V112 -9.375632716853234e-19

R89_113 V89 V113 -3817.4260012280624
L89_113 V89 V113 -1.042342536200973e-12
C89_113 V89 V113 -3.2909232080521913e-19

R89_114 V89 V114 -3051.3299242169755
L89_114 V89 V114 -1.1571547195505255e-12
C89_114 V89 V114 -6.170512552532695e-19

R89_115 V89 V115 67092.30123456095
L89_115 V89 V115 9.492056091344447e-12
C89_115 V89 V115 -5.0001464480541724e-20

R89_116 V89 V116 2644.297256106451
L89_116 V89 V116 9.066952201246998e-13
C89_116 V89 V116 6.418523767737524e-19

R89_117 V89 V117 3275.316771818992
L89_117 V89 V117 9.32371844039504e-13
C89_117 V89 V117 5.59881247179537e-19

R89_118 V89 V118 5183.839612327242
L89_118 V89 V118 1.0569501478486682e-12
C89_118 V89 V118 4.049811581789288e-19

R89_119 V89 V119 4049.5426527193617
L89_119 V89 V119 2.906969587779493e-12
C89_119 V89 V119 6.504424368527283e-19

R89_120 V89 V120 210789.38723571898
L89_120 V89 V120 6.455841162145637e-13
C89_120 V89 V120 2.711022428277655e-19

R89_121 V89 V121 -9089.270644902528
L89_121 V89 V121 -5.404244392808782e-13
C89_121 V89 V121 5.810391039917267e-20

R89_122 V89 V122 -1928.2379084085528
L89_122 V89 V122 -5.353273975307345e-13
C89_122 V89 V122 -1.1397919413342076e-19

R89_123 V89 V123 -9864.100373768284
L89_123 V89 V123 -1.358492445776215e-11
C89_123 V89 V123 9.902404861088475e-20

R89_124 V89 V124 423892.64630107215
L89_124 V89 V124 4.199547645583538e-11
C89_124 V89 V124 1.7176508212344266e-19

R89_125 V89 V125 6179.917923877642
L89_125 V89 V125 4.13195987541578e-13
C89_125 V89 V125 1.1415913728554641e-19

R89_126 V89 V126 2483.2887997239736
L89_126 V89 V126 2.523107325180269e-12
C89_126 V89 V126 -6.627240481339433e-20

R89_127 V89 V127 -4005.647896451885
L89_127 V89 V127 5.83675017957225e-12
C89_127 V89 V127 2.436837212041788e-20

R89_128 V89 V128 94330.10993129207
L89_128 V89 V128 3.270604316376658e-11
C89_128 V89 V128 5.446340404522614e-20

R89_129 V89 V129 -824500.6455423974
L89_129 V89 V129 2.27271845871076e-12
C89_129 V89 V129 2.417196037351665e-19

R89_130 V89 V130 3210.326334938413
L89_130 V89 V130 2.4383126914055263e-12
C89_130 V89 V130 2.9256276103221925e-19

R89_131 V89 V131 5397.137063979581
L89_131 V89 V131 4.225754748257555e-12
C89_131 V89 V131 -2.0353742555834208e-20

R89_132 V89 V132 8492.767195395367
L89_132 V89 V132 3.1774174341294916e-12
C89_132 V89 V132 8.480647462305374e-20

R89_133 V89 V133 -13563.359795522052
L89_133 V89 V133 2.933743794668915e-11
C89_133 V89 V133 -3.238964817015735e-19

R89_134 V89 V134 -56222.50496044316
L89_134 V89 V134 3.5673671614815544e-12
C89_134 V89 V134 -6.78791823393788e-20

R89_135 V89 V135 -4999.808300895134
L89_135 V89 V135 1.7538877105849853e-11
C89_135 V89 V135 4.15434020638458e-20

R89_136 V89 V136 49168.88160880637
L89_136 V89 V136 1.1290617063272182e-11
C89_136 V89 V136 -9.605848912409396e-21

R89_137 V89 V137 4578.8978191322685
L89_137 V89 V137 6.268522531211954e-13
C89_137 V89 V137 2.6485473411381603e-19

R89_138 V89 V138 2164.393958421007
L89_138 V89 V138 1.3085879199715272e-12
C89_138 V89 V138 8.199268688782425e-20

R89_139 V89 V139 -3023.1743531154375
L89_139 V89 V139 5.593635447989144e-12
C89_139 V89 V139 -2.857845536039124e-20

R89_140 V89 V140 5418.37029651324
L89_140 V89 V140 1.6744548684445807e-12
C89_140 V89 V140 1.0621937866728731e-19

R89_141 V89 V141 10582.551235084835
L89_141 V89 V141 3.4267195560752663e-12
C89_141 V89 V141 1.3711090225827538e-20

R89_142 V89 V142 4616.701695098809
L89_142 V89 V142 3.0147230490732863e-12
C89_142 V89 V142 1.594972618730875e-19

R89_143 V89 V143 9715.189611252745
L89_143 V89 V143 -3.477107132992094e-12
C89_143 V89 V143 1.3292933389517308e-21

R89_144 V89 V144 -6830.772495948194
L89_144 V89 V144 -1.886590696930199e-12
C89_144 V89 V144 -1.0006056853324345e-19

R90_90 V90 0 -382.5135882257801
L90_90 V90 0 -6.683465462052533e-13
C90_90 V90 0 -3.328592549317901e-19

R90_91 V90 V91 133466.76184889284
L90_91 V90 V91 -3.2431830409385406e-12
C90_91 V90 V91 -7.599984616631698e-20

R90_92 V90 V92 -13268.013335962867
L90_92 V90 V92 -2.753000485456375e-12
C90_92 V90 V92 -2.44023444759526e-19

R90_93 V90 V93 -18719.258711125945
L90_93 V90 V93 3.6469559897228025e-12
C90_93 V90 V93 7.723906448358151e-20

R90_94 V90 V94 -2403.538672657968
L90_94 V90 V94 -2.7409182597230886e-11
C90_94 V90 V94 -1.8962575486876128e-19

R90_95 V90 V95 35195.14052310943
L90_95 V90 V95 -6.858049742516486e-12
C90_95 V90 V95 -7.653652535084148e-20

R90_96 V90 V96 -38564.348330991495
L90_96 V90 V96 -3.800059745425449e-12
C90_96 V90 V96 -1.8561129091872807e-19

R90_97 V90 V97 -32334.423834315807
L90_97 V90 V97 -9.275762142612055e-13
C90_97 V90 V97 -4.1931614602418725e-19

R90_98 V90 V98 8441.825253178298
L90_98 V90 V98 -1.1938633535390854e-12
C90_98 V90 V98 -2.9353952642306964e-19

R90_99 V90 V99 -2973.2656736702
L90_99 V90 V99 1.6999296008581544e-12
C90_99 V90 V99 9.62791588912623e-20

R90_100 V90 V100 -11545.46569363189
L90_100 V90 V100 -4.929256367919495e-12
C90_100 V90 V100 -1.0374668439949411e-19

R90_101 V90 V101 -5278.254373922578
L90_101 V90 V101 -3.0732470328058384e-12
C90_101 V90 V101 -1.9753069813773442e-19

R90_102 V90 V102 -1680.8731844607885
L90_102 V90 V102 -3.288222878186624e-13
C90_102 V90 V102 -1.6596348127685648e-18

R90_103 V90 V103 1970.0145408391188
L90_103 V90 V103 6.181615180471116e-13
C90_103 V90 V103 1.0315487310987286e-18

R90_104 V90 V104 -6732.1987137662345
L90_104 V90 V104 -1.2252700884859481e-11
C90_104 V90 V104 -1.734882144463687e-19

R90_105 V90 V105 7596.727715563211
L90_105 V90 V105 1.0802735735241208e-12
C90_105 V90 V105 4.287101123002199e-19

R90_106 V90 V106 -1852.4986355372546
L90_106 V90 V106 -7.422846450145315e-13
C90_106 V90 V106 -8.330994269636973e-19

R90_107 V90 V107 -1527.8885504342777
L90_107 V90 V107 -4.1288741316196435e-13
C90_107 V90 V107 -1.376813265002493e-18

R90_108 V90 V108 1349.9628484825546
L90_108 V90 V108 5.344653696594763e-13
C90_108 V90 V108 1.1418633452241767e-18

R90_109 V90 V109 3790.4009691934148
L90_109 V90 V109 1.099814309024483e-12
C90_109 V90 V109 4.944635469324238e-19

R90_110 V90 V110 1443.2842896578516
L90_110 V90 V110 1.8101721424841753e-12
C90_110 V90 V110 4.94378465876777e-19

R90_111 V90 V111 -12488.770868952477
L90_111 V90 V111 8.738731701928573e-13
C90_111 V90 V111 5.38002385893342e-19

R90_112 V90 V112 18806.315702406657
L90_112 V90 V112 -5.037761833703614e-13
C90_112 V90 V112 -8.452016957377429e-19

R90_113 V90 V113 6593.262681668737
L90_113 V90 V113 -1.0570531443084491e-12
C90_113 V90 V113 -3.724334675969576e-19

R90_114 V90 V114 40066.33006077151
L90_114 V90 V114 -1.5112274630382684e-12
C90_114 V90 V114 -2.2055877909622975e-19

R90_115 V90 V115 -7609.2159934803085
L90_115 V90 V115 -6.737922241606961e-13
C90_115 V90 V115 -8.013478797005955e-19

R90_116 V90 V116 10334.74156502443
L90_116 V90 V116 7.169117486139662e-13
C90_116 V90 V116 6.800603384468583e-19

R90_117 V90 V117 1972.3392810757211
L90_117 V90 V117 1.2576243069474184e-12
C90_117 V90 V117 5.924026228063733e-19

R90_118 V90 V118 -26247.38114547293
L90_118 V90 V118 1.2043033328448922e-12
C90_118 V90 V118 3.069514275449322e-19

R90_119 V90 V119 -12662.67252178664
L90_119 V90 V119 1.1684942268187719e-12
C90_119 V90 V119 3.5206522457630153e-19

R90_120 V90 V120 736.5346651178181
L90_120 V90 V120 -1.1932612951784463e-12
C90_120 V90 V120 2.0386071400238876e-19

R90_121 V90 V121 4282.078690630434
L90_121 V90 V121 -1.923679540615403e-12
C90_121 V90 V121 -6.543743709151521e-20

R90_122 V90 V122 503.39826433828483
L90_122 V90 V122 -4.978416101841406e-13
C90_122 V90 V122 -2.6377374085702036e-21

R90_123 V90 V123 2570.4242815013026
L90_123 V90 V123 -2.380108031080096e-12
C90_123 V90 V123 4.293289470787531e-20

R90_124 V90 V124 -11767.810171246121
L90_124 V90 V124 4.963020098067383e-12
C90_124 V90 V124 1.0889386549539659e-19

R90_125 V90 V125 4893.185508665691
L90_125 V90 V125 4.6157664824124356e-12
C90_125 V90 V125 1.0134786786054008e-19

R90_126 V90 V126 -396.60289964714633
L90_126 V90 V126 4.622347904068259e-13
C90_126 V90 V126 -1.437229648631618e-19

R90_127 V90 V127 551.427573506672
L90_127 V90 V127 -5.624524754807406e-13
C90_127 V90 V127 -1.7511381403204045e-20

R90_128 V90 V128 5453.881187250446
L90_128 V90 V128 -1.5203085495277843e-11
C90_128 V90 V128 3.07109831565411e-20

R90_129 V90 V129 1508.1497238296904
L90_129 V90 V129 -1.5668250047586409e-12
C90_129 V90 V129 5.378516621197161e-20

R90_130 V90 V130 -3655.2143470108995
L90_130 V90 V130 7.554292987864022e-13
C90_130 V90 V130 3.684163924878982e-19

R90_131 V90 V131 -1348.882053362292
L90_131 V90 V131 7.774516212565126e-12
C90_131 V90 V131 -3.416229687427409e-19

R90_132 V90 V132 -2235.244408972994
L90_132 V90 V132 1.7716511979599803e-12
C90_132 V90 V132 7.518634982805156e-20

R90_133 V90 V133 -4593.371449878658
L90_133 V90 V133 -6.443006654310681e-12
C90_133 V90 V133 -1.7667968767107274e-19

R90_134 V90 V134 -2557.0653293347673
L90_134 V90 V134 3.8010794338402265e-12
C90_134 V90 V134 -6.977992851264027e-20

R90_135 V90 V135 757.2486334276559
L90_135 V90 V135 -9.763786109230556e-13
C90_135 V90 V135 1.341006264093404e-19

R90_136 V90 V136 27688.46183142983
L90_136 V90 V136 -4.1083877923409904e-11
C90_136 V90 V136 -3.1978800973199975e-20

R90_137 V90 V137 43392.33208202985
L90_137 V90 V137 3.970284280797651e-12
C90_137 V90 V137 6.633464962167641e-20

R90_138 V90 V138 -496.14086116132813
L90_138 V90 V138 4.445931780223486e-13
C90_138 V90 V138 1.1085593058296826e-19

R90_139 V90 V139 443.415838451928
L90_139 V90 V139 -4.1132801851544284e-13
C90_139 V90 V139 -1.2849604913335995e-19

R90_140 V90 V140 -1774.7263831112186
L90_140 V90 V140 1.093376226483569e-12
C90_140 V90 V140 8.034783666581115e-20

R90_141 V90 V141 -2108.1622566484843
L90_141 V90 V141 2.05504727139483e-12
C90_141 V90 V141 2.9375838596638276e-20

R90_142 V90 V142 -1964.0869054954446
L90_142 V90 V142 1.0916265429083676e-12
C90_142 V90 V142 9.694764418195515e-20

R90_143 V90 V143 -1376.7303867444227
L90_143 V90 V143 1.078023481698305e-12
C90_143 V90 V143 9.997784081137478e-20

R90_144 V90 V144 3098.413155313115
L90_144 V90 V144 -1.420672101565482e-12
C90_144 V90 V144 -1.1884826652901544e-19

R91_91 V91 0 -637.8692710525714
L91_91 V91 0 -5.446465969064738e-13
C91_91 V91 0 9.666649505611709e-19

R91_92 V91 V92 -5264.547307765666
L91_92 V91 V92 -9.156003832261994e-13
C91_92 V91 V92 -6.460417495918116e-19

R91_93 V91 V93 26434.835642013524
L91_93 V91 V93 2.4070488292910504e-12
C91_93 V91 V93 1.9882983506845249e-19

R91_94 V91 V94 9206.851520914826
L91_94 V91 V94 9.122827967809544e-13
C91_94 V91 V94 6.584006441689074e-19

R91_95 V91 V95 -2773.3152498764453
L91_95 V91 V95 -5.10649269972613e-13
C91_95 V91 V95 -1.2870605365079603e-18

R91_96 V91 V96 21624.20311600588
L91_96 V91 V96 3.643607616537383e-12
C91_96 V91 V96 4.3804179161275637e-20

R91_97 V91 V97 7656.506483690498
L91_97 V91 V97 1.315934399907853e-12
C91_97 V91 V97 4.891940845071623e-19

R91_98 V91 V98 -4493.544905718216
L91_98 V91 V98 -6.700012190428869e-13
C91_98 V91 V98 -8.505803839510749e-19

R91_99 V91 V99 -9045.376146241177
L91_99 V91 V99 6.185841140704018e-12
C91_99 V91 V99 7.578718399324136e-20

R91_100 V91 V100 -68814.06252617414
L91_100 V91 V100 5.9460598006874595e-12
C91_100 V91 V100 -1.9031095292959495e-20

R91_101 V91 V101 -3240.4099974132746
L91_101 V91 V101 -6.863657621706155e-13
C91_101 V91 V101 -9.174420213209845e-19

R91_102 V91 V102 -3224.927410627616
L91_102 V91 V102 -5.874331567621519e-13
C91_102 V91 V102 -7.749878295446256e-19

R91_103 V91 V103 -24542.39856243622
L91_103 V91 V103 -1.0993336445890485e-11
C91_103 V91 V103 -5.300840764349618e-20

R91_104 V91 V104 5945.317374300474
L91_104 V91 V104 9.804126801390094e-13
C91_104 V91 V104 5.969580347200829e-19

R91_105 V91 V105 2502.6891782735383
L91_105 V91 V105 4.857037026792641e-13
C91_105 V91 V105 1.1998667485390686e-18

R91_106 V91 V106 -1173.3719133559084
L91_106 V91 V106 -2.6883749989939543e-13
C91_106 V91 V106 -2.461310209579972e-18

R91_107 V91 V107 -3672.263325086475
L91_107 V91 V107 -8.367848775953361e-13
C91_107 V91 V107 -6.82923360828547e-19

R91_108 V91 V108 4269.420803206633
L91_108 V91 V108 1.0093013747411118e-12
C91_108 V91 V108 4.59737344034258e-19

R91_109 V91 V109 4943.059723466834
L91_109 V91 V109 1.1656459227244585e-12
C91_109 V91 V109 5.429012174284274e-19

R91_110 V91 V110 1114.7815583408278
L91_110 V91 V110 3.097043142598397e-13
C91_110 V91 V110 2.187072867635831e-18

R91_111 V91 V111 27316.10765193938
L91_111 V91 V111 1.0320678244352532e-12
C91_111 V91 V111 5.612186414475198e-19

R91_112 V91 V112 -6944.553131443082
L91_112 V91 V112 -6.233823391032772e-13
C91_112 V91 V112 -7.976792575284878e-19

R91_113 V91 V113 -12186.590020044656
L91_113 V91 V113 -8.807749657661956e-13
C91_113 V91 V113 -6.266971005619373e-19

R91_114 V91 V114 -2056.7948402327756
L91_114 V91 V114 -6.016441708887651e-13
C91_114 V91 V114 -1.1732345029577632e-18

R91_115 V91 V115 -18100.998065512493
L91_115 V91 V115 -1.4294796266685142e-12
C91_115 V91 V115 -3.416534573284824e-19

R91_116 V91 V116 16324.401292449886
L91_116 V91 V116 1.09846827080274e-12
C91_116 V91 V116 3.800132818861087e-19

R91_117 V91 V117 3501.276888616853
L91_117 V91 V117 9.542872254763167e-13
C91_117 V91 V117 5.887674651276977e-19

R91_118 V91 V118 2752.722615260876
L91_118 V91 V118 4.832602495385751e-13
C91_118 V91 V118 1.3133580409250984e-18

R91_119 V91 V119 2859.660569068052
L91_119 V91 V119 4.95607419314231e-13
C91_119 V91 V119 1.3351158578819763e-18

R91_120 V91 V120 1779.271397377854
L91_120 V91 V120 6.858064307805499e-11
C91_120 V91 V120 1.4430913574734925e-19

R91_121 V91 V121 -12613.085714697361
L91_121 V91 V121 -1.2269950829345042e-12
C91_121 V91 V121 -3.1511586580519354e-19

R91_122 V91 V122 1605.8343787255772
L91_122 V91 V122 -1.7211601898555725e-12
C91_122 V91 V122 -2.922960298317025e-20

R91_123 V91 V123 10046.71528280684
L91_123 V91 V123 2.3983226474063277e-12
C91_123 V91 V123 2.841768492188346e-19

R91_124 V91 V124 -9327.053218298517
L91_124 V91 V124 2.3713643151565384e-12
C91_124 V91 V124 1.8156946009758888e-19

R91_125 V91 V125 5733.289874717285
L91_125 V91 V125 1.9226110565475867e-12
C91_125 V91 V125 2.1507893956141805e-19

R91_126 V91 V126 -1098.9841357574653
L91_126 V91 V126 2.705919260159477e-12
C91_126 V91 V126 -1.684881423524032e-19

R91_127 V91 V127 1463.9265176130025
L91_127 V91 V127 -1.8839684010096095e-12
C91_127 V91 V127 -2.1451161347964218e-20

R91_128 V91 V128 6366.983906650828
L91_128 V91 V128 -8.532115185315673e-12
C91_128 V91 V128 1.486872937636372e-19

R91_129 V91 V129 8011.425987697545
L91_129 V91 V129 4.401492577428043e-11
C91_129 V91 V129 9.467120435522906e-20

R91_130 V91 V130 7853.611624226219
L91_130 V91 V130 3.156855296465354e-12
C91_130 V91 V130 3.2161702298664986e-19

R91_131 V91 V131 -9948.094527068566
L91_131 V91 V131 -4.8175532192637145e-12
C91_131 V91 V131 -8.51787235914318e-20

R91_132 V91 V132 -4917.206265160923
L91_132 V91 V132 -5.160940688624297e-12
C91_132 V91 V132 -1.9611910430482247e-19

R91_133 V91 V133 -3977.0695234804484
L91_133 V91 V133 -7.111751303004695e-13
C91_133 V91 V133 -9.580097804967117e-19

R91_134 V91 V134 -10019.066833158791
L91_134 V91 V134 6.582872297649062e-12
C91_134 V91 V134 1.4805792508629112e-19

R91_135 V91 V135 2085.2573410569894
L91_135 V91 V135 -4.161390598008733e-12
C91_135 V91 V135 -1.1026536135035983e-20

R91_136 V91 V136 15246.894871738376
L91_136 V91 V136 -1.4816291160398833e-11
C91_136 V91 V136 5.15378105933248e-20

R91_137 V91 V137 10235.896990647903
L91_137 V91 V137 1.8417127285305876e-12
C91_137 V91 V137 3.5613497140481705e-19

R91_138 V91 V138 -1678.6590493963326
L91_138 V91 V138 2.9214219627029147e-12
C91_138 V91 V138 -2.36964112487969e-20

R91_139 V91 V139 1218.460255811299
L91_139 V91 V139 -1.4521545479260173e-12
C91_139 V91 V139 -1.572960072160046e-19

R91_140 V91 V140 -6729.766248073532
L91_140 V91 V140 4.292148192081132e-12
C91_140 V91 V140 4.170401316525414e-20

R91_141 V91 V141 -4561.358494907837
L91_141 V91 V141 3.1787725950378215e-12
C91_141 V91 V141 5.157664275424734e-20

R91_142 V91 V142 36387.49165560569
L91_142 V91 V142 1.965408089496359e-12
C91_142 V91 V142 1.339153857714007e-19

R91_143 V91 V143 -4363.423007865603
L91_143 V91 V143 6.134228463175438e-12
C91_143 V91 V143 3.0997914693795636e-20

R91_144 V91 V144 13536.112248075922
L91_144 V91 V144 -3.921081260728689e-12
C91_144 V91 V144 -1.499284998468206e-19

R92_92 V92 0 -1470.532180685512
L92_92 V92 0 -2.0388635601262117e-13
C92_92 V92 0 -4.748371191758455e-19

R92_93 V92 V93 9352.941117309932
L92_93 V92 V93 2.171174422989024e-12
C92_93 V92 V93 2.0852255288517955e-19

R92_94 V92 V94 3383.66623080262
L92_94 V92 V94 6.884548268041374e-13
C92_94 V92 V94 9.240355347099664e-19

R92_95 V92 V95 -8732.362793859256
L92_95 V92 V95 -1.294604920931477e-12
C92_95 V92 V95 -4.936732929635815e-19

R92_96 V92 V96 -1870.9757210601722
L92_96 V92 V96 -3.51953977792008e-13
C92_96 V92 V96 -1.8953353743690435e-18

R92_97 V92 V97 13552.432050516767
L92_97 V92 V97 1.123419794701415e-12
C92_97 V92 V97 5.669067390200028e-19

R92_98 V92 V98 -2914.7121261257194
L92_98 V92 V98 -5.96228314815511e-13
C92_98 V92 V98 -9.611983757579048e-19

R92_99 V92 V99 19931.450656586374
L92_99 V92 V99 2.409507899280395e-12
C92_99 V92 V99 2.7661888451831346e-19

R92_100 V92 V100 5208.684610606293
L92_100 V92 V100 1.0546958617080854e-12
C92_100 V92 V100 7.2873771634408445e-19

R92_101 V92 V101 -3256.7848306397673
L92_101 V92 V101 -6.277927532976118e-13
C92_101 V92 V101 -1.0047623450981822e-18

R92_102 V92 V102 -3347.790779802746
L92_102 V92 V102 -7.877128020046112e-13
C92_102 V92 V102 -7.022202845432049e-19

R92_103 V92 V103 140121.08568516516
L92_103 V92 V103 2.9912968008048097e-12
C92_103 V92 V103 2.3857006592829137e-19

R92_104 V92 V104 -2154.608727218271
L92_104 V92 V104 -6.01830366854835e-13
C92_104 V92 V104 -1.2124260228568638e-18

R92_105 V92 V105 2143.427070748907
L92_105 V92 V105 5.250892018158938e-13
C92_105 V92 V105 1.2565404024697148e-18

R92_106 V92 V106 -1815.2999423184165
L92_106 V92 V106 -4.0539127900083733e-13
C92_106 V92 V106 -1.649661622679024e-18

R92_107 V92 V107 -5164.009672334936
L92_107 V92 V107 -9.382019363008663e-13
C92_107 V92 V107 -6.347242513338805e-19

R92_108 V92 V108 2386.0107558874756
L92_108 V92 V108 5.332579882287772e-13
C92_108 V92 V108 1.2868657228897972e-18

R92_109 V92 V109 -2734.064573265593
L92_109 V92 V109 -9.384792523523211e-13
C92_109 V92 V109 -8.881397908991326e-19

R92_110 V92 V110 2001.1388072474792
L92_110 V92 V110 4.462787368867691e-13
C92_110 V92 V110 1.4104901096190203e-18

R92_111 V92 V111 10363.306663654466
L92_111 V92 V111 9.913047696277997e-13
C92_111 V92 V111 6.732983825008604e-19

R92_112 V92 V112 -2702.999456181436
L92_112 V92 V112 -6.275131995721586e-13
C92_112 V92 V112 -9.120373206839138e-19

R92_113 V92 V113 8774.617617412176
L92_113 V92 V113 -3.823932284608425e-12
C92_113 V92 V113 1.1067118518443322e-20

R92_114 V92 V114 -2336.6704767902406
L92_114 V92 V114 -8.618206132026609e-13
C92_114 V92 V114 -8.470824758742482e-19

R92_115 V92 V115 -8207.631666347215
L92_115 V92 V115 -1.6530543853374962e-12
C92_115 V92 V115 -4.2054397524756287e-19

R92_116 V92 V116 4053.6092159979817
L92_116 V92 V116 7.018740937746697e-13
C92_116 V92 V116 8.551926685775828e-19

R92_117 V92 V117 8765.541625890084
L92_117 V92 V117 2.402017530831062e-12
C92_117 V92 V117 1.5779193487493845e-19

R92_118 V92 V118 8293.830535893938
L92_118 V92 V118 1.4147579568999597e-12
C92_118 V92 V118 3.7112028013227256e-19

R92_119 V92 V119 2769.976517447891
L92_119 V92 V119 5.52421966087355e-13
C92_119 V92 V119 1.2626190622590844e-18

R92_120 V92 V120 2464.379979653167
L92_120 V92 V120 1.2426371648204046e-12
C92_120 V92 V120 5.85115231064039e-19

R92_121 V92 V121 -5954.781108834666
L92_121 V92 V121 -2.888867772479867e-12
C92_121 V92 V121 -7.868186322196226e-20

R92_122 V92 V122 -83474.18062501345
L92_122 V92 V122 -3.2709825388708577e-12
C92_122 V92 V122 -5.526003320602079e-20

R92_123 V92 V123 -6605.4836992247465
L92_123 V92 V123 3.310512260532496e-12
C92_123 V92 V123 9.899152543611987e-20

R92_124 V92 V124 -26434.339832326074
L92_124 V92 V124 1.1410647159371542e-12
C92_124 V92 V124 6.563589429909802e-19

R92_125 V92 V125 5039.319233792833
L92_125 V92 V125 1.745891653673219e-12
C92_125 V92 V125 1.3184924632640176e-19

R92_126 V92 V126 -4514.152140398948
L92_126 V92 V126 2.867505817284027e-11
C92_126 V92 V126 -9.322322807783848e-20

R92_127 V92 V127 3827.0578798505626
L92_127 V92 V127 -8.723544757960949e-12
C92_127 V92 V127 1.0655959912646544e-19

R92_128 V92 V128 6875.162017202066
L92_128 V92 V128 3.3744919267587445e-10
C92_128 V92 V128 9.18167723442056e-21

R92_129 V92 V129 -9041.425857049197
L92_129 V92 V129 3.055586141386937e-12
C92_129 V92 V129 1.8157052047630863e-19

R92_130 V92 V130 2785.1351659001484
L92_130 V92 V130 4.843609814130091e-12
C92_130 V92 V130 2.488529201545368e-19

R92_131 V92 V131 6124.075751842724
L92_131 V92 V131 -2.7112258925936255e-12
C92_131 V92 V131 -1.817309477891236e-19

R92_132 V92 V132 68637.70337799483
L92_132 V92 V132 2.029555717876168e-12
C92_132 V92 V132 2.403751200703193e-19

R92_133 V92 V133 -13245.165399558025
L92_133 V92 V133 -1.1633664258608721e-12
C92_133 V92 V133 -5.474660583735208e-19

R92_134 V92 V134 -33477.73992212808
L92_134 V92 V134 1.152629229511329e-11
C92_134 V92 V134 3.505922776011317e-20

R92_135 V92 V135 5871.1080914113545
L92_135 V92 V135 2.0044260214639786e-10
C92_135 V92 V135 9.078728141322356e-20

R92_136 V92 V136 9650.423095269207
L92_136 V92 V136 1.4602919429325256e-10
C92_136 V92 V136 4.520473846858155e-20

R92_137 V92 V137 6597.2245947183665
L92_137 V92 V137 1.8928874620091016e-12
C92_137 V92 V137 3.549208682421792e-19

R92_138 V92 V138 12538.778317667919
L92_138 V92 V138 7.784112933255947e-12
C92_138 V92 V138 1.7108589401083237e-19

R92_139 V92 V139 3965.0924258420005
L92_139 V92 V139 -3.9094261498764585e-12
C92_139 V92 V139 -9.582392781699886e-20

R92_140 V92 V140 19971.043444601324
L92_140 V92 V140 2.3418366964077745e-12
C92_140 V92 V140 1.5343145937990447e-19

R92_141 V92 V141 -6820.023413712829
L92_141 V92 V141 6.434060861453085e-11
C92_141 V92 V141 -5.2290023468094e-20

R92_142 V92 V142 3576.2116025052624
L92_142 V92 V142 5.9321814028789875e-12
C92_142 V92 V142 2.1661371737684458e-19

R92_143 V92 V143 -138770.46158346088
L92_143 V92 V143 2.203343619271837e-11
C92_143 V92 V143 8.890211191079652e-20

R92_144 V92 V144 -31214.733445271024
L92_144 V92 V144 -2.314448975144993e-12
C92_144 V92 V144 -1.2790623443097944e-19

R93_93 V93 0 -136.5192766177001
L93_93 V93 0 6.717519659575181e-13
C93_93 V93 0 7.783780899396496e-19

R93_94 V93 V94 2211.1750665891013
L93_94 V93 V94 -5.755912183087304e-12
C93_94 V93 V94 5.496848934869636e-21

R93_95 V93 V95 3717.5828378448964
L93_95 V93 V95 4.637476775554221e-12
C93_95 V93 V95 7.503575135262809e-20

R93_96 V93 V96 4609.21665257858
L93_96 V93 V96 2.591833560119301e-12
C93_96 V93 V96 2.392762286915521e-19

R93_97 V93 V97 -1709.128158501776
L93_97 V93 V97 -6.97047513248284e-10
C93_97 V93 V97 -1.0507136416868192e-19

R93_98 V93 V98 -863.4098133240066
L93_98 V93 V98 3.3861683326629553e-12
C93_98 V93 V98 2.772969559059221e-20

R93_99 V93 V99 -188482.26515610993
L93_99 V93 V99 -5.878612107648816e-12
C93_99 V93 V99 -2.850378043532288e-20

R93_100 V93 V100 41851.98605134587
L93_100 V93 V100 -9.55919445447357e-12
C93_100 V93 V100 -7.078656165647583e-20

R93_101 V93 V101 -8250.161332218098
L93_101 V93 V101 1.9612165796341694e-11
C93_101 V93 V101 -2.6440355709356423e-19

R93_102 V93 V102 -10669.459832636323
L93_102 V93 V102 1.5388157832577892e-12
C93_102 V93 V102 9.750906135026882e-20

R93_103 V93 V103 -3080.7111979663127
L93_103 V93 V103 -2.9515418886510453e-12
C93_103 V93 V103 -2.841879902275837e-19

R93_104 V93 V104 3374.5457018560455
L93_104 V93 V104 7.169796380173963e-12
C93_104 V93 V104 6.346255217057299e-20

R93_105 V93 V105 17930.72222834963
L93_105 V93 V105 -2.0781115160531293e-12
C93_105 V93 V105 -2.540366943293424e-19

R93_106 V93 V106 1161.6685515502254
L93_106 V93 V106 1.2411117159372274e-12
C93_106 V93 V106 3.4998298124521147e-19

R93_107 V93 V107 -5941.355691502282
L93_107 V93 V107 1.542779656504192e-12
C93_107 V93 V107 3.985610954498174e-19

R93_108 V93 V108 -1382.605210971943
L93_108 V93 V108 -2.1621564707496913e-12
C93_108 V93 V108 2.4961103613076125e-21

R93_109 V93 V109 -1971.9406328874793
L93_109 V93 V109 -2.8432147258581064e-11
C93_109 V93 V109 1.0161552680415684e-19

R93_110 V93 V110 -42592.943058925826
L93_110 V93 V110 -2.2705436159702882e-12
C93_110 V93 V110 -1.9030824449398212e-19

R93_111 V93 V111 -1160.2378014701555
L93_111 V93 V111 -2.046232054488217e-12
C93_111 V93 V111 -2.8018232505525385e-19

R93_112 V93 V112 -751.0619538339564
L93_112 V93 V112 2.443407736027597e-12
C93_112 V93 V112 -5.832936658878508e-20

R93_113 V93 V113 -1749.7129413586683
L93_113 V93 V113 7.1147393743481284e-12
C93_113 V93 V113 -1.482998518570085e-20

R93_114 V93 V114 6165.46538217616
L93_114 V93 V114 2.282427930755373e-12
C93_114 V93 V114 8.473124732786069e-20

R93_115 V93 V115 3946.3146518917124
L93_115 V93 V115 3.2038033926105158e-12
C93_115 V93 V115 1.840954699908315e-19

R93_116 V93 V116 22329.177170338553
L93_116 V93 V116 -2.108280234272646e-12
C93_116 V93 V116 -8.215799793473849e-20

R93_117 V93 V117 7311.257821987407
L93_117 V93 V117 -8.06266043295958e-12
C93_117 V93 V117 5.608359187192236e-20

R93_118 V93 V118 2869.673924154412
L93_118 V93 V118 -2.754449702011519e-12
C93_118 V93 V118 -1.410558659645501e-19

R93_119 V93 V119 -1148.4351610511542
L93_119 V93 V119 -1.783955957673812e-12
C93_119 V93 V119 -2.1104806022059234e-19

R93_120 V93 V120 880.646190505688
L93_120 V93 V120 5.290788364463089e-12
C93_120 V93 V120 -3.358301772022182e-20

R93_121 V93 V121 -431.13240642198735
L93_121 V93 V121 5.716699457441544e-12
C93_121 V93 V121 1.1577377550400413e-19

R93_122 V93 V122 -428.7223062270375
L93_122 V93 V122 3.602051418839855e-12
C93_122 V93 V122 -7.702328846838873e-20

R93_123 V93 V123 -3233.578901626779
L93_123 V93 V123 6.7190739560074224e-12
C93_123 V93 V123 -3.635369593094267e-20

R93_124 V93 V124 -4154.599541780143
L93_124 V93 V124 -2.268511747360971e-11
C93_124 V93 V124 -9.838983540629633e-20

R93_125 V93 V125 381.3451595022762
L93_125 V93 V125 -1.3554970660707463e-11
C93_125 V93 V125 -9.414966210809215e-20

R93_126 V93 V126 1000.6184822454693
L93_126 V93 V126 -2.147876660253551e-12
C93_126 V93 V126 -9.309728609705028e-21

R93_127 V93 V127 -9105.617019401787
L93_127 V93 V127 2.8764452401411594e-12
C93_127 V93 V127 -2.854960620324779e-21

R93_128 V93 V128 -11732.743623761306
L93_128 V93 V128 -1.0649618789614412e-10
C93_128 V93 V128 8.664437241801257e-22

R93_129 V93 V129 27306.677605721463
L93_129 V93 V129 3.1603874887261282e-12
C93_129 V93 V129 8.815169249589729e-20

R93_130 V93 V130 -35596.1341427635
L93_130 V93 V130 -2.1917308056196236e-12
C93_130 V93 V130 -1.9731387809125832e-20

R93_131 V93 V131 2533.898220110244
L93_131 V93 V131 -6.240656988866677e-12
C93_131 V93 V131 5.953775593767105e-20

R93_132 V93 V132 3839.364151911137
L93_132 V93 V132 -9.476362979273503e-12
C93_132 V93 V132 9.873703562931852e-21

R93_133 V93 V133 1455.21849996411
L93_133 V93 V133 5.703422605021776e-12
C93_133 V93 V133 7.214908086944576e-20

R93_134 V93 V134 1881.5503365489903
L93_134 V93 V134 -2.1504765062886682e-11
C93_134 V93 V134 -9.151671407901666e-20

R93_135 V93 V135 -4474.690693232828
L93_135 V93 V135 4.714879749793935e-12
C93_135 V93 V135 -3.3879649392751116e-20

R93_136 V93 V136 8767.34873021015
L93_136 V93 V136 -1.4436203937980804e-10
C93_136 V93 V136 2.9916280526749015e-22

R93_137 V93 V137 683.0592920200357
L93_137 V93 V137 9.137234950985143e-12
C93_137 V93 V137 5.254723934556985e-20

R93_138 V93 V138 917.5206183165096
L93_138 V93 V138 -2.189017422863527e-12
C93_138 V93 V138 8.337092297191806e-21

R93_139 V93 V139 -10110.180714390799
L93_139 V93 V139 2.0142071602678282e-12
C93_139 V93 V139 6.016673441145668e-20

R93_140 V93 V140 1862.0017333400965
L93_140 V93 V140 -3.784431982084474e-12
C93_140 V93 V140 1.4146599138307647e-20

R93_141 V93 V141 2300.9945252020375
L93_141 V93 V141 -1.879613741210846e-11
C93_141 V93 V141 5.597557648232704e-21

R93_142 V93 V142 13278.251065803106
L93_142 V93 V142 -2.670447055865228e-12
C93_142 V93 V142 -7.110139019121889e-21

R93_143 V93 V143 -4094.967736122417
L93_143 V93 V143 -3.2139140124314432e-12
C93_143 V93 V143 -6.749160957479078e-20

R93_144 V93 V144 -2037.5312489511584
L93_144 V93 V144 2.6264012165765803e-11
C93_144 V93 V144 -6.3890212786786e-20

R94_94 V94 0 611.6082363490672
L94_94 V94 0 2.86055908068085e-13
C94_94 V94 0 3.8791620384561277e-19

R94_95 V94 V95 10960.254214287454
L94_95 V94 V95 1.5603531495236035e-12
C94_95 V94 V95 4.36754764756208e-19

R94_96 V94 V96 4113.724698998987
L94_96 V94 V96 9.087924084813532e-13
C94_96 V94 V96 7.924971961586081e-19

R94_97 V94 V97 -1548.4685400651906
L94_97 V94 V97 -2.1384964154129207e-12
C94_97 V94 V97 -5.109840443405619e-19

R94_98 V94 V98 -1446.9237870898992
L94_98 V94 V98 7.31831990554917e-13
C94_98 V94 V98 5.186746411256617e-19

R94_99 V94 V99 1474.8945899987418
L94_99 V94 V99 -9.585873187569487e-12
C94_99 V94 V99 -1.3022873918289252e-19

R94_100 V94 V100 -31583.79547630566
L94_100 V94 V100 -1.9050801997129707e-12
C94_100 V94 V100 -3.9761895681695563e-19

R94_101 V94 V101 2051.015303134459
L94_101 V94 V101 7.138187475057827e-13
C94_101 V94 V101 6.9648252227704445e-19

R94_102 V94 V102 -2863.231583414859
L94_102 V94 V102 1.920875535939423e-12
C94_102 V94 V102 -1.7554317291082645e-19

R94_103 V94 V103 -54963.9488604602
L94_103 V94 V103 1.9348710370455774e-12
C94_103 V94 V103 4.564017068774862e-19

R94_104 V94 V104 2232.761346211227
L94_104 V94 V104 1.7096567843620863e-12
C94_104 V94 V104 4.81370280637986e-19

R94_105 V94 V105 -152555.69617146943
L94_105 V94 V105 -8.985030695535172e-13
C94_105 V94 V105 -6.422832271120116e-19

R94_106 V94 V106 1225.1913776875915
L94_106 V94 V106 7.610787567506224e-13
C94_106 V94 V106 8.2419040868005475e-19

R94_107 V94 V107 -12867.016073606828
L94_107 V94 V107 5.169612390184889e-12
C94_107 V94 V107 -2.1936631742468654e-19

R94_108 V94 V108 -1130.9053005404617
L94_108 V94 V108 -1.2111821643474089e-12
C94_108 V94 V108 -3.3731894601191724e-19

R94_109 V94 V109 -10718.073433313182
L94_109 V94 V109 1.7951168219709186e-12
C94_109 V94 V109 5.158152174528145e-19

R94_110 V94 V110 -800.1430819697733
L94_110 V94 V110 -5.356454444696874e-13
C94_110 V94 V110 -1.0057627671181268e-18

R94_111 V94 V111 2806.149093383196
L94_111 V94 V111 -2.343496794531095e-11
C94_111 V94 V111 -1.556852783401397e-19

R94_112 V94 V112 -853.6143067413184
L94_112 V94 V112 8.411849388008345e-13
C94_112 V94 V112 2.1463022261825974e-19

R94_113 V94 V113 -1296.66050886387
L94_113 V94 V113 2.6752565365391038e-12
C94_113 V94 V113 -3.841326416926652e-20

R94_114 V94 V114 -29035.99368429476
L94_114 V94 V114 1.1875672712398607e-12
C94_114 V94 V114 5.513557754553571e-19

R94_115 V94 V115 -2423.7271862873354
L94_115 V94 V115 -6.124389112305782e-10
C94_115 V94 V115 -1.257326713296547e-19

R94_116 V94 V116 3778.3277836179877
L94_116 V94 V116 -1.3129747958287884e-12
C94_116 V94 V116 -2.6898115945817373e-19

R94_117 V94 V117 -1975.2650062979312
L94_117 V94 V117 -1.9236431844159216e-12
C94_117 V94 V117 -1.1552049601434695e-20

R94_118 V94 V118 2877.793303051762
L94_118 V94 V118 -1.4479849306165675e-12
C94_118 V94 V118 -2.7771156119070637e-19

R94_119 V94 V119 -36046.513534275604
L94_119 V94 V119 -1.2391949610324836e-12
C94_119 V94 V119 -6.648541708565651e-19

R94_120 V94 V120 -449.87761552544794
L94_120 V94 V120 -9.723178311981867e-13
C94_120 V94 V120 -2.145861656825562e-19

R94_121 V94 V121 -792.4126058982476
L94_121 V94 V121 1.1575773128819667e-12
C94_121 V94 V121 6.150469277810298e-20

R94_122 V94 V122 -217.04571584834883
L94_122 V94 V122 2.0792501256295112e-12
C94_122 V94 V122 3.4924458575942345e-20

R94_123 V94 V123 -1154.9418367123067
L94_123 V94 V123 -5.6315822315063165e-12
C94_123 V94 V123 -1.1134007348237946e-19

R94_124 V94 V124 21587.68679997926
L94_124 V94 V124 -3.4738715573397453e-12
C94_124 V94 V124 -3.0087359260763726e-19

R94_125 V94 V125 2010.137991086505
L94_125 V94 V125 -8.623627623310436e-13
C94_125 V94 V125 -8.459736643142111e-20

R94_126 V94 V126 194.6729229482489
L94_126 V94 V126 6.677578396386816e-12
C94_126 V94 V126 -5.841954166166356e-20

R94_127 V94 V127 -274.83715596461303
L94_127 V94 V127 -3.0257908517641915e-12
C94_127 V94 V127 -4.6687380067185923e-20

R94_128 V94 V128 -2743.6970597219592
L94_128 V94 V128 -1.3193496496794755e-11
C94_128 V94 V128 -7.15568845277457e-20

R94_129 V94 V129 -728.4351184425784
L94_129 V94 V129 -3.0954208768407554e-12
C94_129 V94 V129 -1.2502397436853973e-19

R94_130 V94 V130 1138.0181350361388
L94_130 V94 V130 -1.3241412260367249e-11
C94_130 V94 V130 -2.6983184278229547e-20

R94_131 V94 V131 775.4592217114116
L94_131 V94 V131 -1.3554510323378377e-10
C94_131 V94 V131 -8.221385521698281e-20

R94_132 V94 V132 1039.6229752540537
L94_132 V94 V132 -4.4584997062966126e-12
C94_132 V94 V132 -1.280410645729144e-19

R94_133 V94 V133 1653.5643379950748
L94_133 V94 V133 3.5919166436159763e-12
C94_133 V94 V133 2.3789442212622033e-19

R94_134 V94 V134 1114.3357699443836
L94_134 V94 V134 -2.222764958423136e-11
C94_134 V94 V134 -1.4022071103703444e-20

R94_135 V94 V135 -395.84368371096053
L94_135 V94 V135 -3.576099264575665e-12
C94_135 V94 V135 -2.3801180794882828e-20

R94_136 V94 V136 -298004.9518460331
L94_136 V94 V136 4.9373824652925365e-11
C94_136 V94 V136 3.4739000473140073e-20

R94_137 V94 V137 2358.5765075212785
L94_137 V94 V137 -1.3358201914455305e-12
C94_137 V94 V137 -1.8059933845319755e-19

R94_138 V94 V138 227.5199945097984
L94_138 V94 V138 1.4531716713183128e-11
C94_138 V94 V138 -1.9555985730006173e-20

R94_139 V94 V139 -215.23181986871964
L94_139 V94 V139 -2.336158588803928e-12
C94_139 V94 V139 -1.480536695775388e-20

R94_140 V94 V140 736.0214740605517
L94_140 V94 V140 -7.794365404549418e-12
C94_140 V94 V140 1.7971665863293156e-20

R94_141 V94 V141 924.1183615153285
L94_141 V94 V141 1.782990457077674e-10
C94_141 V94 V141 4.6252922167542795e-20

R94_142 V94 V142 875.4608106731968
L94_142 V94 V142 -5.384692231856503e-12
C94_142 V94 V142 -1.3464691481443338e-19

R94_143 V94 V143 723.9226257689764
L94_143 V94 V143 6.794313846253267e-12
C94_143 V94 V143 -7.75968494931235e-20

R94_144 V94 V144 -1230.651068914517
L94_144 V94 V144 4.40234538026055e-12
C94_144 V94 V144 2.508912603058283e-20

R95_95 V95 0 -563.2024048209897
L95_95 V95 0 -6.272422160510473e-13
C95_95 V95 0 5.868284828538877e-21

R95_96 V95 V96 -235179.00074589698
L95_96 V95 V96 -5.4342707468777495e-12
C95_96 V95 V96 -1.6944932741929252e-19

R95_97 V95 V97 19295.24827326974
L95_97 V95 V97 1.7022992223536352e-12
C95_97 V95 V97 2.8937238916424093e-19

R95_98 V95 V98 -2704.869789488462
L95_98 V95 V98 -1.3245890732750754e-12
C95_98 V95 V98 -5.440881007510047e-19

R95_99 V95 V99 -5317.399259433211
L95_99 V95 V99 6.819237504461082e-12
C95_99 V95 V99 8.425160741482453e-20

R95_100 V95 V100 32363.728972030854
L95_100 V95 V100 5.579405941196964e-12
C95_100 V95 V100 8.237040772378237e-20

R95_101 V95 V101 -4207.057224153573
L95_101 V95 V101 -1.2238883568190342e-12
C95_101 V95 V101 -6.104235486457661e-19

R95_102 V95 V102 -7245.793518651751
L95_102 V95 V102 -1.1695597216636683e-12
C95_102 V95 V102 -5.530169638233825e-19

R95_103 V95 V103 21403.24559265422
L95_103 V95 V103 1.3660528186891713e-11
C95_103 V95 V103 9.665432813836678e-21

R95_104 V95 V104 10684.343731317727
L95_104 V95 V104 3.0339390990226e-12
C95_104 V95 V104 1.731958420896197e-19

R95_105 V95 V105 5112.765470911929
L95_105 V95 V105 8.324455121018948e-13
C95_105 V95 V105 7.458874301283369e-19

R95_106 V95 V106 -3340.772764055706
L95_106 V95 V106 -4.938554122309572e-13
C95_106 V95 V106 -1.3659001822294847e-18

R95_107 V95 V107 -3019.045027610156
L95_107 V95 V107 -1.4474191133201023e-12
C95_107 V95 V107 -4.463374224908728e-19

R95_108 V95 V108 16684.50836657364
L95_108 V95 V108 1.543748544988789e-12
C95_108 V95 V108 4.1972535187984446e-19

R95_109 V95 V109 -19417.763697752926
L95_109 V95 V109 2.614220256427796e-12
C95_109 V95 V109 2.373062094243822e-19

R95_110 V95 V110 1408.6687840241116
L95_110 V95 V110 5.510747104335419e-13
C95_110 V95 V110 1.2750234272818735e-18

R95_111 V95 V111 -3290.88627936742
L95_111 V95 V111 1.3774789535626337e-12
C95_111 V95 V111 3.89676380004836e-19

R95_112 V95 V112 -3273.3683359649435
L95_112 V95 V112 -1.2906603397586345e-12
C95_112 V95 V112 -5.511621876419173e-19

R95_113 V95 V113 -5294.418922898431
L95_113 V95 V113 -2.0403012809305607e-12
C95_113 V95 V113 -3.2264494147281073e-19

R95_114 V95 V114 -25542.4468224239
L95_114 V95 V114 -1.186037681068824e-12
C95_114 V95 V114 -7.332347294060186e-19

R95_115 V95 V115 9041.982706684728
L95_115 V95 V115 -2.6015441171585e-12
C95_115 V95 V115 -2.094321792098515e-19

R95_116 V95 V116 -47445.18740812942
L95_116 V95 V116 1.919204640536252e-12
C95_116 V95 V116 2.9229411801014374e-19

R95_117 V95 V117 2862.3927473393987
L95_117 V95 V117 2.4602427067324327e-12
C95_117 V95 V117 2.979354170835855e-19

R95_118 V95 V118 4039.4486291183
L95_118 V95 V118 1.0189574128234788e-12
C95_118 V95 V118 6.683330733134531e-19

R95_119 V95 V119 -4389.15359086337
L95_119 V95 V119 8.89648290097812e-13
C95_119 V95 V119 7.4945865280448085e-19

R95_120 V95 V120 807.2310236142234
L95_120 V95 V120 -1.4767366508396148e-11
C95_120 V95 V120 1.4071552451069564e-19

R95_121 V95 V121 -1505.6103917541104
L95_121 V95 V121 -4.917109800345435e-12
C95_121 V95 V121 -1.5924949867693184e-19

R95_122 V95 V122 2111.32262871821
L95_122 V95 V122 -3.131287793185915e-11
C95_122 V95 V122 -7.856118867159703e-21

R95_123 V95 V123 4042.3683833377636
L95_123 V95 V123 2.442683222193534e-12
C95_123 V95 V123 1.5883793224804842e-19

R95_124 V95 V124 16316.194071188835
L95_124 V95 V124 2.76606244439593e-12
C95_124 V95 V124 1.501786827434621e-19

R95_125 V95 V125 976.8912214012569
L95_125 V95 V125 1.671615665492256e-11
C95_125 V95 V125 1.0005860325529938e-19

R95_126 V95 V126 -804.8485956618949
L95_126 V95 V126 9.070682380790248e-12
C95_126 V95 V126 -9.104714643737837e-20

R95_127 V95 V127 907.234928554642
L95_127 V95 V127 -3.386998421185858e-12
C95_127 V95 V127 1.4705336112344345e-20

R95_128 V95 V128 -29588.785779545455
L95_128 V95 V128 -1.7138329023000132e-10
C95_128 V95 V128 8.363361650716979e-20

R95_129 V95 V129 1791.3119832452442
L95_129 V95 V129 5.436515644875292e-12
C95_129 V95 V129 1.005995975948803e-19

R95_130 V95 V130 -2634.7361985268763
L95_130 V95 V130 -1.7877814654360965e-11
C95_130 V95 V130 1.7732481390105658e-19

R95_131 V95 V131 -2493.485855743606
L95_131 V95 V131 -2.437724739495198e-12
C95_131 V95 V131 -1.3145511170927398e-19

R95_132 V95 V132 -4093.246149798731
L95_132 V95 V132 -2.5758508055898205e-11
C95_132 V95 V132 -4.6330944533231383e-20

R95_133 V95 V133 -15915.727335918053
L95_133 V95 V133 -1.3303823736809708e-12
C95_133 V95 V133 -4.537037729706596e-19

R95_134 V95 V134 -23171.09226501039
L95_134 V95 V134 5.1342906661113646e-11
C95_134 V95 V134 2.4013519670140802e-20

R95_135 V95 V135 1380.3414000402695
L95_135 V95 V135 -1.027944746074949e-11
C95_135 V95 V135 2.8335877286824324e-20

R95_136 V95 V136 -55935.531091731864
L95_136 V95 V136 -3.488282963410238e-11
C95_136 V95 V136 2.8460939739351683e-20

R95_137 V95 V137 1723.382217920299
L95_137 V95 V137 4.7187834192422015e-12
C95_137 V95 V137 2.174524635050953e-19

R95_138 V95 V138 -1023.4413588417453
L95_138 V95 V138 3.053864826378784e-11
C95_138 V95 V138 6.503462633366926e-20

R95_139 V95 V139 718.5199216919443
L95_139 V95 V139 -2.36072776985035e-12
C95_139 V95 V139 -9.552586668931661e-20

R95_140 V95 V140 -3310.6199230467805
L95_140 V95 V140 2.1706746897485492e-11
C95_140 V95 V140 2.179905606649223e-20

R95_141 V95 V141 -50726.712902674844
L95_141 V95 V141 6.94971572836187e-12
C95_141 V95 V141 3.4268322175380456e-20

R95_142 V95 V142 -2292.764230200003
L95_142 V95 V142 5.72766778751477e-12
C95_142 V95 V142 1.5083315762499023e-19

R95_143 V95 V143 -1724.1153571964314
L95_143 V95 V143 2.2105645676008565e-11
C95_143 V95 V143 2.82233413632293e-21

R95_144 V95 V144 17794.336620580314
L95_144 V95 V144 -6.9559401190549536e-12
C95_144 V95 V144 -8.148472524330835e-20

R96_96 V96 0 4402.410960042257
L96_96 V96 0 -2.4347997214599725e-13
C96_96 V96 0 -7.979924501859927e-19

R96_97 V96 V97 4903.897638484367
L96_97 V96 V97 1.0713096949182892e-12
C96_97 V96 V97 5.3324995169709655e-19

R96_98 V96 V98 -3398.494619030574
L96_98 V96 V98 -9.429533277165211e-13
C96_98 V96 V98 -7.566574597427517e-19

R96_99 V96 V99 77854.58066902183
L96_99 V96 V99 2.352240979790787e-12
C96_99 V96 V99 2.726741276559386e-19

R96_100 V96 V100 4361.111352587258
L96_100 V96 V100 8.450017689539389e-13
C96_100 V96 V100 8.382907616738881e-19

R96_101 V96 V101 -4049.927902726041
L96_101 V96 V101 -9.251175437016636e-13
C96_101 V96 V101 -7.485474751253948e-19

R96_102 V96 V102 -23422.06973044103
L96_102 V96 V102 -1.3844045539697925e-12
C96_102 V96 V102 -4.284397212515201e-19

R96_103 V96 V103 5842.839501083844
L96_103 V96 V103 1.5248832281400003e-12
C96_103 V96 V103 3.3478625377328783e-19

R96_104 V96 V104 -2326.277594406246
L96_104 V96 V104 -4.5033376711939534e-13
C96_104 V96 V104 -1.504451733773863e-18

R96_105 V96 V105 3657.5559805702374
L96_105 V96 V105 6.999835271805548e-13
C96_105 V96 V105 1.0663125185428615e-18

R96_106 V96 V106 -3446.551644867422
L96_106 V96 V106 -6.289380749360379e-13
C96_106 V96 V106 -1.1279668012143092e-18

R96_107 V96 V107 -4160.996968160206
L96_107 V96 V107 -1.1771065554076608e-12
C96_107 V96 V107 -4.846483747528038e-19

R96_108 V96 V108 3434.0741806119795
L96_108 V96 V108 5.838229285420463e-13
C96_108 V96 V108 1.1458219581250248e-18

R96_109 V96 V109 -2492.5384601685596
L96_109 V96 V109 -7.016844226180263e-13
C96_109 V96 V109 -1.1982796539529029e-18

R96_110 V96 V110 2438.6134618674896
L96_110 V96 V110 8.061998849459459e-13
C96_110 V96 V110 8.824905441214098e-19

R96_111 V96 V111 30642.76514482097
L96_111 V96 V111 1.0039830283212094e-12
C96_111 V96 V111 5.847795498129217e-19

R96_112 V96 V112 -3251.1820305245956
L96_112 V96 V112 -1.2360751934471895e-12
C96_112 V96 V112 -6.97172924369993e-19

R96_113 V96 V113 18757.930990068624
L96_113 V96 V113 3.104102192258234e-11
C96_113 V96 V113 2.3212388175561927e-19

R96_114 V96 V114 13026.844583433221
L96_114 V96 V114 -1.5565001605152948e-12
C96_114 V96 V114 -5.694342908448781e-19

R96_115 V96 V115 188899.31323067425
L96_115 V96 V115 -1.9710917361039498e-12
C96_115 V96 V115 -3.4970724167596003e-19

R96_116 V96 V116 4295.156014247214
L96_116 V96 V116 8.716195352302515e-13
C96_116 V96 V116 7.425704119611579e-19

R96_117 V96 V117 39239.29434161336
L96_117 V96 V117 -1.9409756579071414e-10
C96_117 V96 V117 -6.847582069912063e-20

R96_118 V96 V118 -15732.239474852278
L96_118 V96 V118 7.926931792010159e-11
C96_118 V96 V118 1.9135052847409147e-20

R96_119 V96 V119 13683.119313447844
L96_119 V96 V119 7.602780839745193e-13
C96_119 V96 V119 9.468044930537594e-19

R96_120 V96 V120 1547.8811937607065
L96_120 V96 V120 1.7297657555437848e-12
C96_120 V96 V120 5.552362857492785e-19

R96_121 V96 V121 -3558.9813945233595
L96_121 V96 V121 3.986096120048486e-12
C96_121 V96 V121 -3.480092353498058e-20

R96_122 V96 V122 4838.855951397696
L96_122 V96 V122 5.494235970997285e-12
C96_122 V96 V122 -5.827248729161159e-20

R96_123 V96 V123 3173.921385445495
L96_123 V96 V123 6.2446371730993505e-12
C96_123 V96 V123 -1.215377511947721e-20

R96_124 V96 V124 5284.258828066985
L96_124 V96 V124 9.592560740454342e-13
C96_124 V96 V124 6.12718006069417e-19

R96_125 V96 V125 1957.7086140018323
L96_125 V96 V125 -1.6509404201458473e-11
C96_125 V96 V125 6.46394076277409e-20

R96_126 V96 V126 -2154.2916547177538
L96_126 V96 V126 -4.882970196770055e-12
C96_126 V96 V126 -7.089986847438621e-20

R96_127 V96 V127 2429.5697203044556
L96_127 V96 V127 8.534394121186256e-11
C96_127 V96 V127 1.1615435779092047e-19

R96_128 V96 V128 6406.3838592158245
L96_128 V96 V128 -3.718556519043152e-12
C96_128 V96 V128 -2.3869135921321287e-20

R96_129 V96 V129 2228.6278766005
L96_129 V96 V129 2.789893304179703e-12
C96_129 V96 V129 1.4126993578384722e-19

R96_130 V96 V130 -3387.499289106217
L96_130 V96 V130 6.568858013893222e-11
C96_130 V96 V130 1.8337702287314115e-19

R96_131 V96 V131 -2627.808724862357
L96_131 V96 V131 -1.900120843294025e-12
C96_131 V96 V131 -1.7301648702300993e-19

R96_132 V96 V132 10201.52962036901
L96_132 V96 V132 1.6955204546452414e-12
C96_132 V96 V132 2.9337529560919483e-19

R96_133 V96 V133 -10327.030182917248
L96_133 V96 V133 -1.531672304127076e-12
C96_133 V96 V133 -3.518090458314899e-19

R96_134 V96 V134 -43796.596036723226
L96_134 V96 V134 -7.649480722635247e-11
C96_134 V96 V134 5.83072276992055e-21

R96_135 V96 V135 3399.5317698345366
L96_135 V96 V135 1.5066710625228957e-11
C96_135 V96 V135 9.069703848266829e-20

R96_136 V96 V136 126950.91908176418
L96_136 V96 V136 -4.150980080734661e-12
C96_136 V96 V136 -8.685234155829995e-21

R96_137 V96 V137 2769.299200138521
L96_137 V96 V137 6.920128298846574e-12
C96_137 V96 V137 2.8518135552326015e-19

R96_138 V96 V138 -1979.3381820811128
L96_138 V96 V138 -5.1682004476060836e-12
C96_138 V96 V138 1.479029216524654e-19

R96_139 V96 V139 2103.6526780670024
L96_139 V96 V139 -5.432827716899511e-12
C96_139 V96 V139 -1.008818729716084e-19

R96_140 V96 V140 -667886.3987955948
L96_140 V96 V140 6.160837479930359e-12
C96_140 V96 V140 1.2925377943717014e-19

R96_141 V96 V141 -11672.70671004004
L96_141 V96 V141 -4.5405805727857414e-11
C96_141 V96 V141 -9.267605032700418e-20

R96_142 V96 V142 -2898.026045083017
L96_142 V96 V142 -1.056662711037572e-11
C96_142 V96 V142 1.6132270101611848e-19

R96_143 V96 V143 -4062.6983758840647
L96_143 V96 V143 4.0865090591963457e-10
C96_143 V96 V143 6.80482020786164e-20

R96_144 V96 V144 -29608.03476231025
L96_144 V96 V144 -3.727226158144864e-12
C96_144 V96 V144 -7.0292864036674e-20

R97_97 V97 0 -222.08706488893566
L97_97 V97 0 -2.031991004752686e-12
C97_97 V97 0 -1.9427726251860813e-19

R97_98 V97 V98 1434.8236564901945
L97_98 V97 V98 -2.7098511981951118e-12
C97_98 V97 V98 2.2755707926617587e-19

R97_99 V97 V99 -2715.352799750844
L97_99 V97 V99 4.379988561433499e-12
C97_99 V97 V99 -5.0325547228932475e-20

R97_100 V97 V100 -4672.62090789787
L97_100 V97 V100 -1.8149874758810625e-12
C97_100 V97 V100 -3.231339323490857e-19

R97_101 V97 V101 -14816.675920249327
L97_101 V97 V101 1.2280371590089796e-11
C97_101 V97 V101 2.325666774229926e-19

R97_102 V97 V102 -3002.0508501907498
L97_102 V97 V102 -5.427009861468354e-13
C97_102 V97 V102 -6.94403199384911e-19

R97_103 V97 V103 5852.5681198347
L97_103 V97 V103 1.391731501856576e-12
C97_103 V97 V103 5.093043959940611e-19

R97_104 V97 V104 -4434.501922278093
L97_104 V97 V104 2.647719983586299e-12
C97_104 V97 V104 2.1765582271667024e-19

R97_105 V97 V105 -26212.495189664267
L97_105 V97 V105 -3.856584319388551e-12
C97_105 V97 V105 -3.3825340634456993e-19

R97_106 V97 V106 -2148.3823622809327
L97_106 V97 V106 1.4210792963486233e-12
C97_106 V97 V106 3.5872424873998144e-19

R97_107 V97 V107 -9602.627378289939
L97_107 V97 V107 -9.12357336014899e-13
C97_107 V97 V107 -4.815755262953614e-19

R97_108 V97 V108 1285.3177118957478
L97_108 V97 V108 1.3191145311293718e-12
C97_108 V97 V108 3.3489198308314607e-19

R97_109 V97 V109 2355.903430746197
L97_109 V97 V109 1.2917561716965817e-12
C97_109 V97 V109 5.524596268599951e-19

R97_110 V97 V110 3065.8470494944427
L97_110 V97 V110 -1.305506290010502e-12
C97_110 V97 V110 -4.520498117755447e-19

R97_111 V97 V111 24538.395765192192
L97_111 V97 V111 -7.163460451340427e-12
C97_111 V97 V111 4.235737791805222e-22

R97_112 V97 V112 1292.3698161101688
L97_112 V97 V112 -6.910654928484863e-13
C97_112 V97 V112 -1.696207632351572e-19

R97_113 V97 V113 1485.5219318639602
L97_113 V97 V113 -1.6152752837494598e-12
C97_113 V97 V113 -1.7826736521934802e-19

R97_114 V97 V114 -4116.942378702525
L97_114 V97 V114 -1.2176951231504401e-11
C97_114 V97 V114 3.1548663678563523e-19

R97_115 V97 V115 -9157.185216700991
L97_115 V97 V115 -1.7139560472395693e-12
C97_115 V97 V115 -2.6889928066523276e-19

R97_116 V97 V116 -12839.158432261202
L97_116 V97 V116 1.660294183437253e-12
C97_116 V97 V116 1.5365237472213722e-19

R97_117 V97 V117 3701.5414484175412
L97_117 V97 V117 1.8544570452377533e-12
C97_117 V97 V117 2.7699614728642116e-19

R97_118 V97 V118 -3474.8627097858875
L97_118 V97 V118 4.072003058557661e-12
C97_118 V97 V118 -7.108811586021484e-20

R97_119 V97 V119 3401.161049826641
L97_119 V97 V119 -2.1435000997910387e-12
C97_119 V97 V119 -3.487882237045258e-19

R97_120 V97 V120 1731.6819839323655
L97_120 V97 V120 -3.947567561818232e-12
C97_120 V97 V120 -7.279282532081854e-20

R97_121 V97 V121 764.9317176417954
L97_121 V97 V121 -1.1165024118002815e-12
C97_121 V97 V121 7.446797891189452e-20

R97_122 V97 V122 366.720243590932
L97_122 V97 V122 -4.733039856115913e-13
C97_122 V97 V122 2.4262823508659813e-20

R97_123 V97 V123 11768.305434415703
L97_123 V97 V123 -1.1748945086685857e-12
C97_123 V97 V123 -5.439139316869264e-20

R97_124 V97 V124 -1967.266735214215
L97_124 V97 V124 -1.827475833937654e-12
C97_124 V97 V124 -1.6570767636752595e-19

R97_125 V97 V125 -872.7312499760757
L97_125 V97 V125 1.057322420961591e-12
C97_125 V97 V125 4.6748529786369894e-20

R97_126 V97 V126 -380.42960676584266
L97_126 V97 V126 5.767350609414109e-13
C97_126 V97 V126 -1.8057668834543228e-20

R97_127 V97 V127 593.2770708065545
L97_127 V97 V127 -1.005213240200553e-12
C97_127 V97 V127 -4.3021428670484e-20

R97_128 V97 V128 2144.7819871245006
L97_128 V97 V128 2.5166311553844775e-11
C97_128 V97 V128 -1.3948847058501154e-20

R97_129 V97 V129 15247.132346937004
L97_129 V97 V129 -1.194000563028712e-12
C97_129 V97 V129 -7.238279118290417e-20

R97_130 V97 V130 3398.7825891684347
L97_130 V97 V130 7.549509279260759e-13
C97_130 V97 V130 1.4640012484304815e-19

R97_131 V97 V131 -3786.4528412778463
L97_131 V97 V131 1.2660735943484445e-12
C97_131 V97 V131 -8.150375096911073e-20

R97_132 V97 V132 -1872.0962571371706
L97_132 V97 V132 3.163616883978778e-12
C97_132 V97 V132 -2.1032504520513263e-20

R97_133 V97 V133 -4353.485450626004
L97_133 V97 V133 1.4572891747593893e-12
C97_133 V97 V133 1.4859990875904772e-19

R97_134 V97 V134 -1749.7891231632505
L97_134 V97 V134 2.7312051333158535e-12
C97_134 V97 V134 -3.6239490798424004e-20

R97_135 V97 V135 798.1469229226612
L97_135 V97 V135 -1.484408691475667e-12
C97_135 V97 V135 5.72891348736731e-20

R97_136 V97 V136 5298.565294179639
L97_136 V97 V136 6.9872178752613654e-12
C97_136 V97 V136 -2.228200087254547e-20

R97_137 V97 V137 -1152.4513259987073
L97_137 V97 V137 2.046051679736641e-12
C97_137 V97 V137 -7.269862383709193e-20

R97_138 V97 V138 -515.0890907955462
L97_138 V97 V138 4.7677938621765e-13
C97_138 V97 V138 -6.930817978255695e-22

R97_139 V97 V139 469.2485073630977
L97_139 V97 V139 -7.307479440002891e-13
C97_139 V97 V139 -3.301901211931895e-20

R97_140 V97 V140 -1946.6690717127187
L97_140 V97 V140 1.307876702902226e-12
C97_140 V97 V140 1.083163680127802e-20

R97_141 V97 V141 -1067.8300345166674
L97_141 V97 V141 3.330127736195203e-12
C97_141 V97 V141 2.5400192423525002e-20

R97_142 V97 V142 26605.886212726633
L97_142 V97 V142 1.2192044723099732e-12
C97_142 V97 V142 -7.686360260953917e-20

R97_143 V97 V143 -2568.4782562205382
L97_143 V97 V143 1.740178128275282e-12
C97_143 V97 V143 2.8779415171388415e-20

R97_144 V97 V144 2067.9029079556253
L97_144 V97 V144 -2.404170191064562e-12
C97_144 V97 V144 1.7190865946159198e-20

R98_98 V98 0 -244.87336779548383
L98_98 V98 0 -1.7340047577193954e-13
C98_98 V98 0 -1.7360050945798786e-19

R98_99 V98 V99 -2225.758836040472
L98_99 V98 V99 2.354994760960885e-12
C98_99 V98 V99 1.8427054920966617e-19

R98_100 V98 V100 37722.93578326295
L98_100 V98 V100 2.3479595004155308e-12
C98_100 V98 V100 2.776642461196999e-19

R98_101 V98 V101 -1470.39386801369
L98_101 V98 V101 -4.295238669475093e-13
C98_101 V98 V101 -8.728703303550729e-19

R98_102 V98 V102 -4385.611053898464
L98_102 V98 V102 -3.862192510547588e-13
C98_102 V98 V102 -9.758774514877146e-19

R98_103 V98 V103 2699.5326772731864
L98_103 V98 V103 5.6175751423543114e-12
C98_103 V98 V103 2.785515061857841e-19

R98_104 V98 V104 -1930.4797845784983
L98_104 V98 V104 -2.535431718150633e-12
C98_104 V98 V104 -3.6660728622608933e-19

R98_105 V98 V105 6765.323620926364
L98_105 V98 V105 5.763293195517025e-13
C98_105 V98 V105 8.938269730105797e-19

R98_106 V98 V106 -732.6435373526193
L98_106 V98 V106 -4.884660211986082e-13
C98_106 V98 V106 -1.4786953427271413e-18

R98_107 V98 V107 -25114.05050030149
L98_107 V98 V107 -6.969036894200775e-13
C98_107 V98 V107 -7.248809879110394e-19

R98_108 V98 V108 617.5575080235143
L98_108 V98 V108 4.783820909094364e-13
C98_108 V98 V108 1.0546733606296658e-18

R98_109 V98 V109 1487.3820272057242
L98_109 V98 V109 6.46680758669653e-11
C98_109 V98 V109 -8.343831981759832e-21

R98_110 V98 V110 915.7118865048905
L98_110 V98 V110 4.189799600174842e-13
C98_110 V98 V110 1.2987370507080428e-18

R98_111 V98 V111 1637.9139032943633
L98_111 V98 V111 2.7905077670474597e-12
C98_111 V98 V111 5.644237113775596e-19

R98_112 V98 V112 670.1266553590449
L98_112 V98 V112 -3.006301815469249e-13
C98_112 V98 V112 -9.167019209168478e-19

R98_113 V98 V113 1243.7559770868922
L98_113 V98 V113 -8.258560013903886e-13
C98_113 V98 V113 -2.8688802371316505e-19

R98_114 V98 V114 -4371.438422337413
L98_114 V98 V114 -6.782445822001781e-13
C98_114 V98 V114 -7.668825118351952e-19

R98_115 V98 V115 -10026.19295056512
L98_115 V98 V115 -1.6576729507785791e-12
C98_115 V98 V115 -3.9880218456249186e-19

R98_116 V98 V116 -481094.22863954096
L98_116 V98 V116 6.090615124346192e-13
C98_116 V98 V116 6.235565683668767e-19

R98_117 V98 V117 2557.0818581767076
L98_117 V98 V117 8.197048140481037e-13
C98_117 V98 V117 4.0867185983013685e-19

R98_118 V98 V118 -3407.390907274616
L98_118 V98 V118 7.501164939747477e-13
C98_118 V98 V118 5.108209039287191e-19

R98_119 V98 V119 1092.121776168523
L98_119 V98 V119 8.591677821090076e-13
C98_119 V98 V119 8.886967131952954e-19

R98_120 V98 V120 2037.4433107763182
L98_120 V98 V120 8.816615403543837e-13
C98_120 V98 V120 3.365751671121618e-19

R98_121 V98 V121 360.00450702517065
L98_121 V98 V121 -5.423350437953982e-13
C98_121 V98 V121 -1.0157348344549955e-19

R98_122 V98 V122 204.78455867903196
L98_122 V98 V122 -4.2928154789767236e-13
C98_122 V98 V122 -3.7255467230062924e-20

R98_123 V98 V123 1176.2365780648497
L98_123 V98 V123 -3.734475149540032e-12
C98_123 V98 V123 1.19196600376144e-19

R98_124 V98 V124 3777.250960101099
L98_124 V98 V124 6.386673832993354e-12
C98_124 V98 V124 3.137824419678773e-19

R98_125 V98 V125 -395.5612831577075
L98_125 V98 V125 4.581207629406659e-13
C98_125 V98 V125 1.2388077132710798e-19

R98_126 V98 V126 -237.29139372429978
L98_126 V98 V126 9.1123686021584e-13
C98_126 V98 V126 -1.1180864020655202e-19

R98_127 V98 V127 421.51998926925677
L98_127 V98 V127 -1.842384771119347e-12
C98_127 V98 V127 2.209739582372763e-20

R98_128 V98 V128 5447.428212901944
L98_128 V98 V128 1.0821768841284204e-10
C98_128 V98 V128 4.628679515626791e-20

R98_129 V98 V129 1055.3888388519033
L98_129 V98 V129 -3.195034842952555e-11
C98_129 V98 V129 1.4103888320748491e-19

R98_130 V98 V130 -1779.6099741558874
L98_130 V98 V130 1.0725641189815502e-12
C98_130 V98 V130 2.8386580486190053e-19

R98_131 V98 V131 -752.0071274619854
L98_131 V98 V131 3.976814617650918e-12
C98_131 V98 V131 -1.7677052711836302e-19

R98_132 V98 V132 -1230.289275838558
L98_132 V98 V132 1.9984363960605964e-12
C98_132 V98 V132 8.142926857202198e-20

R98_133 V98 V133 -980.0203123418607
L98_133 V98 V133 -3.6056076685857034e-12
C98_133 V98 V133 -4.564038241104949e-19

R98_134 V98 V134 -1089.5080338885084
L98_134 V98 V134 2.5007335064907093e-12
C98_134 V98 V134 -2.1550838121318458e-20

R98_135 V98 V135 543.3085026148631
L98_135 V98 V135 -3.115811567013957e-12
C98_135 V98 V135 9.462301519827802e-20

R98_136 V98 V136 -6029.444377060741
L98_136 V98 V136 6.052165225520558e-12
C98_136 V98 V136 2.5821562278702583e-20

R98_137 V98 V137 -676.8666789604096
L98_137 V98 V137 6.594610779682034e-13
C98_137 V98 V137 2.896714057154529e-19

R98_138 V98 V138 -268.08566078384126
L98_138 V98 V138 6.460005923227424e-13
C98_138 V98 V138 1.0642961570465597e-19

R98_139 V98 V139 341.4342509552316
L98_139 V98 V139 -1.2190520150788273e-12
C98_139 V98 V139 -1.2803023943288652e-19

R98_140 V98 V140 -828.9832680576377
L98_140 V98 V140 1.052237255908965e-12
C98_140 V98 V140 1.1133492208620545e-19

R98_141 V98 V141 -985.8776148992374
L98_141 V98 V141 2.823255075644003e-12
C98_141 V98 V141 1.8406772826685457e-20

R98_142 V98 V142 -1318.2649516035601
L98_142 V98 V142 1.1778343594133514e-12
C98_142 V98 V142 1.8990585103165638e-19

R98_143 V98 V143 -1398.0386038220236
L98_143 V98 V143 1.2880826993968072e-11
C98_143 V98 V143 1.285519717382117e-20

R98_144 V98 V144 1041.4439592269805
L98_144 V98 V144 -1.329675361496106e-12
C98_144 V98 V144 -8.918686401090251e-20

R99_99 V99 0 218.81463005472148
L99_99 V99 0 1.1429465747431886e-12
C99_99 V99 0 1.6364119173846674e-19

R99_100 V99 V100 13352.127862332363
L99_100 V99 V100 -2.28975965051375e-11
C99_100 V99 V100 -9.94611542653098e-20

R99_101 V99 V101 3996.9205951030117
L99_101 V99 V101 5.351729060308522e-12
C99_101 V99 V101 1.6916421997497902e-19

R99_102 V99 V102 -4427.496845776493
L99_102 V99 V102 8.321361645010041e-13
C99_102 V99 V102 2.5605440911813507e-19

R99_103 V99 V103 -4082.8033730930547
L99_103 V99 V103 -1.4924806491973495e-12
C99_103 V99 V103 -1.0130705474872688e-19

R99_104 V99 V104 3536.4423315465356
L99_104 V99 V104 4.8897434687025756e-12
C99_104 V99 V104 1.8277379964259278e-19

R99_105 V99 V105 11626.799788814016
L99_105 V99 V105 -1.7601311284575067e-12
C99_105 V99 V105 -2.3144562934461705e-19

R99_106 V99 V106 2296.1968030186217
L99_106 V99 V106 1.2249726155405805e-12
C99_106 V99 V106 3.260904572355225e-19

R99_107 V99 V107 2625.8096977165524
L99_107 V99 V107 8.816762276351498e-13
C99_107 V99 V107 2.602417771782183e-19

R99_108 V99 V108 -1540.1098373253965
L99_108 V99 V108 -1.0923213001814236e-12
C99_108 V99 V108 -3.11468329944429e-19

R99_109 V99 V109 -220100.45304716763
L99_109 V99 V109 -3.850414908622458e-12
C99_109 V99 V109 6.015733117898889e-20

R99_110 V99 V110 -733.884429709975
L99_110 V99 V110 -2.356822402314493e-12
C99_110 V99 V110 -2.8606161219337006e-19

R99_111 V99 V111 1131.350198453741
L99_111 V99 V111 -1.4327986047798988e-12
C99_111 V99 V111 -1.8638730260511716e-19

R99_112 V99 V112 -1144.236602343658
L99_112 V99 V112 1.2151914411886817e-12
C99_112 V99 V112 2.2279392348482026e-19

R99_113 V99 V113 -1580.4701471202554
L99_113 V99 V113 3.173463876073925e-12
C99_113 V99 V113 3.208575351334673e-20

R99_114 V99 V114 -2725.257290046892
L99_114 V99 V114 2.6735121052716043e-12
C99_114 V99 V114 1.7326919631423977e-19

R99_115 V99 V115 -2015.6698907836292
L99_115 V99 V115 1.5511572779033642e-12
C99_115 V99 V115 1.361258881551644e-19

R99_116 V99 V116 2502.2333926824713
L99_116 V99 V116 -1.6680054323938917e-12
C99_116 V99 V116 -1.6646043155441535e-19

R99_117 V99 V117 -1301.1314851125553
L99_117 V99 V117 -4.072107935185256e-12
C99_117 V99 V117 -7.363981248811261e-20

R99_118 V99 V118 3120.1303140046653
L99_118 V99 V118 -3.1008946839650958e-12
C99_118 V99 V118 -7.064123551413821e-20

R99_119 V99 V119 1414.114177659485
L99_119 V99 V119 -1.895248896552425e-12
C99_119 V99 V119 -1.963164915595707e-19

R99_120 V99 V120 -279.44925942041186
L99_120 V99 V120 2.858081476972785e-12
C99_120 V99 V120 -1.0407717632686412e-19

R99_121 V99 V121 -3800.828262239785
L99_121 V99 V121 8.24339333404406e-12
C99_121 V99 V121 2.7900681062503124e-20

R99_122 V99 V122 -209.09050849108115
L99_122 V99 V122 1.63267719289859e-12
C99_122 V99 V122 -9.465640356207304e-21

R99_123 V99 V123 -997.7736937090232
L99_123 V99 V123 1.1525102914338507e-11
C99_123 V99 V123 -2.44083275698434e-20

R99_124 V99 V124 5740.5265485532755
L99_124 V99 V124 -5.037207214026417e-12
C99_124 V99 V124 -1.1049723348841448e-19

R99_125 V99 V125 -1092.7019840908722
L99_125 V99 V125 2.020294004583211e-11
C99_125 V99 V125 -2.5597390618361836e-20

R99_126 V99 V126 160.22886084136366
L99_126 V99 V126 -1.2077577932217202e-12
C99_126 V99 V126 2.146460352648687e-21

R99_127 V99 V127 -210.9753041403841
L99_127 V99 V127 1.358683280227731e-12
C99_127 V99 V127 -9.761639398581697e-22

R99_128 V99 V128 -2779.3273314731387
L99_128 V99 V128 2.680283574924012e-10
C99_128 V99 V128 -1.245816265873816e-20

R99_129 V99 V129 -545.0413229482947
L99_129 V99 V129 4.647009413270082e-12
C99_129 V99 V129 -3.020336023312269e-20

R99_130 V99 V130 788.3111442899508
L99_130 V99 V130 -2.016901441435593e-12
C99_130 V99 V130 -7.336078266774424e-20

R99_131 V99 V131 610.1099719788962
L99_131 V99 V131 3.616889887997399e-11
C99_131 V99 V131 3.643309112912159e-20

R99_132 V99 V132 852.8713297932817
L99_132 V99 V132 -3.8736525042315365e-12
C99_132 V99 V132 -5.417534664661009e-20

R99_133 V99 V133 2984.019195161707
L99_133 V99 V133 4.991220259346005e-12
C99_133 V99 V133 8.219853695433217e-20

R99_134 V99 V134 1140.902195336092
L99_134 V99 V134 -3.588114457606173e-11
C99_134 V99 V134 2.9725809761772786e-20

R99_135 V99 V135 -307.6555355069868
L99_135 V99 V135 2.7814788832361676e-12
C99_135 V99 V135 -6.410047156487928e-20

R99_136 V99 V136 -22908.587664796796
L99_136 V99 V136 1.3636427463454212e-10
C99_136 V99 V136 4.370732820871097e-21

R99_137 V99 V137 -3726.6401158044932
L99_137 V99 V137 -1.017086647032159e-11
C99_137 V99 V137 -7.813021158983521e-20

R99_138 V99 V138 191.70505173349747
L99_138 V99 V138 -1.3097199639769405e-12
C99_138 V99 V138 -1.5791470784681985e-20

R99_139 V99 V139 -164.74325208879569
L99_139 V99 V139 9.712697170534617e-13
C99_139 V99 V139 5.288483110851321e-20

R99_140 V99 V140 640.5319821329936
L99_140 V99 V140 -2.735202457297359e-12
C99_140 V99 V140 -1.681016654314273e-20

R99_141 V99 V141 912.2077052687237
L99_141 V99 V141 -5.70586414375775e-12
C99_141 V99 V141 1.502502178123823e-21

R99_142 V99 V142 617.82630004114
L99_142 V99 V142 -2.560134173886293e-12
C99_142 V99 V142 -6.586217426553356e-20

R99_143 V99 V143 499.5687518536569
L99_143 V99 V143 -3.1343152868980323e-12
C99_143 V99 V143 -9.352792683453349e-22

R99_144 V99 V144 -1243.586708020894
L99_144 V99 V144 3.6357843177060625e-12
C99_144 V99 V144 1.5936661263201895e-20

R100_100 V100 0 919.7562110024622
L100_100 V100 0 6.342986789385959e-13
C100_100 V100 0 3.0475506779593486e-19

R100_101 V100 V101 5386.358357560495
L100_101 V100 V101 1.7308179295913545e-12
C100_101 V100 V101 3.2860327823528795e-19

R100_102 V100 V102 -5619.197104591065
L100_102 V100 V102 -2.259816930081932e-11
C100_102 V100 V102 -1.0359642916327024e-19

R100_103 V100 V103 -15961.082128018432
L100_103 V100 V103 9.29873598011575e-12
C100_103 V100 V103 7.75622319846479e-20

R100_104 V100 V104 5374.739388481149
L100_104 V100 V104 1.8159191184882419e-12
C100_104 V100 V104 5.694587583084614e-19

R100_105 V100 V105 -18778.72168543281
L100_105 V100 V105 -1.9394351146473125e-12
C100_105 V100 V105 -3.915560982742346e-19

R100_106 V100 V106 8897.524872819897
L100_106 V100 V106 1.5563033188510716e-12
C100_106 V100 V106 3.6049805812654533e-19

R100_107 V100 V107 135944.51901283476
L100_107 V100 V107 -2.5502301497964964e-11
C100_107 V100 V107 -6.424395789271619e-20

R100_108 V100 V108 -6642.890965866485
L100_108 V100 V108 -2.6457193061706686e-12
C100_108 V100 V108 -2.9095785564256883e-19

R100_109 V100 V109 6591.988052162745
L100_109 V100 V109 2.087455365780126e-12
C100_109 V100 V109 5.572375711924862e-19

R100_110 V100 V110 -3670.208199017985
L100_110 V100 V110 -1.4323279635457841e-12
C100_110 V100 V110 -3.5017618553127584e-19

R100_111 V100 V111 -76546.50731524739
L100_111 V100 V111 -6.379574553956346e-12
C100_111 V100 V111 -1.598678392593638e-19

R100_112 V100 V112 -26863.37230205911
L100_112 V100 V112 9.489742014056572e-12
C100_112 V100 V112 1.620074625758376e-19

R100_113 V100 V113 -7493.0393157848885
L100_113 V100 V113 5.76868556732046e-12
C100_113 V100 V113 -1.344231531658038e-19

R100_114 V100 V114 -3797.6075066639
L100_114 V100 V114 2.7392936304406547e-12
C100_114 V100 V114 2.569700281579578e-19

R100_115 V100 V115 -8288.762785684969
L100_115 V100 V115 -1.1972638899529783e-11
C100_115 V100 V115 -2.633313252117512e-20

R100_116 V100 V116 -16733.496192946655
L100_116 V100 V116 -5.1456443339016266e-12
C100_116 V100 V116 -1.6085260730153785e-19

R100_117 V100 V117 81773.62353246516
L100_117 V100 V117 -1.9755295028760824e-11
C100_117 V100 V117 1.1781695785664148e-19

R100_118 V100 V118 9367.481947413948
L100_118 V100 V118 -7.689295890205573e-12
C100_118 V100 V118 1.662880690065078e-20

R100_119 V100 V119 30775.34058016269
L100_119 V100 V119 -2.6954706095045734e-12
C100_119 V100 V119 -3.3760918188698183e-19

R100_120 V100 V120 -2818.718411642498
L100_120 V100 V120 -2.359591869512164e-12
C100_120 V100 V120 -1.7587752236669453e-19

R100_121 V100 V121 -14256.83248257666
L100_121 V100 V121 1.280457046906376e-10
C100_121 V100 V121 2.8317215809067446e-20

R100_122 V100 V122 -1602.491436578426
L100_122 V100 V122 -4.037699815698859e-12
C100_122 V100 V122 1.9436411577349952e-20

R100_123 V100 V123 -2043.172071129487
L100_123 V100 V123 -1.3355791459502774e-11
C100_123 V100 V123 -1.2846588287458704e-20

R100_124 V100 V124 -6293.471325643863
L100_124 V100 V124 -2.3068391119275448e-12
C100_124 V100 V124 -2.0782359277734958e-19

R100_125 V100 V125 -7542.485452187418
L100_125 V100 V125 -9.287966000202758e-12
C100_125 V100 V125 -9.083806074770639e-21

R100_126 V100 V126 1544.6628261870537
L100_126 V100 V126 2.34617885314024e-12
C100_126 V100 V126 -5.3179421920192215e-21

R100_127 V100 V127 -2476.6390745197073
L100_127 V100 V127 -3.052715598444603e-12
C100_127 V100 V127 -4.822287893923622e-20

R100_128 V100 V128 -5703.679229147514
L100_128 V100 V128 2.681694556393091e-12
C100_128 V100 V128 1.0347635998171722e-20

R100_129 V100 V129 -1775.1822282041458
L100_129 V100 V129 -4.11483286218741e-12
C100_129 V100 V129 -5.64240887460942e-20

R100_130 V100 V130 1909.4937683237085
L100_130 V100 V130 4.835626316478197e-12
C100_130 V100 V130 2.8264536204068255e-21

R100_131 V100 V131 1866.188369284277
L100_131 V100 V131 4.714543990108505e-12
C100_131 V100 V131 1.9301091228172427e-20

R100_132 V100 V132 22679.542112212883
L100_132 V100 V132 -9.300722107295172e-12
C100_132 V100 V132 -1.0983833325042958e-19

R100_133 V100 V133 8414.48953374713
L100_133 V100 V133 3.85661394080254e-12
C100_133 V100 V133 8.675906943223952e-20

R100_134 V100 V134 11760.029588300325
L100_134 V100 V134 2.8549663703786045e-11
C100_134 V100 V134 1.0848153769608074e-21

R100_135 V100 V135 -3122.7218969089786
L100_135 V100 V135 -4.291562377303305e-12
C100_135 V100 V135 -2.494559232908307e-20

R100_136 V100 V136 318451.8905807358
L100_136 V100 V136 4.020871311554224e-12
C100_136 V100 V136 1.5460739007064332e-20

R100_137 V100 V137 -10327.271883450532
L100_137 V100 V137 -8.08682185870545e-12
C100_137 V100 V137 -1.0413569394431403e-19

R100_138 V100 V138 1183.4721765293573
L100_138 V100 V138 2.4019584971041783e-12
C100_138 V100 V138 -4.9920489282599914e-20

R100_139 V100 V139 -1947.7305745407825
L100_139 V100 V139 -2.8738200889935518e-12
C100_139 V100 V139 1.920916351834957e-20

R100_140 V100 V140 12157.29032503263
L100_140 V100 V140 6.04503700131635e-12
C100_140 V100 V140 -3.862320390940038e-20

R100_141 V100 V141 9994.752201517844
L100_141 V100 V141 -1.4722043171058332e-11
C100_141 V100 V141 3.322080971412879e-20

R100_142 V100 V142 1980.0671323197496
L100_142 V100 V142 7.937663929429947e-12
C100_142 V100 V142 -7.560398511726049e-20

R100_143 V100 V143 3604.2610387952705
L100_143 V100 V143 4.6910471972099076e-12
C100_143 V100 V143 -4.306444127727653e-21

R100_144 V100 V144 -16175.745077449601
L100_144 V100 V144 -1.876164325611291e-11
C100_144 V100 V144 5.6149311446353396e-21

R101_101 V101 0 -3789.3896757169346
L101_101 V101 0 -2.345370777970541e-13
C101_101 V101 0 6.294688827675308e-19

R101_102 V101 V102 -2069.2881414949143
L101_102 V101 V102 -6.020530479055814e-13
C101_102 V101 V102 -9.504595044723406e-19

R101_103 V101 V103 -20317.884201516023
L101_103 V101 V103 -4.554304039144283e-12
C101_103 V101 V103 -2.6154981687895946e-20

R101_104 V101 V104 103904.46244251628
L101_104 V101 V104 -2.350132865264774e-12
C101_104 V101 V104 -4.2230410836259795e-19

R101_105 V101 V105 3663.8410930502882
L101_105 V101 V105 6.806051338634436e-13
C101_105 V101 V105 8.615754166709673e-19

R101_106 V101 V106 -4037.3910696460593
L101_106 V101 V106 -5.671589441603507e-13
C101_106 V101 V106 -1.4755632215816579e-18

R101_107 V101 V107 -17332.87133774135
L101_107 V101 V107 -1.4174109769281207e-12
C101_107 V101 V107 -3.111696021518231e-19

R101_108 V101 V108 2212.0860698596116
L101_108 V101 V108 6.152873414314216e-13
C101_108 V101 V108 1.2843578673702061e-18

R101_109 V101 V109 18226.80864965431
L101_109 V101 V109 -3.626205728214976e-12
C101_109 V101 V109 3.1186054400893874e-21

R101_110 V101 V110 3022.889252607962
L101_110 V101 V110 4.22313598366946e-13
C101_110 V101 V110 1.4230284271127214e-18

R101_111 V101 V111 5047.002146859521
L101_111 V101 V111 -4.3833292704265694e-10
C101_111 V101 V111 3.6241582922538594e-19

R101_112 V101 V112 -1078.353804400717
L101_112 V101 V112 -3.4875239340832137e-13
C101_112 V101 V112 -1.168987018898909e-18

R101_113 V101 V113 -1691.0372537105513
L101_113 V101 V113 -9.513108600586437e-13
C101_113 V101 V113 -3.5056276690112107e-19

R101_114 V101 V114 -7682.0799143043505
L101_114 V101 V114 -9.120534719861583e-13
C101_114 V101 V114 -8.781042377277443e-19

R101_115 V101 V115 -13273.525730549216
L101_115 V101 V115 -1.871097606114296e-11
C101_115 V101 V115 -1.736031265248466e-19

R101_116 V101 V116 2210.2359423067937
L101_116 V101 V116 7.689535566051421e-13
C101_116 V101 V116 7.133267815912396e-19

R101_117 V101 V117 5102.241603854677
L101_117 V101 V117 9.251738584709652e-13
C101_117 V101 V117 5.651270551657754e-19

R101_118 V101 V118 2865.483191258377
L101_118 V101 V118 8.914930212519219e-13
C101_118 V101 V118 5.228961617639489e-19

R101_119 V101 V119 3866.7619085992533
L101_119 V101 V119 1.274915995015097e-12
C101_119 V101 V119 8.978920240585167e-19

R101_120 V101 V120 -2207.402431354128
L101_120 V101 V120 7.234383474881253e-13
C101_120 V101 V120 3.6079477413627455e-19

R101_121 V101 V121 -3140.4979630763473
L101_121 V101 V121 -5.832267863019492e-13
C101_121 V101 V121 -2.4839506560231294e-20

R101_122 V101 V122 -735.9925904070218
L101_122 V101 V122 -6.261987576533872e-13
C101_122 V101 V122 -1.3607978612305823e-19

R101_123 V101 V123 16577.155514746482
L101_123 V101 V123 1.378222794777259e-11
C101_123 V101 V123 6.009111477432439e-20

R101_124 V101 V124 2157.5944206124323
L101_124 V101 V124 3.809498059843916e-12
C101_124 V101 V124 2.3548879218496175e-19

R101_125 V101 V125 3484.151329418823
L101_125 V101 V125 4.794252791645963e-13
C101_125 V101 V125 8.725601601442287e-20

R101_126 V101 V126 723.8558368651155
L101_126 V101 V126 3.7633696826578654e-12
C101_126 V101 V126 -1.4295894109791009e-19

R101_127 V101 V127 -938.9635683611376
L101_127 V101 V127 2.5581350159457065e-11
C101_127 V101 V127 4.4806929953778466e-20

R101_128 V101 V128 -2896.4864512660974
L101_128 V101 V128 -2.5587312706828442e-11
C101_128 V101 V128 6.211801176656768e-20

R101_129 V101 V129 8691.714206419876
L101_129 V101 V129 1.4090607040574944e-12
C101_129 V101 V129 2.9501707955563116e-19

R101_130 V101 V130 -14795.746974934915
L101_130 V101 V130 4.380467135265056e-12
C101_130 V101 V130 3.4723564549528758e-19

R101_131 V101 V131 -23215.321734103727
L101_131 V101 V131 -5.233432492298414e-12
C101_131 V101 V131 -1.1995537366195664e-19

R101_132 V101 V132 3003.4786624051653
L101_132 V101 V132 3.065212613052016e-12
C101_132 V101 V132 8.74172465122713e-20

R101_133 V101 V133 -8956.204117888283
L101_133 V101 V133 -2.7365213211141253e-12
C101_133 V101 V133 -4.889709219292441e-19

R101_134 V101 V134 3429.571698486269
L101_134 V101 V134 6.423981685561233e-12
C101_134 V101 V134 -7.977097862681077e-20

R101_135 V101 V135 -1422.1626406184073
L101_135 V101 V135 -9.424757907985566e-11
C101_135 V101 V135 4.931298705001172e-20

R101_136 V101 V136 -5670.534781694945
L101_136 V101 V136 1.1205282544411078e-10
C101_136 V101 V136 6.857045518130561e-21

R101_137 V101 V137 2520.2923903265014
L101_137 V101 V137 6.480115116363815e-13
C101_137 V101 V137 3.5432497664935854e-19

R101_138 V101 V138 991.5169589245613
L101_138 V101 V138 2.0774472288381494e-12
C101_138 V101 V138 9.130250586037213e-20

R101_139 V101 V139 -702.0194934880006
L101_139 V101 V139 -8.370014358406932e-12
C101_139 V101 V139 -1.3078874436499205e-19

R101_140 V101 V140 3100.9668295839765
L101_140 V101 V140 1.6750403772980407e-12
C101_140 V101 V140 1.2336466486128041e-19

R101_141 V101 V141 1827.4673112736525
L101_141 V101 V141 2.970007497064598e-12
C101_141 V101 V141 2.4470117586378683e-21

R101_142 V101 V142 27110.79737591517
L101_142 V101 V142 4.436976454892209e-12
C101_142 V101 V142 2.1618365358442905e-19

R101_143 V101 V143 3942.2772388180874
L101_143 V101 V143 -2.5205102814959474e-12
C101_143 V101 V143 -5.927980139667473e-20

R101_144 V101 V144 -4050.7372644266698
L101_144 V101 V144 -1.7711400510549759e-12
C101_144 V101 V144 -1.4412769919502295e-19

R102_102 V102 0 -202.18804503151952
L102_102 V102 0 -1.8631475143425856e-13
C102_102 V102 0 -8.591089153720095e-19

R102_103 V102 V103 1338.1424250336593
L102_103 V102 V103 3.5198261842552505e-13
C102_103 V102 V103 2.052993278602533e-18

R102_104 V102 V104 -4514.989282682254
L102_104 V102 V104 2.197971971297442e-11
C102_104 V102 V104 -2.1224457195963464e-19

R102_105 V102 V105 1848.3730388785418
L102_105 V102 V105 3.779655010771812e-13
C102_105 V102 V105 1.289113663296454e-18

R102_106 V102 V106 -861.9837511432297
L102_106 V102 V106 -2.6089908524651904e-13
C102_106 V102 V106 -2.50129637417748e-18

R102_107 V102 V107 -811.9134787428281
L102_107 V102 V107 -2.0564905354955398e-13
C102_107 V102 V107 -2.9722838796118645e-18

R102_108 V102 V108 720.3129896864987
L102_108 V102 V108 2.4311628292588837e-13
C102_108 V102 V108 2.6832705669468864e-18

R102_109 V102 V109 1847.2190209861774
L102_109 V102 V109 5.50305876589172e-13
C102_109 V102 V109 1.2390551596262282e-18

R102_110 V102 V110 925.2219652160641
L102_110 V102 V110 4.2001718457998353e-13
C102_110 V102 V110 1.754192220809105e-18

R102_111 V102 V111 4762.2538229540905
L102_111 V102 V111 4.154719658472837e-13
C102_111 V102 V111 1.4022631987854426e-18

R102_112 V102 V112 -1502.7870327907415
L102_112 V102 V112 -2.0117936722901384e-13
C102_112 V102 V112 -2.2323384826131672e-18

R102_113 V102 V113 16287.84822233017
L102_113 V102 V113 -4.343352103909877e-13
C102_113 V102 V113 -1.0003284570586982e-18

R102_114 V102 V114 -1598.0936132005415
L102_114 V102 V114 -4.4351893390079676e-13
C102_114 V102 V114 -1.011635106541577e-18

R102_115 V102 V115 -1731.1498780020381
L102_115 V102 V115 -3.698441046180512e-13
C102_115 V102 V115 -1.620902025646081e-18

R102_116 V102 V116 1945.4933358752376
L102_116 V102 V116 3.368377770986841e-13
C102_116 V102 V116 1.505926289891802e-18

R102_117 V102 V117 1275.393056377419
L102_117 V102 V117 5.339412807169299e-13
C102_117 V102 V117 1.3903179049607723e-18

R102_118 V102 V118 4058.4129186058194
L102_118 V102 V118 4.488772415648879e-13
C102_118 V102 V118 9.450872084573432e-19

R102_119 V102 V119 2142.6811219188644
L102_119 V102 V119 4.549086100437725e-13
C102_119 V102 V119 1.116392572319361e-18

R102_120 V102 V120 767.8623874904252
L102_120 V102 V120 -9.46621090583719e-13
C102_120 V102 V120 5.065378043421736e-19

R102_121 V102 V121 6580.709529366518
L102_121 V102 V121 -5.748782687610993e-13
C102_121 V102 V121 -2.2173635239629697e-19

R102_122 V102 V122 616.4868142336707
L102_122 V102 V122 -2.299697636474921e-13
C102_122 V102 V122 1.0342072056177228e-21

R102_123 V102 V123 30811.320990434946
L102_123 V102 V123 -1.2439502857208891e-12
C102_123 V102 V123 2.1979320769330096e-19

R102_124 V102 V124 -2010.5775833118123
L102_124 V102 V124 2.5007185018246524e-12
C102_124 V102 V124 2.595020042356318e-19

R102_125 V102 V125 6013.086306440714
L102_125 V102 V125 8.513696928795546e-13
C102_125 V102 V125 2.627747172341523e-19

R102_126 V102 V126 -449.1091878466406
L102_126 V102 V126 2.445394177502384e-13
C102_126 V102 V126 -3.912852825851301e-19

R102_127 V102 V127 633.4310395115798
L102_127 V102 V127 -3.0254612639611593e-13
C102_127 V102 V127 -4.4671614287631465e-20

R102_128 V102 V128 1870.274856178189
L102_128 V102 V128 -3.661881425960846e-12
C102_128 V102 V128 8.04209137304233e-20

R102_129 V102 V129 8743.741540777
L102_129 V102 V129 -8.782492309370792e-13
C102_129 V102 V129 2.028761984690082e-19

R102_130 V102 V130 1754.0329108264407
L102_130 V102 V130 3.6146110508732403e-13
C102_130 V102 V130 8.833738698241003e-19

R102_131 V102 V131 -2997.3011519346524
L102_131 V102 V131 3.7284111921692025e-12
C102_131 V102 V131 -7.955654583618172e-19

R102_132 V102 V132 -2902.324852143466
L102_132 V102 V132 9.30871007205734e-13
C102_132 V102 V132 1.0788652250762704e-19

R102_133 V102 V133 -4029.972729589686
L102_133 V102 V133 -1.7107231529668707e-12
C102_133 V102 V133 -6.125206058188849e-19

R102_134 V102 V134 -2766.908424532908
L102_134 V102 V134 1.7293415747055878e-12
C102_134 V102 V134 -1.4850799539304118e-19

R102_135 V102 V135 825.8464281752645
L102_135 V102 V135 -5.178933231543223e-13
C102_135 V102 V135 3.069039443193879e-19

R102_136 V102 V136 3889.1269875054745
L102_136 V102 V136 -2.7277584682345688e-11
C102_136 V102 V136 -5.482293272801322e-20

R102_137 V102 V137 -21907.535231943748
L102_137 V102 V137 9.286531324910018e-13
C102_137 V102 V137 3.034923194554039e-19

R102_138 V102 V138 -783.9290788607176
L102_138 V102 V138 2.1532293609949736e-13
C102_138 V102 V138 3.2763160260810213e-19

R102_139 V102 V139 523.1341763529167
L102_139 V102 V139 -2.154321654685964e-13
C102_139 V102 V139 -3.8095081234500137e-19

R102_140 V102 V140 -5457.411381905899
L102_140 V102 V140 4.961432184100668e-13
C102_140 V102 V140 2.617696892049525e-19

R102_141 V102 V141 -1362.6128333161712
L102_141 V102 V141 8.889086235958419e-13
C102_141 V102 V141 1.29099247317535e-19

R102_142 V102 V142 5618.1716204533295
L102_142 V102 V142 4.630691438718857e-13
C102_142 V102 V142 3.5374654193786893e-19

R102_143 V102 V143 -2299.3141907834147
L102_143 V102 V143 6.95668002869527e-13
C102_143 V102 V143 3.951510797646617e-20

R102_144 V102 V144 6111.159779850832
L102_144 V102 V144 -7.475817613977801e-13
C102_144 V102 V144 -1.5693322072430586e-19

R103_103 V103 0 -341.3845426044673
L103_103 V103 0 1.5403844179684988e-12
C103_103 V103 0 9.20981373803157e-19

R103_104 V103 V104 -8012.721262734356
L103_104 V103 V104 3.452609260216155e-12
C103_104 V103 V104 2.179421066825109e-19

R103_105 V103 V105 -8178.0155440046765
L103_105 V103 V105 -1.1201789100199285e-12
C103_105 V103 V105 -5.62171695230807e-19

R103_106 V103 V106 5844.351004121956
L103_106 V103 V106 6.160531446943657e-13
C103_106 V103 V106 1.0993985482180268e-18

R103_107 V103 V107 1121.6253530320162
L103_107 V103 V107 3.796778916038296e-13
C103_107 V103 V107 1.886032211850438e-18

R103_108 V103 V108 -3880.5574156549997
L103_108 V103 V108 -5.1413767725981e-13
C103_108 V103 V108 -1.3078647258515325e-18

R103_109 V103 V109 -4632.11319236794
L103_109 V103 V109 -1.0464625521555764e-12
C103_109 V103 V109 -5.436113059977572e-19

R103_110 V103 V110 21194.560055950136
L103_110 V103 V110 -1.1574108369464673e-11
C103_110 V103 V110 -4.2905879491034004e-19

R103_111 V103 V111 -2088.216601629851
L103_111 V103 V111 -5.385870222385952e-13
C103_111 V103 V111 -8.120375740100317e-19

R103_112 V103 V112 1364.1495643534827
L103_112 V103 V112 7.399234415760207e-13
C103_112 V103 V112 1.0363825224749704e-18

R103_113 V103 V113 1439.0500872200364
L103_113 V103 V113 1.4839866152138765e-12
C103_113 V103 V113 4.1736001799777466e-19

R103_114 V103 V114 -2855.6678915513635
L103_114 V103 V114 3.2647666638181807e-12
C103_114 V103 V114 2.2206088570119404e-19

R103_115 V103 V115 2305.516823874632
L103_115 V103 V115 5.941265407894132e-13
C103_115 V103 V115 1.082199496989335e-18

R103_116 V103 V116 -2605.616094647192
L103_116 V103 V116 -7.683485283920825e-13
C103_116 V103 V116 -7.746978881671995e-19

R103_117 V103 V117 -5878.304232961915
L103_117 V103 V117 -2.3740496219326783e-12
C103_117 V103 V117 -6.099688057819611e-19

R103_118 V103 V118 -3584.4860088657874
L103_118 V103 V118 -2.0031740668517255e-12
C103_118 V103 V118 -3.0882145474462243e-19

R103_119 V103 V119 7891.798202949945
L103_119 V103 V119 -9.81282938762858e-13
C103_119 V103 V119 -3.74116216534974e-19

R103_120 V103 V120 2557.277626217983
L103_120 V103 V120 5.853546214701467e-13
C103_120 V103 V120 -2.1989386986957973e-19

R103_121 V103 V121 1875.7016966945878
L103_121 V103 V121 -2.539990226508176e-12
C103_121 V103 V121 1.2322922813806772e-19

R103_122 V103 V122 822.1297401960887
L103_122 V103 V122 8.242773376322652e-13
C103_122 V103 V122 -1.1136205699050775e-20

R103_123 V103 V123 -3823.245440737129
L103_123 V103 V123 4.484174449310781e-12
C103_123 V103 V123 4.131544338314105e-20

R103_124 V103 V124 -1465.8073391143198
L103_124 V103 V124 -2.3597135003743944e-12
C103_124 V103 V124 -6.921864180723032e-20

R103_125 V103 V125 -2051.4322422146365
L103_125 V103 V125 1.1442689220013014e-12
C103_125 V103 V125 -1.3414575361134447e-19

R103_126 V103 V126 -785.2352811941465
L103_126 V103 V126 -4.855041415673667e-13
C103_126 V103 V126 2.5939716564316154e-19

R103_127 V103 V127 984.350482263298
L103_127 V103 V127 4.621599153158802e-13
C103_127 V103 V127 2.8609839093735545e-20

R103_128 V103 V128 1986.9288178566553
L103_128 V103 V128 6.089789064642137e-12
C103_128 V103 V128 6.95987166144481e-21

R103_129 V103 V129 -3033.653138495313
L103_129 V103 V129 1.5970143236824135e-12
C103_129 V103 V129 4.1869547496309413e-20

R103_130 V103 V130 2486.819943113936
L103_130 V103 V130 -1.0403967133551923e-12
C103_130 V103 V130 -4.5297960414000235e-19

R103_131 V103 V131 1982.6117667493365
L103_131 V103 V131 2.302336041114616e-12
C103_131 V103 V131 5.197219748819184e-19

R103_132 V103 V132 -3731.2506632999352
L103_132 V103 V132 -1.9913180569218875e-12
C103_132 V103 V132 -4.3629189798662106e-20

R103_133 V103 V133 11241.136463433832
L103_133 V103 V133 2.111464318936233e-12
C103_133 V103 V133 2.39052921974977e-19

R103_134 V103 V134 -4070.629155305708
L103_134 V103 V134 -4.73990179662256e-12
C103_134 V103 V134 2.810547148625118e-20

R103_135 V103 V135 1650.7359214858388
L103_135 V103 V135 7.93011496414265e-13
C103_135 V103 V135 -1.3578819660630678e-19

R103_136 V103 V136 3411.888670325792
L103_136 V103 V136 6.2279109937313095e-12
C103_136 V103 V136 2.7090724026248036e-20

R103_137 V103 V137 -2170.6375037738762
L103_137 V103 V137 2.5073034594363387e-12
C103_137 V103 V137 -6.690297678786919e-20

R103_138 V103 V138 -1324.2316064802649
L103_138 V103 V138 -5.419583258078774e-13
C103_138 V103 V138 -1.4079133370233315e-19

R103_139 V103 V139 715.581759067469
L103_139 V103 V139 3.352096606515839e-13
C103_139 V103 V139 2.3888122364511987e-19

R103_140 V103 V140 -6377.163823697953
L103_140 V103 V140 -1.2696225072989509e-12
C103_140 V103 V140 -1.2370790353194165e-19

R103_141 V103 V141 -1290.5893272293442
L103_141 V103 V141 -1.894302095415236e-12
C103_141 V103 V141 -5.603495426796099e-20

R103_142 V103 V142 2543.912265586887
L103_142 V103 V142 -2.0203913070179514e-12
C103_142 V103 V142 -3.1074819192146697e-20

R103_143 V103 V143 -6760.080691409479
L103_143 V103 V143 -9.744586344306372e-13
C103_143 V103 V143 -7.572955802277438e-20

R103_144 V103 V144 4877.029611350582
L103_144 V103 V144 2.258605251098314e-12
C103_144 V103 V144 4.2099340100943155e-20

R104_104 V104 0 1104.9082666999784
L104_104 V104 0 -6.034305355045999e-13
C104_104 V104 0 -5.410716343136265e-19

R104_105 V104 V105 3307.8022020713443
L104_105 V104 V105 1.655573345125423e-12
C104_105 V104 V105 5.791018061565831e-19

R104_106 V104 V106 6890.957554547848
L104_106 V104 V106 -4.8561224450254795e-12
C104_106 V104 V106 -3.0909573139448676e-19

R104_107 V104 V107 -69867.97460777989
L104_107 V104 V107 -1.771520608453642e-11
C104_107 V104 V107 -1.3714592984972563e-19

R104_108 V104 V108 -15897.800049854448
L104_108 V104 V108 1.2075117240945458e-12
C104_108 V104 V108 8.008443495354161e-19

R104_109 V104 V109 -1681.902861140197
L104_109 V104 V109 -6.680425035834679e-13
C104_109 V104 V109 -1.065377630633656e-18

R104_110 V104 V110 -3582.9129728570506
L104_110 V104 V110 5.821550138873088e-12
C104_110 V104 V110 1.9973739209643138e-19

R104_111 V104 V111 67963.15332007877
L104_111 V104 V111 3.801713965952618e-12
C104_111 V104 V111 2.3494689403983037e-19

R104_112 V104 V112 -1462.0095205742691
L104_112 V104 V112 -4.798998383208711e-12
C104_112 V104 V112 -3.196866205400327e-19

R104_113 V104 V113 -14510.915119289786
L104_113 V104 V113 1.7420660714485188e-12
C104_113 V104 V113 2.837059083734666e-19

R104_114 V104 V114 -2517.549222212636
L104_114 V104 V114 8.252318475950722e-12
C104_114 V104 V114 -7.115562759859454e-20

R104_115 V104 V115 -5917.25614337209
L104_115 V104 V115 -1.4285028859110387e-11
C104_115 V104 V115 -1.523756506927805e-19

R104_116 V104 V116 4640.431805601681
L104_116 V104 V116 1.9222398645640705e-12
C104_116 V104 V116 4.952276798878088e-19

R104_117 V104 V117 -8314.598020225312
L104_117 V104 V117 -6.1396307976590355e-12
C104_117 V104 V117 -6.009666719517338e-20

R104_118 V104 V118 7915.7685151344895
L104_118 V104 V118 -1.9285648343331374e-12
C104_118 V104 V118 -2.7074191202053532e-19

R104_119 V104 V119 7238.855191487849
L104_119 V104 V119 3.1178513785394037e-12
C104_119 V104 V119 3.3649555354361557e-19

R104_120 V104 V120 -3320.457686347518
L104_120 V104 V120 2.095487539711194e-12
C104_120 V104 V120 3.42823126200376e-19

R104_121 V104 V121 -1380.2676134761493
L104_121 V104 V121 4.822756194204728e-12
C104_121 V104 V121 4.397039640718487e-20

R104_122 V104 V122 -550.4833011658386
L104_122 V104 V122 4.158237699302358e-12
C104_122 V104 V122 -7.265283607325564e-20

R104_123 V104 V123 -1410.011741200843
L104_123 V104 V123 9.080706671985889e-12
C104_123 V104 V123 -7.422452634564443e-20

R104_124 V104 V124 -8005.151700510543
L104_124 V104 V124 3.190122180840683e-12
C104_124 V104 V124 3.796030900469882e-19

R104_125 V104 V125 2095.0876347389526
L104_125 V104 V125 2.3111142717472147e-11
C104_125 V104 V125 1.2160888127729303e-20

R104_126 V104 V126 605.4795400456434
L104_126 V104 V126 -2.9804523987784764e-12
C104_126 V104 V126 -2.4696342699600473e-20

R104_127 V104 V127 -1047.199620084315
L104_127 V104 V127 5.153078146961943e-12
C104_127 V104 V127 6.834321316122218e-20

R104_128 V104 V128 -166387.53885011174
L104_128 V104 V128 2.3570245335902543e-12
C104_128 V104 V128 6.167320467365234e-20

R104_129 V104 V129 -1300.461646895088
L104_129 V104 V129 3.4418821314169367e-12
C104_129 V104 V129 1.220895803801969e-19

R104_130 V104 V130 1277.2957623857078
L104_130 V104 V130 9.742211142919106e-12
C104_130 V104 V130 1.812585948782281e-19

R104_131 V104 V131 1147.5972554644404
L104_131 V104 V131 -8.066576905047958e-12
C104_131 V104 V131 -3.3378753621156586e-20

R104_132 V104 V132 3048.54172860563
L104_132 V104 V132 2.0445640892041474e-12
C104_132 V104 V132 3.692123699256023e-19

R104_133 V104 V133 3343.188591165882
L104_133 V104 V133 -6.289406454988249e-12
C104_133 V104 V133 -1.2652942120350598e-19

R104_134 V104 V134 3371.282236519536
L104_134 V104 V134 -3.536837815071239e-11
C104_134 V104 V134 -3.526604405936343e-20

R104_135 V104 V135 -1345.361796239471
L104_135 V104 V135 5.732115721446454e-12
C104_135 V104 V135 7.455468757907403e-20

R104_136 V104 V136 10146.358678125756
L104_136 V104 V136 -5.964521533779381e-12
C104_136 V104 V136 -1.8568000388949193e-19

R104_137 V104 V137 3117.119682136525
L104_137 V104 V137 1.6601261351347192e-11
C104_137 V104 V137 1.4132255087453554e-19

R104_138 V104 V138 545.7383212863891
L104_138 V104 V138 -2.5418244053733122e-12
C104_138 V104 V138 4.3131300148318515e-20

R104_139 V104 V139 -795.7824857609903
L104_139 V104 V139 7.198369778844759e-12
C104_139 V104 V139 -6.951266871131424e-20

R104_140 V104 V140 1995.0121106735508
L104_140 V104 V140 2.3831857673741545e-11
C104_140 V104 V140 1.559986460479584e-20

R104_141 V104 V141 4480.658401393304
L104_141 V104 V141 -3.680187927597561e-12
C104_141 V104 V141 -9.651666575646959e-20

R104_142 V104 V142 1261.4395672676999
L104_142 V104 V142 -4.622137802442368e-12
C104_142 V104 V142 9.034545489992613e-20

R104_143 V104 V143 2006.2147210288847
L104_143 V104 V143 -1.1254470419962126e-11
C104_143 V104 V143 3.8174826077622565e-20

R104_144 V104 V144 -3151.3654677717773
L104_144 V104 V144 -2.057380514350661e-11
C104_144 V104 V144 5.362722834758656e-20

R105_105 V105 0 264.3809894161899
L105_105 V105 0 2.1137381541172184e-13
C105_105 V105 0 3.1126048497964584e-19

R105_106 V105 V106 1175.5518703460893
L105_106 V105 V106 2.9724919272130797e-13
C105_106 V105 V106 2.0951309192174786e-18

R105_107 V105 V107 2593.161551231622
L105_107 V105 V107 4.843922119681818e-13
C105_107 V105 V107 1.1449658699411116e-18

R105_108 V105 V108 -1644.1891340855195
L105_108 V105 V108 -4.72921951097128e-13
C105_108 V105 V108 -1.21578806436033e-18

R105_109 V105 V109 39687.73511391151
L105_109 V105 V109 -7.346599099652428e-12
C105_109 V105 V109 1.4306266021125354e-19

R105_110 V105 V110 -1352.438958589725
L105_110 V105 V110 -3.8157544703978113e-13
C105_110 V105 V110 -1.730451628026087e-18

R105_111 V105 V111 -5164.341526899828
L105_111 V105 V111 -6.768428844612114e-13
C105_111 V105 V111 -8.470343862156715e-19

R105_112 V105 V112 7894.606029193393
L105_112 V105 V112 4.3877532467911607e-13
C105_112 V105 V112 1.0496132232023799e-18

R105_113 V105 V113 -4318.194554129054
L105_113 V105 V113 1.0810263649768694e-12
C105_113 V105 V113 3.452034924663703e-19

R105_114 V105 V114 1704.115796691682
L105_114 V105 V114 6.086659782499883e-13
C105_114 V105 V114 9.784627338522167e-19

R105_115 V105 V115 4015.4056172759892
L105_115 V105 V115 9.662333042149888e-13
C105_115 V105 V115 6.002605551353907e-19

R105_116 V105 V116 -5514.757892704089
L105_116 V105 V116 -6.27160348290081e-13
C105_116 V105 V116 -7.608452130814284e-19

R105_117 V105 V117 -4356.073525042678
L105_117 V105 V117 -1.139204095082181e-12
C105_117 V105 V117 -4.597919707144864e-19

R105_118 V105 V118 -5975.702490979508
L105_118 V105 V118 -6.782420869637498e-13
C105_118 V105 V118 -7.490644863080403e-19

R105_119 V105 V119 -1812.3281517907026
L105_119 V105 V119 -5.356661440822652e-13
C105_119 V105 V119 -1.146811279579453e-18

R105_120 V105 V120 -2122.783716783921
L105_120 V105 V120 1.1611773188161446e-11
C105_120 V105 V120 -3.8485915090943486e-19

R105_121 V105 V121 -4064.491945108482
L105_121 V105 V121 1.2971859427377467e-12
C105_121 V105 V121 2.250362175065995e-19

R105_122 V105 V122 -1147.1549857089533
L105_122 V105 V122 8.368796085961864e-13
C105_122 V105 V122 2.095699098102284e-20

R105_123 V105 V123 10149.362583752349
L105_123 V105 V123 9.519263466087674e-11
C105_123 V105 V123 -1.496687383578819e-19

R105_124 V105 V124 4452.711286713753
L105_124 V105 V124 -1.9737933177981465e-12
C105_124 V105 V124 -3.891417218954881e-19

R105_125 V105 V125 4271.965157005606
L105_125 V105 V125 -1.8703079928463526e-12
C105_125 V105 V125 -1.6941829859931906e-19

R105_126 V105 V126 972.4868052144676
L105_126 V105 V126 -9.043839951076361e-13
C105_126 V105 V126 1.659242055966623e-19

R105_127 V105 V127 -1407.7201385593955
L105_127 V105 V127 9.884837887853872e-13
C105_127 V105 V127 -3.705395856750054e-20

R105_128 V105 V128 -3366.934182470262
L105_128 V105 V128 -1.4491628403892214e-11
C105_128 V105 V128 -1.5162593510506716e-19

R105_129 V105 V129 6322.2701535977585
L105_129 V105 V129 7.212230911192128e-12
C105_129 V105 V129 -1.5205098682931428e-19

R105_130 V105 V130 -2108.6744640710444
L105_130 V105 V130 -9.554375964914135e-13
C105_130 V105 V130 -4.387985151054176e-19

R105_131 V105 V131 -19006.73544471612
L105_131 V105 V131 5.234158578122394e-12
C105_131 V105 V131 3.1329508204488337e-19

R105_132 V105 V132 5858.3261124144165
L105_132 V105 V132 -2.0324231998798772e-12
C105_132 V105 V132 -1.61792829615424e-19

R105_133 V105 V133 4952.318772076208
L105_133 V105 V133 1.0286064980246309e-12
C105_133 V105 V133 6.699005009814034e-19

R105_134 V105 V134 6652.287764515622
L105_134 V105 V134 -1.2578775465001916e-11
C105_134 V105 V134 -4.9324001855297735e-21

R105_135 V105 V135 -1845.931490323797
L105_135 V105 V135 1.914186084770119e-12
C105_135 V105 V135 -1.3354932487594742e-19

R105_136 V105 V136 -6415.423426887715
L105_136 V105 V136 5.139743417125092e-12
C105_136 V105 V136 1.0444998150354664e-19

R105_137 V105 V137 5409.727414587801
L105_137 V105 V137 -1.8461000336168923e-12
C105_137 V105 V137 -3.313344197067984e-19

R105_138 V105 V138 1997.8056532242424
L105_138 V105 V138 -8.566607985516862e-13
C105_138 V105 V138 -1.0017966389979252e-19

R105_139 V105 V139 -1235.6857056718075
L105_139 V105 V139 6.437540688934394e-13
C105_139 V105 V139 2.341189148929324e-19

R105_140 V105 V140 10982.546779006056
L105_140 V105 V140 -1.4684561407006554e-12
C105_140 V105 V140 -6.249721249156603e-20

R105_141 V105 V141 2177.247911448336
L105_141 V105 V141 -2.866648477460163e-12
C105_141 V105 V141 -9.081568120137588e-21

R105_142 V105 V142 -2884.1348142596617
L105_142 V105 V142 -1.1649832384305045e-12
C105_142 V105 V142 -2.5952673760611805e-19

R105_143 V105 V143 10510.008298594368
L105_143 V105 V143 -2.4791720775104695e-12
C105_143 V105 V143 -2.2877729445104264e-20

R105_144 V105 V144 -7372.115308478185
L105_144 V105 V144 2.4125065538131005e-12
C105_144 V105 V144 3.552598773616155e-20

R106_106 V106 0 401.78279948076363
L106_106 V106 0 -2.2363486145941614e-13
C106_106 V106 0 -1.5209423883675023e-19

R106_107 V106 V107 -1089.7449052376505
L106_107 V106 V107 -3.132913754189523e-13
C106_107 V106 V107 -2.144896239840476e-18

R106_108 V106 V108 -93074.86685237239
L106_108 V106 V108 3.38634419831565e-13
C106_108 V106 V108 2.055552148072592e-18

R106_109 V106 V109 -4400.096439844528
L106_109 V106 V109 1.2530866728094395e-12
C106_109 V106 V109 4.2058578195114135e-19

R106_110 V106 V110 1642.9047000999722
L106_110 V106 V110 2.508313105030047e-13
C106_110 V106 V110 3.0294960220490432e-18

R106_111 V106 V111 6260.468973646704
L106_111 V106 V111 3.7737864634631903e-13
C106_111 V106 V111 1.4177523481766098e-18

R106_112 V106 V112 -519.9685555437829
L106_112 V106 V112 -3.6404849427988546e-13
C106_112 V106 V112 -1.9470188421312163e-18

R106_113 V106 V113 -1191.262316254971
L106_113 V106 V113 -7.018904873794548e-13
C106_113 V106 V113 -8.538904062210604e-19

R106_114 V106 V114 -1288.4755533963223
L106_114 V106 V114 -4.190511266404649e-13
C106_114 V106 V114 -1.745929812863271e-18

R106_115 V106 V115 -2059.911316389497
L106_115 V106 V115 -5.295494338629127e-13
C106_115 V106 V115 -1.148129111672157e-18

R106_116 V106 V116 1577.674922611499
L106_116 V106 V116 4.941853692659836e-13
C106_116 V106 V116 1.2353248258520203e-18

R106_117 V106 V117 3644.3488720426562
L106_117 V106 V117 7.98083201070872e-13
C106_117 V106 V117 1.048884654194511e-18

R106_118 V106 V118 1232.377702376754
L106_118 V106 V118 4.4083852979246654e-13
C106_118 V106 V118 1.4957048355533966e-18

R106_119 V106 V119 3504.1920895206886
L106_119 V106 V119 3.163440994729737e-13
C106_119 V106 V119 1.989829279885634e-18

R106_120 V106 V120 33032.844460187145
L106_120 V106 V120 -1.3107556152319605e-12
C106_120 V106 V120 5.785554590826404e-19

R106_121 V106 V121 -502.4559582040968
L106_121 V106 V121 -2.337856818424516e-12
C106_121 V106 V121 -3.919683314717603e-19

R106_122 V106 V122 -305.5626935699395
L106_122 V106 V122 -8.33750817700729e-13
C106_122 V106 V122 -5.927543089308783e-20

R106_123 V106 V123 -1624.983131253282
L106_123 V106 V123 2.648155927936675e-12
C106_123 V106 V123 2.7804807271654723e-19

R106_124 V106 V124 -8012.563537694962
L106_124 V106 V124 9.896684945416174e-13
C106_124 V106 V124 4.944353300914671e-19

R106_125 V106 V125 554.8833090133093
L106_125 V106 V125 -8.04616200896411e-12
C106_125 V106 V125 3.315092589651105e-19

R106_126 V106 V126 385.6594274704363
L106_126 V106 V126 6.399376394014111e-13
C106_126 V106 V126 -3.3502428865876273e-19

R106_127 V106 V127 -686.9738740781371
L106_127 V106 V127 -5.302510741022796e-13
C106_127 V106 V127 -1.4058821279790154e-20

R106_128 V106 V128 52388.85677407857
L106_128 V106 V128 -6.622290182046362e-12
C106_128 V106 V128 1.8882810813322165e-19

R106_129 V106 V129 -1363.0207821744748
L106_129 V106 V129 -4.314639129957926e-12
C106_129 V106 V129 1.9297972476187377e-19

R106_130 V106 V130 948.6081145608177
L106_130 V106 V130 1.008257137650594e-12
C106_130 V106 V130 7.447597378396465e-19

R106_131 V106 V131 1118.9132191621763
L106_131 V106 V131 -1.5104862400865231e-12
C106_131 V106 V131 -5.057872655834369e-19

R106_132 V106 V132 1791.153028563419
L106_132 V106 V132 2.108518046554798e-12
C106_132 V106 V132 6.294256461629631e-20

R106_133 V106 V133 3680.0451211434774
L106_133 V106 V133 -5.517560723524374e-13
C106_133 V106 V133 -1.1950483886801409e-18

R106_134 V106 V134 1818.075413623453
L106_134 V106 V134 5.901016660591829e-12
C106_134 V106 V134 4.63719729539689e-20

R106_135 V106 V135 -956.6189381977989
L106_135 V106 V135 -1.142133553381762e-12
C106_135 V106 V135 1.9602085279775234e-19

R106_136 V106 V136 5067.973576078986
L106_136 V106 V136 -3.423169867020582e-12
C106_136 V106 V136 -3.361212137971228e-20

R106_137 V106 V137 838.770155356871
L106_137 V106 V137 2.8406857130421846e-12
C106_137 V106 V137 5.695586676208436e-19

R106_138 V106 V138 372.6149428486404
L106_138 V106 V138 7.353175176773108e-13
C106_138 V106 V138 1.2538969133621616e-19

R106_139 V106 V139 -501.8526812667598
L106_139 V106 V139 -3.793512100407691e-13
C106_139 V106 V139 -4.026417973120249e-19

R106_140 V106 V140 1096.3145138281523
L106_140 V106 V140 1.2630337920993141e-12
C106_140 V106 V140 1.8594305767748635e-19

R106_141 V106 V141 1674.3196513992211
L106_141 V106 V141 1.6892998227713452e-12
C106_141 V106 V141 7.685219041210798e-20

R106_142 V106 V142 1050.75415768145
L106_142 V106 V142 1.1278499958688753e-12
C106_142 V106 V142 3.1033435121636344e-19

R106_143 V106 V143 1849.5120013988615
L106_143 V106 V143 1.4302983752423398e-12
C106_143 V106 V143 4.7484536491056285e-20

R106_144 V106 V144 -1391.3853256983332
L106_144 V106 V144 -1.7908114869124198e-12
C106_144 V106 V144 -1.4280373773655747e-19

R107_107 V107 0 593.4836215919837
L107_107 V107 0 -2.7438437615204927e-13
C107_107 V107 0 -9.718542352174429e-19

R107_108 V107 V108 1156.2096041933228
L107_108 V107 V108 3.020671813192234e-13
C107_108 V107 V108 1.9895275449227926e-18

R107_109 V107 V109 1660.8533770755644
L107_109 V107 V109 6.39974442412306e-13
C107_109 V107 V109 9.167444548190247e-19

R107_110 V107 V110 11531.698705510598
L107_110 V107 V110 6.241240607763761e-13
C107_110 V107 V110 1.378043064996206e-18

R107_111 V107 V111 878.7204407440853
L107_111 V107 V111 3.95672331508105e-13
C107_111 V107 V111 1.3432152574701216e-18

R107_112 V107 V112 -2219.215813290199
L107_112 V107 V112 -3.173356374014218e-13
C107_112 V107 V112 -1.6211441984666523e-18

R107_113 V107 V113 -2559.6333830381295
L107_113 V107 V113 -6.633050125821045e-13
C107_113 V107 V113 -7.192026755268145e-19

R107_114 V107 V114 -3269.134372305529
L107_114 V107 V114 -6.572043323137555e-13
C107_114 V107 V114 -7.952877328833571e-19

R107_115 V107 V115 -1227.1825213105205
L107_115 V107 V115 -4.1502844877382466e-13
C107_115 V107 V115 -1.5228233306988916e-18

R107_116 V107 V116 1696.6443443078144
L107_116 V107 V116 4.49478392492985e-13
C107_116 V107 V116 1.1321428033588415e-18

R107_117 V107 V117 10314.397190303727
L107_117 V107 V117 8.770609118565007e-13
C107_117 V107 V117 9.497668234181747e-19

R107_118 V107 V118 2992.90830041417
L107_118 V107 V118 6.401518103368779e-13
C107_118 V107 V118 8.123685604416719e-19

R107_119 V107 V119 1216.7347568275316
L107_119 V107 V119 4.956789241191448e-13
C107_119 V107 V119 9.507186588357209e-19

R107_120 V107 V120 -715.0594649488403
L107_120 V107 V120 -6.617422818266809e-13
C107_120 V107 V120 4.197331091900641e-19

R107_121 V107 V121 1579.9120620993924
L107_121 V107 V121 -1.9853546240579334e-12
C107_121 V107 V121 -2.5808416350509513e-19

R107_122 V107 V122 -1600.4065372142536
L107_122 V107 V122 -3.80912141070746e-13
C107_122 V107 V122 8.523015446189263e-20

R107_123 V107 V123 -80992.74398958492
L107_123 V107 V123 -2.501830501469878e-12
C107_123 V107 V123 1.5328378978625885e-19

R107_124 V107 V124 2325.517748508449
L107_124 V107 V124 1.6079301479238222e-12
C107_124 V107 V124 2.8634222213313695e-19

R107_125 V107 V125 -914.9292570656723
L107_125 V107 V125 -1.3358287744328667e-11
C107_125 V107 V125 2.2590004512307993e-19

R107_126 V107 V126 672.6745732378375
L107_126 V107 V126 3.0286545171554285e-13
C107_126 V107 V126 -2.5650375609714984e-19

R107_127 V107 V127 -662.6731630297057
L107_127 V107 V127 -3.42584335190469e-13
C107_127 V107 V127 -4.6451759414613675e-20

R107_128 V107 V128 -4431.63996260088
L107_128 V107 V128 -4.730011662312441e-12
C107_128 V107 V128 4.877823761022118e-20

R107_129 V107 V129 -2951.2949913572284
L107_129 V107 V129 -1.0184965664378218e-12
C107_129 V107 V129 2.780956955539193e-20

R107_130 V107 V130 2481.3194398251653
L107_130 V107 V130 5.395564967061383e-13
C107_130 V107 V130 6.63725835919685e-19

R107_131 V107 V131 -7981.249096747109
L107_131 V107 V131 -1.338016952424636e-11
C107_131 V107 V131 -6.618745791121892e-19

R107_132 V107 V132 3265.781089954771
L107_132 V107 V132 1.2375053457805618e-12
C107_132 V107 V132 5.481062401483941e-20

R107_133 V107 V133 -2470.4852544126634
L107_133 V107 V133 -1.3905322801912145e-12
C107_133 V107 V133 -5.235927321347387e-19

R107_134 V107 V134 13487.94503115139
L107_134 V107 V134 2.5756648708866246e-12
C107_134 V107 V134 -8.604334691477702e-20

R107_135 V107 V135 -1164.3084898259845
L107_135 V107 V135 -6.374434737328951e-13
C107_135 V107 V135 3.2289629460189786e-19

R107_136 V107 V136 -6030.137335846848
L107_136 V107 V136 -2.8989958455493948e-11
C107_136 V107 V136 1.6830071637521283e-20

R107_137 V107 V137 -2160.0453162918398
L107_137 V107 V137 3.707239101718665e-12
C107_137 V107 V137 2.268513624760317e-19

R107_138 V107 V138 845.2450128090142
L107_138 V107 V138 3.125431788587819e-13
C107_138 V107 V138 1.760660353179858e-19

R107_139 V107 V139 -483.6315050170972
L107_139 V107 V139 -2.4720213914425544e-13
C107_139 V107 V139 -3.768499351781731e-19

R107_140 V107 V140 2933.627360085198
L107_140 V107 V140 7.214027663691805e-13
C107_140 V107 V140 1.6896360980269873e-19

R107_141 V107 V141 2632.8348686157074
L107_141 V107 V141 1.2579541158255892e-12
C107_141 V107 V141 9.808190363680954e-20

R107_142 V107 V142 2899.8374099845346
L107_142 V107 V142 6.693964670910764e-13
C107_142 V107 V142 2.577071158217451e-19

R107_143 V107 V143 1464.116909034656
L107_143 V107 V143 7.44487247407141e-13
C107_143 V107 V143 7.561059915233281e-20

R107_144 V107 V144 -9434.292658408682
L107_144 V107 V144 -9.936589180480074e-13
C107_144 V107 V144 -1.5508218655962862e-19

R108_108 V108 0 -640.7529179875007
L108_108 V108 0 1.9883108543396707e-13
C108_108 V108 0 7.834093223753015e-19

R108_109 V108 V109 3788.4254200913792
L108_109 V108 V109 -1.7751013513819978e-12
C108_109 V108 V109 -3.546102004344488e-19

R108_110 V108 V110 12477.329433188788
L108_110 V108 V110 -4.908079870687116e-13
C108_110 V108 V110 -1.564761533403124e-18

R108_111 V108 V111 -4741.991552539593
L108_111 V108 V111 -5.206464983400431e-13
C108_111 V108 V111 -1.0768240400220204e-18

R108_112 V108 V112 404.56567966779346
L108_112 V108 V112 2.887111019708964e-13
C108_112 V108 V112 1.949364924874979e-18

R108_113 V108 V113 874.6298146378655
L108_113 V108 V113 7.593286177693836e-13
C108_113 V108 V113 5.760275944837757e-19

R108_114 V108 V114 2251.8613790262893
L108_114 V108 V114 7.326372625183179e-13
C108_114 V108 V114 9.028173519737643e-19

R108_115 V108 V115 1798.1025509811657
L108_115 V108 V115 5.758032882972737e-13
C108_115 V108 V115 1.1142511447696155e-18

R108_116 V108 V116 -1165.576637542545
L108_116 V108 V116 -4.1472791893570316e-13
C108_116 V108 V116 -1.4909315456739466e-18

R108_117 V108 V117 -4905.82234575322
L108_117 V108 V117 -8.725905662671769e-13
C108_117 V108 V117 -9.950445335710697e-19

R108_118 V108 V118 -1339.3361891555548
L108_118 V108 V118 -6.985620379591085e-13
C108_118 V108 V118 -6.504911560782584e-19

R108_119 V108 V119 -11554.770775469373
L108_119 V108 V119 -5.438510812907509e-13
C108_119 V108 V119 -1.1562259635686593e-18

R108_120 V108 V120 1483.1833900652314
L108_120 V108 V120 2.184383555705104e-12
C108_120 V108 V120 -6.037150344477218e-19

R108_121 V108 V121 458.0151311545499
L108_121 V108 V121 1.1084178736943952e-12
C108_121 V108 V121 6.274657654807268e-20

R108_122 V108 V122 215.6743819038185
L108_122 V108 V122 4.296023441837826e-13
C108_122 V108 V122 4.156262345495276e-20

R108_123 V108 V123 1313.1172024512357
L108_123 V108 V123 5.901778223058187e-12
C108_123 V108 V123 -9.114548362692724e-20

R108_124 V108 V124 -9049.713995222886
L108_124 V108 V124 -1.3984900719359274e-12
C108_124 V108 V124 -4.040857531698981e-19

R108_125 V108 V125 -523.3050283648776
L108_125 V108 V125 -1.1698869946510807e-12
C108_125 V108 V125 -2.8127803405365864e-19

R108_126 V108 V126 -241.22432179936285
L108_126 V108 V126 -4.1439661103450146e-13
C108_126 V108 V126 2.087593198761166e-19

R108_127 V108 V127 377.5957212013984
L108_127 V108 V127 4.869094405701198e-13
C108_127 V108 V127 -1.2325636740570174e-20

R108_128 V108 V128 3654.2743612267077
L108_128 V108 V128 5.087290288268261e-12
C108_128 V108 V128 -1.8815193933872938e-20

R108_129 V108 V129 1143.6181826824552
L108_129 V108 V129 2.551577445626953e-12
C108_129 V108 V129 -1.5074905186203223e-19

R108_130 V108 V130 -1078.4312944058183
L108_130 V108 V130 -7.400619628947189e-13
C108_130 V108 V130 -7.034769786684689e-19

R108_131 V108 V131 -1026.066014089024
L108_131 V108 V131 4.117678834106769e-12
C108_131 V108 V131 4.806232230526536e-19

R108_132 V108 V132 -1127.2676416854767
L108_132 V108 V132 -1.2809797794361572e-12
C108_132 V108 V132 -1.8973420192909794e-19

R108_133 V108 V133 -2034.597034351385
L108_133 V108 V133 1.4625472946378925e-12
C108_133 V108 V133 5.434133461630379e-19

R108_134 V108 V134 -1146.7734459844887
L108_134 V108 V134 -2.684917663142552e-12
C108_134 V108 V134 1.0148907179640132e-19

R108_135 V108 V135 537.8070975375804
L108_135 V108 V135 9.251750541155094e-13
C108_135 V108 V135 -2.739748724318411e-19

R108_136 V108 V136 -13561.091410298432
L108_136 V108 V136 1.010993207838535e-11
C108_136 V108 V136 2.172446173118467e-20

R108_137 V108 V137 -763.5246129683486
L108_137 V108 V137 -1.3841746086848267e-12
C108_137 V108 V137 -3.58808206432293e-19

R108_138 V108 V138 -258.4781273168577
L108_138 V108 V138 -4.480632091595369e-13
C108_138 V108 V138 -1.8232787101909144e-19

R108_139 V108 V139 288.9686571225979
L108_139 V108 V139 3.4654724781824873e-13
C108_139 V108 V139 2.7277184170341736e-19

R108_140 V108 V140 -769.849862950693
L108_140 V108 V140 -7.89403194212219e-13
C108_140 V108 V140 -2.2870153027167377e-19

R108_141 V108 V141 -948.0512660038493
L108_141 V108 V141 -1.2869590387976576e-12
C108_141 V108 V141 -7.486207178546928e-20

R108_142 V108 V142 -1017.6113058537691
L108_142 V108 V142 -1.111486214456291e-12
C108_142 V108 V142 -2.615534470695297e-19

R108_143 V108 V143 -1111.0634110165984
L108_143 V108 V143 -1.1690740772355288e-12
C108_143 V108 V143 -9.806421194767005e-20

R108_144 V108 V144 1049.6034201415794
L108_144 V108 V144 1.1978583547064886e-12
C108_144 V108 V144 1.2879269191222815e-19

R109_109 V109 0 1379.068787655916
L109_109 V109 0 -1.442445502639998e-12
C109_109 V109 0 -5.869203523324992e-20

R109_110 V109 V110 -5742.886023084308
L109_110 V109 V110 -5.298786176223715e-12
C109_110 V109 V110 -3.1425314616086416e-19

R109_111 V109 V111 2842.8346753993274
L109_111 V109 V111 -1.2545873471608795e-12
C109_111 V109 V111 -2.2545503455523583e-19

R109_112 V109 V112 983.4681133249294
L109_112 V109 V112 1.2845376000451324e-12
C109_112 V109 V112 5.113871889338106e-19

R109_113 V109 V113 1390.1569437228964
L109_113 V109 V113 1.0431553894113619e-12
C109_113 V109 V113 6.426757050497326e-19

R109_114 V109 V114 -5489.808445292497
L109_114 V109 V114 2.8046165996300385e-12
C109_114 V109 V114 1.7381425563920821e-19

R109_115 V109 V115 20855.267584000463
L109_115 V109 V115 1.1623152114610415e-12
C109_115 V109 V115 4.242831297663467e-19

R109_116 V109 V116 -6647.422805079385
L109_116 V109 V116 -2.5067481614244876e-12
C109_116 V109 V116 -1.4572592221671925e-19

R109_117 V109 V117 -3068.9672695268027
L109_117 V109 V117 -2.198265576344741e-12
C109_117 V109 V117 -6.181350936321481e-19

R109_118 V109 V118 -2791.649755212183
L109_118 V109 V118 -1.2335695913844217e-12
C109_118 V109 V118 -5.025446662732353e-19

R109_119 V109 V119 1843.7915596413852
L109_119 V109 V119 -3.1783464405439928e-12
C109_119 V109 V119 6.811624029748297e-20

R109_120 V109 V120 -1453.3412474782565
L109_120 V109 V120 8.300379492475387e-13
C109_120 V109 V120 1.4917914756167204e-19

R109_121 V109 V121 705.1748010538028
L109_121 V109 V121 7.909505355261396e-12
C109_121 V109 V121 6.954638448867846e-20

R109_122 V109 V122 759.1337247889188
L109_122 V109 V122 1.0415472554295392e-12
C109_122 V109 V122 -6.325017184844546e-20

R109_123 V109 V123 -15636.103931491843
L109_123 V109 V123 9.763196826659328e-12
C109_123 V109 V123 -1.1362671043253098e-19

R109_124 V109 V124 25587.574504435033
L109_124 V109 V124 -7.454394447978555e-11
C109_124 V109 V124 2.758030482495837e-19

R109_125 V109 V125 -597.4102958496063
L109_125 V109 V125 3.0251944082499792e-12
C109_125 V109 V125 -8.840354554753794e-20

R109_126 V109 V126 -1870.445059400878
L109_126 V109 V126 -6.595297385248364e-13
C109_126 V109 V126 9.744241229695979e-20

R109_127 V109 V127 9048.872186653161
L109_127 V109 V127 7.37830978134102e-13
C109_127 V109 V127 8.892869167229961e-20

R109_128 V109 V128 7909.251401868986
L109_128 V109 V128 3.427872117911423e-12
C109_128 V109 V128 -7.60091443774644e-21

R109_129 V109 V129 -4171.342199624756
L109_129 V109 V129 2.064797761765156e-12
C109_129 V109 V129 2.986473868394794e-20

R109_130 V109 V130 4995.479713603133
L109_130 V109 V130 -1.860848414040526e-12
C109_130 V109 V130 -1.990714780789444e-19

R109_131 V109 V131 8650.671543148886
L109_131 V109 V131 1.2776040350993055e-11
C109_131 V109 V131 2.1882404986596153e-19

R109_132 V109 V132 -6345.593442574112
L109_132 V109 V132 -2.575699822716667e-10
C109_132 V109 V132 2.3679199653445067e-19

R109_133 V109 V133 -3797.140756630414
L109_133 V109 V133 9.72622696602994e-12
C109_133 V109 V133 2.9577866418130737e-20

R109_134 V109 V134 -3352.303738172504
L109_134 V109 V134 -1.1525832517625299e-11
C109_134 V109 V134 6.336659629673673e-20

R109_135 V109 V135 9838.352789380451
L109_135 V109 V135 1.2997739131798349e-12
C109_135 V109 V135 -7.11776669275856e-20

R109_136 V109 V136 49784.59588337634
L109_136 V109 V136 -2.8787827373997947e-11
C109_136 V109 V136 -9.863681245452583e-20

R109_137 V109 V137 -1044.3650795228093
L109_137 V109 V137 8.684085347657877e-12
C109_137 V109 V137 4.2631245208951503e-20

R109_138 V109 V138 -2115.338473659082
L109_138 V109 V138 -7.149203380969249e-13
C109_138 V109 V138 -4.498675951468295e-20

R109_139 V109 V139 8663.627795557342
L109_139 V109 V139 5.640749077327094e-13
C109_139 V109 V139 7.927509241557188e-20

R109_140 V109 V140 -3856.4145466614914
L109_140 V109 V140 -2.113604292940109e-12
C109_140 V109 V140 -6.585958940022958e-20

R109_141 V109 V141 -2563.223919640643
L109_141 V109 V141 -2.086906078256609e-12
C109_141 V109 V141 -1.1063140615415368e-19

R109_142 V109 V142 4353.892331529497
L109_142 V109 V142 -1.6822410283273814e-12
C109_142 V109 V142 -4.464526821794629e-20

R109_143 V109 V143 4753.432927111287
L109_143 V109 V143 -1.6135605293135534e-12
C109_143 V109 V143 9.903961916212003e-21

R109_144 V109 V144 3015.532157954642
L109_144 V109 V144 3.58967553951701e-12
C109_144 V109 V144 8.583649748476176e-20

R110_110 V110 0 -123.02675104714424
L110_110 V110 0 1.660662567910417e-13
C110_110 V110 0 6.914926994809222e-19

R110_111 V110 V111 -615.0358219435549
L110_111 V110 V111 -8.204377994273323e-13
C110_111 V110 V111 -1.058078146840199e-18

R110_112 V110 V112 555.8990896473836
L110_112 V110 V112 3.9211866501209783e-13
C110_112 V110 V112 1.4529333320001144e-18

R110_113 V110 V113 803.7272219616617
L110_113 V110 V113 8.441128897694415e-13
C110_113 V110 V113 6.684707088143985e-19

R110_114 V110 V114 985.6534879848725
L110_114 V110 V114 4.956738647493544e-13
C110_114 V110 V114 1.5936517557366877e-18

R110_115 V110 V115 1062.187486311922
L110_115 V110 V115 1.4458033782137286e-12
C110_115 V110 V115 6.909971973782033e-19

R110_116 V110 V116 -1014.0229272148442
L110_116 V110 V116 -5.9287408625737e-13
C110_116 V110 V116 -1.0274529686184903e-18

R110_117 V110 V117 1624.4729873776282
L110_117 V110 V117 -8.601496925869422e-13
C110_117 V110 V117 -7.965859366741861e-19

R110_118 V110 V118 -1089.3888398132185
L110_118 V110 V118 -5.137438420006108e-13
C110_118 V110 V118 -1.3024195140382253e-18

R110_119 V110 V119 -651.606510513768
L110_119 V110 V119 -4.647325793006544e-13
C110_119 V110 V119 -1.693562582213112e-18

R110_120 V110 V120 217.92030988781227
L110_120 V110 V120 -1.6373122527839988e-12
C110_120 V110 V120 -4.64870014085523e-19

R110_121 V110 V121 2480.0444935959254
L110_121 V110 V121 8.350160808383096e-13
C110_121 V110 V121 3.1841856775532155e-19

R110_122 V110 V122 156.5344350928265
L110_122 V110 V122 1.012002959352216e-12
C110_122 V110 V122 2.4794220883360918e-20

R110_123 V110 V123 857.489751259228
L110_123 V110 V123 -1.827130800499891e-12
C110_123 V110 V123 -3.3064169483582215e-19

R110_124 V110 V124 -1589.5506333585834
L110_124 V110 V124 -1.4807722285732278e-12
C110_124 V110 V124 -4.367606993497207e-19

R110_125 V110 V125 875.4456582406497
L110_125 V110 V125 -7.868668444818868e-13
C110_125 V110 V125 -3.097587275674633e-19

R110_126 V110 V126 -121.29176640947101
L110_126 V110 V126 -1.785306821283171e-12
C110_126 V110 V126 1.868034798183864e-19

R110_127 V110 V127 158.07018464423973
L110_127 V110 V127 1.820256079236473e-12
C110_127 V110 V127 4.269288380846754e-22

R110_128 V110 V128 1534.0594366406456
L110_128 V110 V128 5.93487197451224e-11
C110_128 V110 V128 -1.7599233860280284e-19

R110_129 V110 V129 454.7743741575345
L110_129 V110 V129 -2.5976127436914637e-12
C110_129 V110 V129 -2.1619201683056344e-19

R110_130 V110 V130 -562.8309848196141
L110_130 V110 V130 -3.261272751298087e-12
C110_130 V110 V130 -4.913494224570693e-19

R110_131 V110 V131 -522.7869061282794
L110_131 V110 V131 2.195913682642936e-12
C110_131 V110 V131 3.226861934032756e-19

R110_132 V110 V132 -632.6241188495125
L110_132 V110 V132 -3.1020661172899817e-12
C110_132 V110 V132 -7.198612777758031e-20

R110_133 V110 V133 -23801.827543314634
L110_133 V110 V133 9.975847194843599e-13
C110_133 V110 V133 8.534646221211662e-19

R110_134 V110 V134 -878.131884510415
L110_134 V110 V134 -8.50793424016984e-12
C110_134 V110 V134 -1.3016778653710961e-20

R110_135 V110 V135 233.37989952708747
L110_135 V110 V135 8.425978033213932e-12
C110_135 V110 V135 -1.6600057026462694e-19

R110_136 V110 V136 5503.49846075681
L110_136 V110 V136 6.4464656664674006e-12
C110_136 V110 V136 3.3428401863187924e-20

R110_137 V110 V137 7212.583902740247
L110_137 V110 V137 -1.1431015651821028e-12
C110_137 V110 V137 -4.072505866005463e-19

R110_138 V110 V138 -143.84513565542684
L110_138 V110 V138 -2.058339224254041e-12
C110_138 V110 V138 -1.365451405387071e-19

R110_139 V110 V139 121.44598860649529
L110_139 V110 V139 1.2720316429187183e-12
C110_139 V110 V139 2.4424826705653725e-19

R110_140 V110 V140 -493.7125466637611
L110_140 V110 V140 -2.0963987873876104e-12
C110_140 V110 V140 -9.917547859582973e-20

R110_141 V110 V141 -600.4604964775874
L110_141 V110 V141 -2.3774912367502243e-12
C110_141 V110 V141 -7.18807966047971e-20

R110_142 V110 V142 -470.81846104230544
L110_142 V110 V142 -1.9785098095056612e-12
C110_142 V110 V142 -3.372186195469095e-19

R110_143 V110 V143 -378.13383214801775
L110_143 V110 V143 -7.170822823200932e-12
C110_143 V110 V143 -1.1389103428129762e-19

R110_144 V110 V144 901.9567454182325
L110_144 V110 V144 2.519029242213738e-12
C110_144 V110 V144 1.1410700706061612e-19

R111_111 V111 0 119.14046778802242
L111_111 V111 0 3.6873904234840395e-13
C111_111 V111 0 1.2710437534446685e-18

R111_112 V111 V112 2672.7467586341195
L111_112 V111 V112 1.0169492089199588e-12
C111_112 V111 V112 9.071657881258515e-19

R111_113 V111 V113 10316.471495663864
L111_113 V111 V113 2.1572836621566162e-12
C111_113 V111 V113 3.051438885563491e-19

R111_114 V111 V114 -1864.0154198857488
L111_114 V111 V114 1.1824339324251166e-12
C111_114 V111 V114 6.640015780563817e-19

R111_115 V111 V115 -2436.634279385773
L111_115 V111 V115 6.937285957269996e-13
C111_115 V111 V115 6.767620874776908e-19

R111_116 V111 V116 4094.853118947714
L111_116 V111 V116 -8.053010000094394e-13
C111_116 V111 V116 -6.420417159476969e-19

R111_117 V111 V117 -995.2708471270543
L111_117 V111 V117 -3.821087667665392e-12
C111_117 V111 V117 -4.021533600022009e-19

R111_118 V111 V118 -6467.503099521733
L111_118 V111 V118 -1.2581496071224003e-12
C111_118 V111 V118 -4.733599726628839e-19

R111_119 V111 V119 728.3181390194263
L111_119 V111 V119 -5.777118498029272e-13
C111_119 V111 V119 -7.575020537128121e-19

R111_120 V111 V120 -217.1259459456322
L111_120 V111 V120 6.55248902902176e-13
C111_120 V111 V120 -2.9808889929700266e-19

R111_121 V111 V121 555.1062509851114
L111_121 V111 V121 -1.6466944298385739e-12
C111_121 V111 V121 1.8658724897638797e-19

R111_122 V111 V122 -352.9470411190333
L111_122 V111 V122 4.916476128202125e-12
C111_122 V111 V122 -6.228672566540968e-20

R111_123 V111 V123 -1039.387991271728
L111_123 V111 V123 -2.8598444891213288e-12
C111_123 V111 V123 -1.3580182919055717e-19

R111_124 V111 V124 -63513.36207257276
L111_124 V111 V124 -1.2748529432340995e-12
C111_124 V111 V124 -2.5921084922719376e-19

R111_125 V111 V125 -308.7626031431965
L111_125 V111 V125 8.854212950105792e-13
C111_125 V111 V125 -1.6242591133660924e-19

R111_126 V111 V126 184.51492624789742
L111_126 V111 V126 -6.575269163914446e-13
C111_126 V111 V126 1.161286664466086e-19

R111_127 V111 V127 -217.4676891115384
L111_127 V111 V127 5.585429111243918e-13
C111_127 V111 V127 2.1768055559199675e-21

R111_128 V111 V128 -34250.18592728585
L111_128 V111 V128 8.143330973326202e-12
C111_128 V111 V128 -2.2201444774204767e-20

R111_129 V111 V129 -477.3603489578406
L111_129 V111 V129 3.3269580804675103e-12
C111_129 V111 V129 -4.0645500406783134e-20

R111_130 V111 V130 646.6145480451729
L111_130 V111 V130 -1.866610310753815e-12
C111_130 V111 V130 -3.1893644729994056e-19

R111_131 V111 V131 581.3009408546474
L111_131 V111 V131 1.4791241396015376e-12
C111_131 V111 V131 3.3593295012977228e-19

R111_132 V111 V132 1023.8672092647664
L111_132 V111 V132 -2.834134134902093e-12
C111_132 V111 V132 -5.91659744935948e-20

R111_133 V111 V133 -14760.730788623761
L111_133 V111 V133 1.1481183862875316e-12
C111_133 V111 V133 3.3436120603930936e-19

R111_134 V111 V134 2533.73453869951
L111_134 V111 V134 -4.7855604158505963e-11
C111_134 V111 V134 1.1357820676297025e-20

R111_135 V111 V135 -321.6157489630624
L111_135 V111 V135 1.1490680424504901e-12
C111_135 V111 V135 -1.727345759679937e-19

R111_136 V111 V136 236619.49303831183
L111_136 V111 V136 6.724665646309171e-12
C111_136 V111 V136 -1.0394906392243471e-22

R111_137 V111 V137 -616.9827092905673
L111_137 V111 V137 1.7589047208996e-12
C111_137 V111 V137 -1.4857647144453122e-19

R111_138 V111 V138 226.39557775812983
L111_138 V111 V138 -9.670018050048125e-13
C111_138 V111 V138 -1.2544610573396665e-19

R111_139 V111 V139 -171.2343225818569
L111_139 V111 V139 4.039233764958264e-13
C111_139 V111 V139 2.1086392938873443e-19

R111_140 V111 V140 784.1196737414517
L111_140 V111 V140 -1.8376126214170225e-12
C111_140 V111 V140 -9.604548640943538e-20

R111_141 V111 V141 2190.392889145243
L111_141 V111 V141 -2.1471835678781815e-12
C111_141 V111 V141 -7.542462678965242e-20

R111_142 V111 V142 539.3334983823836
L111_142 V111 V142 -2.0817494988128575e-12
C111_142 V111 V142 -2.1675168502748562e-19

R111_143 V111 V143 440.79555685519205
L111_143 V111 V143 -1.2462701674600454e-12
C111_143 V111 V143 -1.849288230279702e-20

R111_144 V111 V144 -2392.3851686067183
L111_144 V111 V144 4.683164553035404e-12
C111_144 V111 V144 -8.87944495099526e-21

R112_112 V112 0 -391.7864072857301
L112_112 V112 0 -1.6663663631505884e-13
C112_112 V112 0 3.2093650804095344e-20

R112_113 V112 V113 995.6657480620814
L112_113 V112 V113 -5.497545947351771e-13
C112_113 V112 V113 -5.564820906897676e-19

R112_114 V112 V114 -3366.9002866156593
L112_114 V112 V114 -5.182770709372908e-13
C112_114 V112 V114 -9.18715673507288e-19

R112_115 V112 V115 -9361.528477825475
L112_115 V112 V115 -6.498820842883481e-13
C112_115 V112 V115 -9.167860829235558e-19

R112_116 V112 V116 -29104.09038801087
L112_116 V112 V116 3.9155658525163575e-13
C112_116 V112 V116 1.0482627385258091e-18

R112_117 V112 V117 972.8522544016779
L112_117 V112 V117 5.66764834672067e-13
C112_117 V112 V117 8.392118061298458e-19

R112_118 V112 V118 -2296.0159154960147
L112_118 V112 V118 5.426062120922645e-13
C112_118 V112 V118 6.343581515153178e-19

R112_119 V112 V119 1286.561365765996
L112_119 V112 V119 6.460444957035509e-13
C112_119 V112 V119 1.047546410996481e-18

R112_120 V112 V120 474.4505330158753
L112_120 V112 V120 1.4618533078826297e-12
C112_120 V112 V120 4.723081499835516e-19

R112_121 V112 V121 296.9492806600537
L112_121 V112 V121 -3.7696927571608304e-13
C112_121 V112 V121 -1.0625216807798544e-19

R112_122 V112 V122 133.01413370890728
L112_122 V112 V122 -2.355122697522754e-13
C112_122 V112 V122 -6.749056666238896e-20

R112_123 V112 V123 882.7201613126318
L112_123 V112 V123 -1.5636625475507922e-12
C112_123 V112 V123 9.27968273456738e-20

R112_124 V112 V124 4452.728979294351
L112_124 V112 V124 -5.065032376867164e-12
C112_124 V112 V124 2.699115483721552e-19

R112_125 V112 V125 -385.82531047989943
L112_125 V112 V125 3.622024653899104e-13
C112_125 V112 V125 1.4074603974456537e-19

R112_126 V112 V126 -134.10407753065172
L112_126 V112 V126 3.57390689874557e-13
C112_126 V112 V126 -2.5693443283139675e-19

R112_127 V112 V127 210.44675327293956
L112_127 V112 V127 -5.267920530993502e-13
C112_127 V112 V127 1.9687014570577278e-20

R112_128 V112 V128 5987.791149028518
L112_128 V112 V128 3.72303855379482e-12
C112_128 V112 V128 1.145349051439943e-21

R112_129 V112 V129 603.8516396924343
L112_129 V112 V129 -2.011143099142426e-12
C112_129 V112 V129 1.8569812050000253e-19

R112_130 V112 V130 -1215.2366366848632
L112_130 V112 V130 5.07034930107932e-13
C112_130 V112 V130 5.548882688919466e-19

R112_131 V112 V131 -486.54884055673585
L112_131 V112 V131 2.6865445871391697e-12
C112_131 V112 V131 -4.670332450377192e-19

R112_132 V112 V132 -689.4823762079329
L112_132 V112 V132 1.2292752266091226e-12
C112_132 V112 V132 5.3819766856088717e-20

R112_133 V112 V133 -754.277679269321
L112_133 V112 V133 -4.219834895950042e-12
C112_133 V112 V133 -5.787023666505751e-19

R112_134 V112 V134 -666.3494440670587
L112_134 V112 V134 1.5779331775795974e-12
C112_134 V112 V134 -1.018450181548928e-19

R112_135 V112 V135 285.14206473045465
L112_135 V112 V135 -8.326360733116058e-13
C112_135 V112 V135 1.7075064900499663e-19

R112_136 V112 V136 -4990.842906786333
L112_136 V112 V136 2.2003966113734417e-12
C112_136 V112 V136 5.3135133314947035e-20

R112_137 V112 V137 -629.5692612116894
L112_137 V112 V137 4.78606810254265e-13
C112_137 V112 V137 4.050030498423526e-19

R112_138 V112 V138 -160.02215814488352
L112_138 V112 V138 2.8829165237343535e-13
C112_138 V112 V138 2.144627315804472e-19

R112_139 V112 V139 168.92594425673144
L112_139 V112 V139 -3.7354293748966324e-13
C112_139 V112 V139 -2.473821300066001e-19

R112_140 V112 V140 -461.59752663861343
L112_140 V112 V140 5.090363176025934e-13
C112_140 V112 V140 2.0167082346327763e-19

R112_141 V112 V141 -640.1720562423345
L112_141 V112 V141 1.4644088737103258e-12
C112_141 V112 V141 1.0150600328145477e-19

R112_142 V112 V142 -752.14040188556
L112_142 V112 V142 6.337339794946495e-13
C112_142 V112 V142 2.5184466114465007e-19

R112_143 V112 V143 -622.3204971573574
L112_143 V112 V143 1.8843236889315527e-12
C112_143 V112 V143 -4.4132328945743646e-20

R112_144 V112 V144 690.4306173811999
L112_144 V112 V144 -6.759807184958841e-13
C112_144 V112 V144 -1.772004837258547e-19

R113_113 V113 0 -1391.5139794605104
L113_113 V113 0 -9.43576773056646e-13
C113_113 V113 0 -1.1139611224986152e-19

R113_114 V113 V114 1146.3658543895065
L113_114 V113 V114 -1.2333343141003738e-12
C113_114 V113 V114 -3.2037364007262975e-19

R113_115 V113 V115 3838.5826306190806
L113_115 V113 V115 -1.382968702822604e-12
C113_115 V113 V115 -3.4697771963964276e-19

R113_116 V113 V116 -15017.927760119066
L113_116 V113 V116 1.0530777588854286e-12
C113_116 V113 V116 2.955692629789956e-19

R113_117 V113 V117 1596.7834508811422
L113_117 V113 V117 9.656539003776553e-13
C113_117 V113 V117 5.52502711870804e-19

R113_118 V113 V118 -3074.1510311775123
L113_118 V113 V118 8.413354205333398e-13
C113_118 V113 V118 5.010641278589665e-19

R113_119 V113 V119 -4697.611925843294
L113_119 V113 V119 1.940664755600447e-12
C113_119 V113 V119 2.6275266168533287e-19

R113_120 V113 V120 592.5230129217997
L113_120 V113 V120 -1.4818430454875532e-11
C113_120 V113 V120 6.039095689279985e-21

R113_121 V113 V121 655.4003844871232
L113_121 V113 V121 -1.0718634847968227e-12
C113_121 V113 V121 -8.182801182171655e-20

R113_122 V113 V122 210.88951574860016
L113_122 V113 V122 -5.677259316932793e-13
C113_122 V113 V122 -2.60879567759331e-21

R113_123 V113 V123 528.794877977992
L113_123 V113 V123 -2.7472315728392393e-12
C113_123 V113 V123 8.575683766992413e-20

R113_124 V113 V124 1702.6594051557145
L113_124 V113 V124 2.1615852334055654e-12
C113_124 V113 V124 -2.0693620347525444e-20

R113_125 V113 V125 -1630.0600538772135
L113_125 V113 V125 1.15434952201298e-12
C113_125 V113 V125 1.0940655878713454e-19

R113_126 V113 V126 -207.47855167706527
L113_126 V113 V126 7.920927871905912e-13
C113_126 V113 V126 -1.1250868101302944e-19

R113_127 V113 V127 333.68390899268644
L113_127 V113 V127 -1.113904291246788e-12
C113_127 V113 V127 -4.662101807567207e-20

R113_128 V113 V128 4464.835289195873
L113_128 V113 V128 -1.5004041618455553e-12
C113_128 V113 V128 9.529253893687929e-20

R113_129 V113 V129 424.9380831394714
L113_129 V113 V129 -5.425568497356647e-12
C113_129 V113 V129 4.4320976659286266e-20

R113_130 V113 V130 -495.566545756536
L113_130 V113 V130 1.3225281592347685e-12
C113_130 V113 V130 2.9430555439764905e-19

R113_131 V113 V131 -400.2687469851739
L113_131 V113 V131 2.3091970375632792e-11
C113_131 V113 V131 -1.6141312035621769e-19

R113_132 V113 V132 -1121.7922388479199
L113_132 V113 V132 3.0328418152137603e-12
C113_132 V113 V132 -4.9280467245212616e-20

R113_133 V113 V133 -1179.2138750776032
L113_133 V113 V133 -2.957322353807796e-12
C113_133 V113 V133 -2.6072420521758793e-19

R113_134 V113 V134 -1177.2626751384082
L113_134 V113 V134 3.4191618126906288e-12
C113_134 V113 V134 -1.359313625525187e-20

R113_135 V113 V135 437.6737409640402
L113_135 V113 V135 -1.826324113333768e-12
C113_135 V113 V135 5.500387649620046e-20

R113_136 V113 V136 -3982.200602806349
L113_136 V113 V136 -2.9411514409591533e-12
C113_136 V113 V136 -1.2527228217743849e-20

R113_137 V113 V137 -2746.4845284840167
L113_137 V113 V137 1.3353767283726444e-12
C113_137 V113 V137 9.07933123682815e-20

R113_138 V113 V138 -200.893417483221
L113_138 V113 V138 7.032537586000924e-13
C113_138 V113 V138 1.2863368968151822e-20

R113_139 V113 V139 261.09434510018895
L113_139 V113 V139 -7.518689731268505e-13
C113_139 V113 V139 -1.0568511284454066e-19

R113_140 V113 V140 -745.3970089953614
L113_140 V113 V140 2.228288796332802e-12
C113_140 V113 V140 8.689232697755045e-20

R113_141 V113 V141 -1688.414676743454
L113_141 V113 V141 1.5965116004503467e-12
C113_141 V113 V141 -5.540177982547214e-21

R113_142 V113 V142 -444.49282010487144
L113_142 V113 V142 1.5553553734578008e-12
C113_142 V113 V142 7.98755199092845e-20

R113_143 V113 V143 -659.1205777689372
L113_143 V113 V143 3.2931211780667663e-12
C113_143 V113 V143 7.781762289537185e-21

R113_144 V113 V144 1295.299053340693
L113_144 V113 V144 -3.098547182055625e-12
C113_144 V113 V144 -2.722856811253139e-20

R114_114 V114 0 -150.4738798111121
L114_114 V114 0 -2.4520633271472696e-13
C114_114 V114 0 -3.1714884003672273e-19

R114_115 V114 V115 -8703.062054937407
L114_115 V114 V115 -1.2249353750971408e-12
C114_115 V114 V115 -3.8300981940572253e-19

R114_116 V114 V116 -77340.68088061658
L114_116 V114 V116 1.0025679349653912e-12
C114_116 V114 V116 5.1838235560988e-19

R114_117 V114 V117 2598.2752604566936
L114_117 V114 V117 1.4857020261645263e-12
C114_117 V114 V117 3.554062187547961e-19

R114_118 V114 V118 10146.39450917041
L114_118 V114 V118 8.087343526814079e-13
C114_118 V114 V118 6.903184030993867e-19

R114_119 V114 V119 1776.1275535263176
L114_119 V114 V119 6.98087130692516e-13
C114_119 V114 V119 1.035063206636014e-18

R114_120 V114 V120 504.07907719833815
L114_120 V114 V120 3.1624438031031674e-12
C114_120 V114 V120 3.3508689289635865e-19

R114_121 V114 V121 -2846.1991487824225
L114_121 V114 V121 -1.0360020649122618e-12
C114_121 V114 V121 -1.7586523994526406e-19

R114_122 V114 V122 622.2535039607094
L114_122 V114 V122 -6.948030232760169e-13
C114_122 V114 V122 -1.2146549263125215e-20

R114_123 V114 V123 -1318.6044235243653
L114_123 V114 V123 -1.919933022240252e-12
C114_123 V114 V123 1.898261505017884e-19

R114_124 V114 V124 -577.2126998579348
L114_124 V114 V124 1.3793680266613147e-11
C114_124 V114 V124 2.7318056441147596e-19

R114_125 V114 V125 1675.6009687639444
L114_125 V114 V125 1.456548060548797e-12
C114_125 V114 V125 1.2481215945981208e-19

R114_126 V114 V126 -371.041275672592
L114_126 V114 V126 1.0309588522263671e-12
C114_126 V114 V126 -1.2023423781120349e-19

R114_127 V114 V127 420.4777092745274
L114_127 V114 V127 -1.6284629371129017e-12
C114_127 V114 V127 1.8323443394326005e-20

R114_128 V114 V128 683.1105843498665
L114_128 V114 V128 -3.574783019255304e-12
C114_128 V114 V128 3.8199738902032994e-20

R114_129 V114 V129 -1122.2323118744678
L114_129 V114 V129 -1.5782980937501837e-12
C114_129 V114 V129 1.596319982109227e-19

R114_130 V114 V130 634.7258625545002
L114_130 V114 V130 8.495457807520523e-13
C114_130 V114 V130 2.2130527041915244e-19

R114_131 V114 V131 1006.1471915337298
L114_131 V114 V131 2.367351912306446e-12
C114_131 V114 V131 -2.3927026176723617e-19

R114_132 V114 V132 -2161.7186304213
L114_132 V114 V132 3.894266083405928e-12
C114_132 V114 V132 1.1400229679047642e-20

R114_133 V114 V133 5076.460306829367
L114_133 V114 V133 -2.8804163207337278e-12
C114_133 V114 V133 -4.598621160856926e-19

R114_134 V114 V134 -2872.4716680616857
L114_134 V114 V134 8.116627229232212e-12
C114_134 V114 V134 -1.767634353730004e-20

R114_135 V114 V135 657.9022769053436
L114_135 V114 V135 -3.0065160460665572e-12
C114_135 V114 V135 1.0514657792876396e-19

R114_136 V114 V136 1167.4488551124568
L114_136 V114 V136 1.2322900027897087e-11
C114_136 V114 V136 6.860313397095259e-20

R114_137 V114 V137 -10530.264420822787
L114_137 V114 V137 1.9211507334842362e-12
C114_137 V114 V137 2.903782904154834e-19

R114_138 V114 V138 -1150.0382048593642
L114_138 V114 V138 6.303220735033944e-13
C114_138 V114 V138 1.51752984578693e-19

R114_139 V114 V139 320.6587934102229
L114_139 V114 V139 -1.0424242465607651e-12
C114_139 V114 V139 -1.6789867876630791e-19

R114_140 V114 V140 9201.76679296835
L114_140 V114 V140 1.6654855948059074e-12
C114_140 V114 V140 1.0403572911394456e-19

R114_141 V114 V141 -599.5496072827532
L114_141 V114 V141 3.049728408540781e-12
C114_141 V114 V141 7.733188280540646e-20

R114_142 V114 V142 874.240676381632
L114_142 V114 V142 8.167296927184583e-13
C114_142 V114 V142 2.1631914529691622e-19

R114_143 V114 V143 -2754.9334143175624
L114_143 V114 V143 3.252176508957881e-12
C114_143 V114 V143 -2.8110031382032773e-20

R114_144 V114 V144 20686.00278690269
L114_144 V114 V144 -2.1447309742080445e-12
C114_144 V114 V144 -1.0486396433219628e-19

R115_115 V115 0 -179.53531371831613
L115_115 V115 0 -2.6993338843624714e-12
C115_115 V115 0 -1.1311263448097833e-19

R115_116 V115 V116 -122113.55926399652
L115_116 V115 V116 7.973263369321364e-13
C115_116 V115 V116 6.440347290374472e-19

R115_117 V115 V117 1695.746676656245
L115_117 V115 V117 1.8101709405361776e-12
C115_117 V115 V117 5.162978845141175e-19

R115_118 V115 V118 50625.51715586727
L115_118 V115 V118 1.2185933968553858e-12
C115_118 V115 V118 3.874153932414121e-19

R115_119 V115 V119 -4114.904765414535
L115_119 V115 V119 8.372194631004879e-13
C115_119 V115 V119 5.418137308662714e-19

R115_120 V115 V120 446.194368298763
L115_120 V115 V120 -9.41045546357354e-13
C115_120 V115 V120 2.632266875215146e-19

R115_121 V115 V121 -3001.8729838862796
L115_121 V115 V121 -8.780152091979262e-12
C115_121 V115 V121 -1.1722337337386456e-19

R115_122 V115 V122 457.8959938575269
L115_122 V115 V122 -7.223320479508108e-13
C115_122 V115 V122 1.4878089347328245e-21

R115_123 V115 V123 3333.7843543876834
L115_123 V115 V123 -2.7595230809513897e-12
C115_123 V115 V123 5.383753341415795e-20

R115_124 V115 V124 -2388.085960339204
L115_124 V115 V124 2.9545581102628185e-12
C115_124 V115 V124 1.7262270077434797e-19

R115_125 V115 V125 1051.3616721056158
L115_125 V115 V125 -2.488753631555803e-12
C115_125 V115 V125 8.061418142021017e-20

R115_126 V115 V126 -302.84647726159915
L115_126 V115 V126 5.291026851229902e-13
C115_126 V115 V126 -1.7661783111903177e-19

R115_127 V115 V127 385.2630394812019
L115_127 V115 V127 -5.87865471391969e-13
C115_127 V115 V127 -1.9966042658678473e-20

R115_128 V115 V128 2272.8896283915897
L115_128 V115 V128 -6.131356843221277e-12
C115_128 V115 V128 1.0443288508748792e-21

R115_129 V115 V129 1540.730073860485
L115_129 V115 V129 -1.5943358907361057e-12
C115_129 V115 V129 2.6664595425177722e-20

R115_130 V115 V130 -5124.0522448300735
L115_130 V115 V130 8.749366446305137e-13
C115_130 V115 V130 3.43500960482574e-19

R115_131 V115 V131 -1497.3211684252835
L115_131 V115 V131 1.143653738735295e-11
C115_131 V115 V131 -3.674566073960945e-19

R115_132 V115 V132 -1720.2280583136776
L115_132 V115 V132 2.324216716997135e-12
C115_132 V115 V132 3.37689855698244e-20

R115_133 V115 V133 -14827.932991381524
L115_133 V115 V133 -1.991812166343719e-12
C115_133 V115 V133 -3.1385561841853296e-19

R115_134 V115 V134 -2697.4879289689525
L115_134 V115 V134 2.415114627430571e-11
C115_134 V115 V134 -5.766512079916924e-20

R115_135 V115 V135 548.3922557275972
L115_135 V115 V135 -9.882326517116484e-13
C115_135 V115 V135 1.474162388431612e-19

R115_136 V115 V136 4974.8846404944
L115_136 V115 V136 -1.3080318987242657e-10
C115_136 V115 V136 3.020993859038143e-20

R115_137 V115 V137 3118.686524474772
L115_137 V115 V137 -5.950840638644562e-11
C115_137 V115 V137 1.5170845391999417e-19

R115_138 V115 V138 -421.3817444130977
L115_138 V115 V138 5.377678099174053e-13
C115_138 V115 V138 1.119429722172684e-19

R115_139 V115 V139 305.36256659744924
L115_139 V115 V139 -4.3229020110675527e-13
C115_139 V115 V139 -1.7241498840363524e-19

R115_140 V115 V140 -1679.3004565051674
L115_140 V115 V140 1.2916308584541919e-12
C115_140 V115 V140 1.0596373351456298e-19

R115_141 V115 V141 -1319.6812580947624
L115_141 V115 V141 2.219473236282502e-12
C115_141 V115 V141 4.920980130482824e-20

R115_142 V115 V142 -2005.403472131729
L115_142 V115 V142 1.210567733478981e-12
C115_142 V115 V142 9.686329032319888e-20

R115_143 V115 V143 -993.7799531386817
L115_143 V115 V143 1.0940320166774853e-12
C115_143 V115 V143 6.608595862874914e-20

R115_144 V115 V144 3269.324974620704
L115_144 V115 V144 -1.5469079785109903e-12
C115_144 V115 V144 -1.667692105687878e-19

R116_116 V116 0 371.5549032306537
L116_116 V116 0 2.2238103987506218e-13
C116_116 V116 0 1.1865879779411622e-18

R116_117 V116 V117 -1599.6111832393233
L116_117 V116 V117 -1.188338487867191e-12
C116_117 V116 V117 -5.456724182105055e-19

R116_118 V116 V118 50624.27820356332
L116_118 V116 V118 -8.612911379961018e-13
C116_118 V116 V118 -4.454322670242336e-19

R116_119 V116 V119 6344.4988786122085
L116_119 V116 V119 -7.038551199669142e-13
C116_119 V116 V119 -7.725732120875248e-19

R116_120 V116 V120 -522.5898387313877
L116_120 V116 V120 7.170960621385788e-12
C116_120 V116 V120 -3.591457712142308e-19

R116_121 V116 V121 -11199.54586428978
L116_121 V116 V121 1.3270759068344906e-12
C116_121 V116 V121 4.381319268759097e-20

R116_122 V116 V122 -444.9216138786121
L116_122 V116 V122 5.522329242830802e-13
C116_122 V116 V122 -9.459830369265282e-21

R116_123 V116 V123 -1992.4404178942314
L116_123 V116 V123 1.0459521958383885e-11
C116_123 V116 V123 -6.441202697335594e-20

R116_124 V116 V124 -14045.951068250797
L116_124 V116 V124 -2.563110854645921e-12
C116_124 V116 V124 -2.8553805073581954e-19

R116_125 V116 V125 -1803.1828421116002
L116_125 V116 V125 -1.0124971406182008e-12
C116_125 V116 V125 -2.5597836790288984e-19

R116_126 V116 V126 324.36558419990513
L116_126 V116 V126 -5.730292134817366e-13
C116_126 V116 V126 1.0435168407206929e-19

R116_127 V116 V127 -430.51628863027065
L116_127 V116 V127 7.047533988130924e-13
C116_127 V116 V127 -2.8495164930116174e-20

R116_128 V116 V128 -28595.914863296104
L116_128 V116 V128 7.614102919900151e-11
C116_128 V116 V128 8.616822195981053e-21

R116_129 V116 V129 -1020.6880119561558
L116_129 V116 V129 2.1814258657090225e-12
C116_129 V116 V129 -5.096141826545221e-20

R116_130 V116 V130 1969.6818507599835
L116_130 V116 V130 -1.100748139997766e-12
C116_130 V116 V130 -3.7768910309751543e-19

R116_131 V116 V131 1070.6852280851233
L116_131 V116 V131 1.3139307063084319e-11
C116_131 V116 V131 2.6563747089094024e-19

R116_132 V116 V132 2035.5131250091674
L116_132 V116 V132 -1.8090577315412824e-12
C116_132 V116 V132 -9.976671413859232e-20

R116_133 V116 V133 3751.3699062208325
L116_133 V116 V133 3.2622946636769024e-12
C116_133 V116 V133 2.8661238198272393e-19

R116_134 V116 V134 2282.14561856463
L116_134 V116 V134 -1.7958830615997445e-12
C116_134 V116 V134 -1.0042724456054441e-20

R116_135 V116 V135 -606.3271306166532
L116_135 V116 V135 1.3264861778305441e-12
C116_135 V116 V135 -1.2869502353056137e-19

R116_136 V116 V136 17167.71420742351
L116_136 V116 V136 -1.0991306841505822e-11
C116_136 V116 V136 -3.374978145590449e-21

R116_137 V116 V137 -3772.975737327728
L116_137 V116 V137 -1.8970400834338e-12
C116_137 V116 V137 -1.4118557825701463e-19

R116_138 V116 V138 397.615874896514
L116_138 V116 V138 -5.633698323629242e-13
C116_138 V116 V138 -1.4595418875862758e-19

R116_139 V116 V139 -344.71255704054073
L116_139 V116 V139 5.121128984483917e-13
C116_139 V116 V139 1.1459906480705504e-19

R116_140 V116 V140 1337.552518250572
L116_140 V116 V140 -1.0913359233559926e-12
C116_140 V116 V140 -1.0458127315359815e-19

R116_141 V116 V141 2196.652057484249
L116_141 V116 V141 -2.609509220371814e-12
C116_141 V116 V141 -3.102383891334714e-20

R116_142 V116 V142 1308.5708596856432
L116_142 V116 V142 -1.549276523908475e-12
C116_142 V116 V142 -1.1964094656506627e-19

R116_143 V116 V143 1006.714923083607
L116_143 V116 V143 -1.3216726164924236e-12
C116_143 V116 V143 -1.7304014412212344e-19

R116_144 V116 V144 -2709.304870478691
L116_144 V116 V144 1.613035861943525e-12
C116_144 V116 V144 4.94226675283913e-20

R117_117 V117 0 -138.66190948684235
L117_117 V117 0 1.2431466852589839e-12
C117_117 V117 0 -2.531449822441048e-20

R117_118 V117 V118 -2515.8929029880487
L117_118 V117 V118 -1.0768167748607996e-12
C117_118 V117 V118 -4.947009238455512e-19

R117_119 V117 V119 -1290.6838920836879
L117_119 V117 V119 -1.95134778737025e-12
C117_119 V117 V119 -4.039372923068937e-19

R117_120 V117 V120 361.7956554283538
L117_120 V117 V120 -5.363141185614054e-12
C117_120 V117 V120 -1.1288669837140915e-19

R117_121 V117 V121 -14757.486882727819
L117_121 V117 V121 1.0203496992866048e-12
C117_121 V117 V121 8.097568032837311e-20

R117_122 V117 V122 299.8463784891527
L117_122 V117 V122 6.393376861350754e-13
C117_122 V117 V122 5.749719173851631e-20

R117_123 V117 V123 1997.1277420649608
L117_123 V117 V123 4.321732115478533e-12
C117_123 V117 V123 -8.243648951842933e-20

R117_124 V117 V124 -3529.480176214254
L117_124 V117 V124 -7.428500935206354e-12
C117_124 V117 V124 -1.819167424376483e-20

R117_125 V117 V125 1129.6649169750085
L117_125 V117 V125 -1.0200612379575085e-12
C117_125 V117 V125 -1.3401931778929526e-19

R117_126 V117 V126 -219.28941778606313
L117_126 V117 V126 -1.0314946531539009e-12
C117_126 V117 V126 1.3522569428529703e-19

R117_127 V117 V127 276.05686996947225
L117_127 V117 V127 1.4706122204574898e-12
C117_127 V117 V127 5.478135904403077e-20

R117_128 V117 V128 5166.864996680195
L117_128 V117 V128 6.3873817700397945e-12
C117_128 V117 V128 -1.0657115861102334e-19

R117_129 V117 V129 894.6185915783826
L117_129 V117 V129 6.9691725327830394e-12
C117_129 V117 V129 -8.463557159534177e-20

R117_130 V117 V130 -1066.0009149156558
L117_130 V117 V130 -1.5220658128454782e-12
C117_130 V117 V130 -3.9354228900613004e-19

R117_131 V117 V131 -1108.603635000182
L117_131 V117 V131 -5.518916773849751e-12
C117_131 V117 V131 1.9335616061481755e-19

R117_132 V117 V132 -1234.6360254846873
L117_132 V117 V132 -3.3975355102072956e-12
C117_132 V117 V132 -2.825057340720027e-20

R117_133 V117 V133 -115020.3470962603
L117_133 V117 V133 4.543500744761514e-12
C117_133 V117 V133 3.04880719448199e-19

R117_134 V117 V134 -1907.577758997341
L117_134 V117 V134 -3.547440225858547e-12
C117_134 V117 V134 3.7187493399924237e-20

R117_135 V117 V135 414.59946846031244
L117_135 V117 V135 2.459606565413815e-12
C117_135 V117 V135 -8.248607390159268e-20

R117_136 V117 V136 25100.432724165712
L117_136 V117 V136 5.991411034290093e-12
C117_136 V117 V136 7.473569372455058e-20

R117_137 V117 V137 4498.322581106973
L117_137 V117 V137 -1.5141341404881709e-12
C117_137 V117 V137 -8.746693591134066e-20

R117_138 V117 V138 -266.68120412986724
L117_138 V117 V138 -9.655018203744045e-13
C117_138 V117 V138 8.41449527178164e-21

R117_139 V117 V139 214.1928073347926
L117_139 V117 V139 1.0960031426308292e-12
C117_139 V117 V139 1.1077696261689342e-19

R117_140 V117 V140 -878.6596593280558
L117_140 V117 V140 -2.1488293112720454e-12
C117_140 V117 V140 -9.354413320509423e-20

R117_141 V117 V141 -1109.4108251292412
L117_141 V117 V141 -2.4969396212449448e-12
C117_141 V117 V141 -2.5545567758031072e-20

R117_142 V117 V142 -968.9659126413526
L117_142 V117 V142 -1.858133975853699e-12
C117_142 V117 V142 -1.1608759331213883e-19

R117_143 V117 V143 -668.0000896688753
L117_143 V117 V143 -4.034644158319769e-12
C117_143 V117 V143 -5.2548652473141486e-20

R117_144 V117 V144 1590.4750779257724
L117_144 V117 V144 2.986187791324857e-12
C117_144 V117 V144 4.866886381831228e-20

R118_118 V118 0 271.1950646470928
L118_118 V118 0 3.5272294026611415e-13
C118_118 V118 0 1.8565395592332158e-19

R118_119 V118 V119 -3691.8893897930275
L118_119 V118 V119 -8.245689914084008e-13
C118_119 V118 V119 -7.3871001392692135e-19

R118_120 V118 V120 -1109.9791921062933
L118_120 V118 V120 1.0707651739703628e-11
C118_120 V118 V120 -1.0211535890127289e-19

R118_121 V118 V121 -1240.3565493126919
L118_121 V118 V121 1.1621057240004487e-12
C118_121 V118 V121 1.6138110671694415e-19

R118_122 V118 V122 -397.1430462599627
L118_122 V118 V122 7.237189559083094e-13
C118_122 V118 V122 -3.096919224374383e-20

R118_123 V118 V123 -1685.7486596066278
L118_123 V118 V123 6.106524054944576e-12
C118_123 V118 V123 -1.5123241329028187e-19

R118_124 V118 V124 -1852531.5088180793
L118_124 V118 V124 -3.5711336195061548e-12
C118_124 V118 V124 -1.0651645041186093e-19

R118_125 V118 V125 2013.3920090667739
L118_125 V118 V125 -1.1856655253865538e-12
C118_125 V118 V125 -2.1423219256427932e-19

R118_126 V118 V126 379.4642702714141
L118_126 V118 V126 -8.500825974073631e-13
C118_126 V118 V126 9.004496554460081e-20

R118_127 V118 V127 -592.9929163416987
L118_127 V118 V127 1.1294152419916284e-12
C118_127 V118 V127 2.065579196257463e-20

R118_128 V118 V128 -3595.372435286732
L118_128 V118 V128 3.702671422204897e-12
C118_128 V118 V128 -1.013578882185212e-19

R118_129 V118 V129 -1350.8183133587172
L118_129 V118 V129 2.5895536244411822e-12
C118_129 V118 V129 -1.9179586497229708e-20

R118_130 V118 V130 2208.316888515251
L118_130 V118 V130 -1.245140344252044e-12
C118_130 V118 V130 -3.0677379578322998e-19

R118_131 V118 V131 1171.0325955779779
L118_131 V118 V131 -1.168554077407052e-11
C118_131 V118 V131 1.487265217252734e-19

R118_132 V118 V132 1737.4353634441186
L118_132 V118 V132 -5.570595887482486e-12
C118_132 V118 V132 7.477126093950964e-20

R118_133 V118 V133 2107.9112267428222
L118_133 V118 V133 1.7621920976241448e-12
C118_133 V118 V133 4.836542274795666e-19

R118_134 V118 V134 2225.597313935729
L118_134 V118 V134 -2.9536027677587477e-12
C118_134 V118 V134 -6.849637003036871e-20

R118_135 V118 V135 -805.1618383593442
L118_135 V118 V135 2.1518445318329626e-12
C118_135 V118 V135 -6.955674888999413e-20

R118_136 V118 V136 -74474.69037078823
L118_136 V118 V136 1.0450304860634893e-11
C118_136 V118 V136 -2.098073252681497e-20

R118_137 V118 V137 2688.652502850957
L118_137 V118 V137 -1.7269646842736808e-12
C118_137 V118 V137 -1.8984969527110277e-19

R118_138 V118 V138 439.6788269472195
L118_138 V118 V138 -7.978245956472194e-13
C118_138 V118 V138 -1.2425166083909752e-20

R118_139 V118 V139 -465.79149058303597
L118_139 V118 V139 7.834327943875414e-13
C118_139 V118 V139 1.4699374207650888e-19

R118_140 V118 V140 1648.594080659355
L118_140 V118 V140 -2.1043795873938868e-12
C118_140 V118 V140 -4.61510336038419e-20

R118_141 V118 V141 1898.1851411937403
L118_141 V118 V141 -2.392924609366501e-12
C118_141 V118 V141 -1.1679933927925742e-20

R118_142 V118 V142 1618.8783588793578
L118_142 V118 V142 -1.4794755925563361e-12
C118_142 V118 V142 -6.965666155824553e-20

R118_143 V118 V143 1557.5385586971831
L118_143 V118 V143 -2.288659884743131e-12
C118_143 V118 V143 -7.248129604279829e-20

R118_144 V118 V144 -2411.2480541282853
L118_144 V118 V144 2.8750039024152648e-12
C118_144 V118 V144 6.383459848934823e-20

R119_119 V119 0 92.0987838575315
L119_119 V119 0 2.6086842035128073e-13
C119_119 V119 0 4.261737301931084e-19

R119_120 V119 V120 -238.62334059659565
L119_120 V119 V120 2.0849571497236627e-12
C119_120 V119 V120 -4.552514727421929e-19

R119_121 V119 V121 502.74822595338634
L119_121 V119 V121 1.075821755489888e-11
C119_121 V119 V121 1.7691385904759205e-19

R119_122 V119 V122 -593.1654905207131
L119_122 V119 V122 1.98782117360595e-12
C119_122 V119 V122 3.8959577217310023e-20

R119_123 V119 V123 4791.554535508928
L119_123 V119 V123 -4.226343555250645e-12
C119_123 V119 V123 -2.0385258026953714e-19

R119_124 V119 V124 927.4437710985959
L119_124 V119 V124 -1.7524250564617998e-12
C119_124 V119 V124 -4.1816492854279016e-19

R119_125 V119 V125 -330.80379699816666
L119_125 V119 V125 5.223927494113943e-12
C119_125 V119 V125 -1.9796079498291572e-19

R119_126 V119 V126 233.7298138923442
L119_126 V119 V126 -9.850334736908965e-13
C119_126 V119 V126 1.2344570834781315e-19

R119_127 V119 V127 -250.73119254258148
L119_127 V119 V127 8.956039626939494e-13
C119_127 V119 V127 -3.862602891971693e-20

R119_128 V119 V128 -1375.6590171054827
L119_128 V119 V128 1.0732255834736201e-10
C119_128 V119 V128 -3.0292262175593445e-21

R119_129 V119 V129 -2271.925208133375
L119_129 V119 V129 2.964515617162461e-12
C119_129 V119 V129 -1.0871596773768577e-19

R119_130 V119 V130 -5255.639186581371
L119_130 V119 V130 -1.577288539506119e-12
C119_130 V119 V130 -2.679382623436755e-19

R119_131 V119 V131 16532.017748796166
L119_131 V119 V131 3.3971113939353e-12
C119_131 V119 V131 2.4739927307761788e-19

R119_132 V119 V132 1515.8312148877837
L119_132 V119 V132 -3.8528147718623565e-12
C119_132 V119 V132 -3.0985685077305646e-20

R119_133 V119 V133 -2903.82170295399
L119_133 V119 V133 1.034602452994045e-12
C119_133 V119 V133 6.049874037809745e-19

R119_134 V119 V134 6224.48563451366
L119_134 V119 V134 -8.025408401537226e-12
C119_134 V119 V134 -7.157485739656414e-20

R119_135 V119 V135 -390.08989881379046
L119_135 V119 V135 1.7294956064813066e-12
C119_135 V119 V135 -8.314296610647154e-20

R119_136 V119 V136 -2047.23418389099
L119_136 V119 V136 -1.17791640591802e-11
C119_136 V119 V136 -7.624878435611735e-20

R119_137 V119 V137 -738.8497360766688
L119_137 V119 V137 9.477715776977267e-12
C119_137 V119 V137 -2.8446726620261824e-19

R119_138 V119 V138 398.59025421338106
L119_138 V119 V138 -1.0972036026285248e-12
C119_138 V119 V138 -1.3010037616384196e-19

R119_139 V119 V139 -196.47504060334649
L119_139 V119 V139 6.836009846255033e-13
C119_139 V119 V139 1.1131915911325085e-19

R119_140 V119 V140 1825.047404276262
L119_140 V119 V140 -1.5060577609375058e-12
C119_140 V119 V140 -1.3982568958793007e-19

R119_141 V119 V141 857.3131011415492
L119_141 V119 V141 -3.81069423301881e-12
C119_141 V119 V141 -8.58554816328099e-20

R119_142 V119 V142 8585.807709548546
L119_142 V119 V142 -1.5409362716020167e-12
C119_142 V119 V142 -1.9378222689838156e-19

R119_143 V119 V143 656.3822649472994
L119_143 V119 V143 -1.5159506568208227e-12
C119_143 V119 V143 -9.262092950118192e-20

R119_144 V119 V144 -7568.892744684605
L119_144 V119 V144 2.4348534845755727e-12
C119_144 V119 V144 1.314577879293619e-19

R120_120 V120 0 -35.570452881683345
L120_120 V120 0 5.4291107567944e-13
C120_120 V120 0 1.7499460422578848e-19

R120_121 V120 V121 -480.23989088193866
L120_121 V120 V121 7.709203588304925e-13
C120_121 V120 V121 1.8524647002735297e-20

R120_122 V120 V122 68.03859834014818
L120_122 V120 V122 2.3643689044542025e-12
C120_122 V120 V122 1.5808943003545472e-20

R120_123 V120 V123 293.49346015437584
L120_123 V120 V123 4.325905532721399e-12
C120_123 V120 V123 -3.522418509589183e-20

R120_124 V120 V124 -1033.893487470803
L120_124 V120 V124 4.143250226391128e-12
C120_124 V120 V124 -2.1759454906595614e-19

R120_125 V120 V125 146.19723414380522
L120_125 V120 V125 -5.168538958437563e-13
C120_125 V120 V125 -3.3677826864110206e-20

R120_126 V120 V126 -45.81363034105781
L120_126 V120 V126 8.402371359308281e-13
C120_126 V120 V126 5.018651529445156e-20

R120_127 V120 V127 57.4902942237443
L120_127 V120 V127 -6.260144041092648e-13
C120_127 V120 V127 -3.270575093241781e-20

R120_128 V120 V128 924.234052712467
L120_128 V120 V128 1.750490633493032e-11
C120_128 V120 V128 3.692905992816094e-20

R120_129 V120 V129 148.01328783792505
L120_129 V120 V129 -1.9722015829130615e-12
C120_129 V120 V129 -7.386421289346667e-20

R120_130 V120 V130 -196.920386764708
L120_130 V120 V130 3.843474451911025e-12
C120_130 V120 V130 -1.0220414390818963e-19

R120_131 V120 V131 -177.5247821928216
L120_131 V120 V131 -1.9495562575815254e-12
C120_131 V120 V131 1.0997409573416195e-19

R120_132 V120 V132 -243.30548479304647
L120_132 V120 V132 1.6096485349691895e-11
C120_132 V120 V132 -6.383694570157074e-20

R120_133 V120 V133 -7387.46173125066
L120_133 V120 V133 -2.3680541157910844e-12
C120_133 V120 V133 1.631620347781497e-19

R120_134 V120 V134 -421.9104160216376
L120_134 V120 V134 -3.5581575245314925e-11
C120_134 V120 V134 2.049157983029558e-20

R120_135 V120 V135 84.69756564631994
L120_135 V120 V135 -1.214779046460753e-12
C120_135 V120 V135 -6.206159206003911e-20

R120_136 V120 V136 3317.9651404954348
L120_136 V120 V136 -5.569948717368931e-12
C120_136 V120 V136 -5.177306840481918e-20

R120_137 V120 V137 354.5052388905702
L120_137 V120 V137 -8.668198433123652e-13
C120_137 V120 V137 -1.4266715539230185e-19

R120_138 V120 V138 -55.21391895685029
L120_138 V120 V138 1.6584985755414649e-12
C120_138 V120 V138 -9.686644992872894e-20

R120_139 V120 V139 44.773066974640024
L120_139 V120 V139 -4.761704996029088e-13
C120_139 V120 V139 6.288464917565367e-20

R120_140 V120 V140 -188.9590980842649
L120_140 V120 V140 7.941172271634764e-12
C120_140 V120 V140 -6.897075045443204e-20

R120_141 V120 V141 -291.06199838885374
L120_141 V120 V141 6.083172859135727e-12
C120_141 V120 V141 -1.876011202589298e-20

R120_142 V120 V142 -164.94776071677043
L120_142 V120 V142 9.203080446968545e-12
C120_142 V120 V142 -7.483137560416627e-20

R120_143 V120 V143 -128.02813673914136
L120_143 V120 V143 1.1934093641597091e-12
C120_143 V120 V143 -1.0007657228896693e-20

R120_144 V120 V144 411.05453693468456
L120_144 V120 V144 1.3172208192115902e-11
C120_144 V120 V144 7.425085497362487e-20

R121_121 V121 0 206.35812666607848
L121_121 V121 0 -3.090348050816306e-13
C121_121 V121 0 -1.4635097930916712e-19

R121_122 V121 V122 145.34879367480175
L121_122 V121 V122 -4.017072941476061e-13
C121_122 V121 V122 9.678362320068543e-21

R121_123 V121 V123 1071.3687772223298
L121_123 V121 V123 -1.7226184557493563e-12
C121_123 V121 V123 6.876373268975384e-20

R121_124 V121 V124 1897.4170203113467
L121_124 V121 V124 -1.6128356294103523e-12
C121_124 V121 V124 2.0727767129980652e-20

R121_125 V121 V125 -156.67416965857527
L121_125 V121 V125 4.194748499309972e-13
C121_125 V121 V125 2.0595049481570706e-20

R121_126 V121 V126 -251.81371651516753
L121_126 V121 V126 1.1575675103402214e-12
C121_126 V121 V126 -3.152388988786227e-20

R121_127 V121 V127 731.9973907253852
L121_127 V121 V127 -7.15827165822683e-12
C121_127 V121 V127 -1.1662363304800731e-20

R121_128 V121 V128 5927.825904808108
L121_128 V121 V128 4.503616519652692e-12
C121_128 V121 V128 3.467144864870956e-20

R121_129 V121 V129 2002.7140330578343
L121_129 V121 V129 -2.971142481513626e-12
C121_129 V121 V129 1.8786087278479808e-20

R121_130 V121 V130 -4788.680825314476
L121_130 V121 V130 1.0219718968149788e-12
C121_130 V121 V130 4.3562935262618293e-20

R121_131 V121 V131 -755.1855689017451
L121_131 V121 V131 1.3138101566054184e-12
C121_131 V121 V131 -6.471900359643509e-20

R121_132 V121 V132 -1101.6789925905266
L121_132 V121 V132 3.4887981640193922e-12
C121_132 V121 V132 -2.536403363413189e-21

R121_133 V121 V133 -579.3821590408502
L121_133 V121 V133 2.3829283210408014e-12
C121_133 V121 V133 -9.351464901603398e-20

R121_134 V121 V134 -640.8832645089565
L121_134 V121 V134 1.948181016939348e-12
C121_134 V121 V134 7.218845134637121e-21

R121_135 V121 V135 782.6812548563767
L121_135 V121 V135 -6.290975704180912e-12
C121_135 V121 V135 2.2102252332143025e-20

R121_136 V121 V136 -2929.997319033796
L121_136 V121 V136 3.704866174992294e-12
C121_136 V121 V136 -4.091185645996068e-20

R121_137 V121 V137 -279.15431816928896
L121_137 V121 V137 6.952936535370325e-13
C121_137 V121 V137 -1.0965919898605918e-20

R121_138 V121 V138 -253.85688488456125
L121_138 V121 V138 6.315243886298318e-13
C121_138 V121 V138 3.1029544672843155e-21

R121_139 V121 V139 612.0006108083026
L121_139 V121 V139 -4.8121569201785954e-12
C121_139 V121 V139 -4.270843600959797e-20

R121_140 V121 V140 -657.9764426993158
L121_140 V121 V140 1.2790990250156176e-12
C121_140 V121 V140 -7.798074571945867e-21

R121_141 V121 V141 -766.4949007426469
L121_141 V121 V141 7.780623852241129e-12
C121_141 V121 V141 2.3440225912752888e-20

R121_142 V121 V142 -2119.099519546881
L121_142 V121 V142 1.0465453173277735e-12
C121_142 V121 V142 7.704001201414806e-20

R121_143 V121 V143 9868.486762342685
L121_143 V121 V143 -1.2786468483724138e-11
C121_143 V121 V143 2.7752004394331426e-21

R121_144 V121 V144 686.7832589522354
L121_144 V121 V144 -1.5835382883560208e-12
C121_144 V121 V144 1.1255514940815456e-20

R122_122 V122 0 -41.40662616206168
L122_122 V122 0 -4.1119288365104555e-13
C122_122 V122 0 4.100383716013942e-19

R122_123 V122 V123 179.56102154609988
L122_123 V122 V123 -7.075966844265469e-13
C122_123 V122 V123 -3.839099565345133e-20

R122_124 V122 V124 -1159.6455586329505
L122_124 V122 V124 -1.9302019671971204e-12
C122_124 V122 V124 -6.658463068610309e-21

R122_125 V122 V125 -559.7943508887614
L122_125 V122 V125 4.146502337528446e-13
C122_125 V122 V125 -4.120293851646996e-20

R122_126 V122 V126 -30.25158566120376
L122_126 V122 V126 3.4649801634583646e-13
C122_126 V122 V126 -3.646001209482313e-20

R122_127 V122 V127 42.55089445119195
L122_127 V122 V127 -5.90044654371425e-13
C122_127 V122 V127 -9.443481680691853e-23

R122_128 V122 V128 442.1835148674448
L122_128 V122 V128 -8.831823317264115e-12
C122_128 V122 V128 1.0708892489290935e-20

R122_129 V122 V129 113.85322825965822
L122_129 V122 V129 -9.16650552958387e-13
C122_129 V122 V129 4.493863797931535e-20

R122_130 V122 V130 -165.20349530212846
L122_130 V122 V130 4.1712244105204597e-13
C122_130 V122 V130 2.0391694143756943e-20

R122_131 V122 V131 -115.09461843743784
L122_131 V122 V131 8.798419202565547e-13
C122_131 V122 V131 1.181649440649331e-20

R122_132 V122 V132 -156.51511464039075
L122_132 V122 V132 1.3491433830889869e-12
C122_132 V122 V132 1.8027427442964427e-20

R122_133 V122 V133 -350.7151710800617
L122_133 V122 V133 2.681952568862068e-12
C122_133 V122 V133 -4.9829240723712273e-20

R122_134 V122 V134 -183.84315627694085
L122_134 V122 V134 1.657566748884823e-12
C122_134 V122 V134 -1.4856014135428596e-20

R122_135 V122 V135 60.550688990615896
L122_135 V122 V135 -8.233615890732112e-13
C122_135 V122 V135 -3.961396561241715e-20

R122_136 V122 V136 6324.3927708465735
L122_136 V122 V136 4.653310892735055e-12
C122_136 V122 V136 -1.6256333904503344e-20

R122_137 V122 V137 -428.96811666628116
L122_137 V122 V137 5.960211380267689e-13
C122_137 V122 V137 5.568821483027867e-20

R122_138 V122 V138 -35.41216969543673
L122_138 V122 V138 2.616671094036477e-13
C122_138 V122 V138 -8.917497905886164e-21

R122_139 V122 V139 33.28998381576252
L122_139 V122 V139 -4.1820704803875397e-13
C122_139 V122 V139 9.782614001010768e-21

R122_140 V122 V140 -116.79001319880933
L122_140 V122 V140 6.261964260816156e-13
C122_140 V122 V140 6.883250293351364e-21

R122_141 V122 V141 -148.3814533879306
L122_141 V122 V141 1.453864008672294e-12
C122_141 V122 V141 -2.0973563042992544e-20

R122_142 V122 V142 -127.95576673145334
L122_142 V122 V142 5.568209156161724e-13
C122_142 V122 V142 -3.3282352793645476e-20

R122_143 V122 V143 -107.98679793694089
L122_143 V122 V143 1.3267746974526792e-12
C122_143 V122 V143 -1.305696940330993e-20

R122_144 V122 V144 194.6493282067632
L122_144 V122 V144 -8.194159294068901e-13
C122_144 V122 V144 -3.380983569537306e-20

R123_123 V123 0 -96.96214548005908
L123_123 V123 0 -4.417392821569349e-12
C123_123 V123 0 4.501535960472026e-19

R123_124 V123 V124 -471.72657443678344
L123_124 V123 V124 -2.0975037475894875e-12
C123_124 V123 V124 -7.107932735911689e-20

R123_125 V123 V125 -8368.588293988498
L123_125 V123 V125 2.183469004889478e-12
C123_125 V123 V125 -4.202757661983682e-20

R123_126 V123 V126 -147.05857251773378
L123_126 V123 V126 1.4720235109892651e-12
C123_126 V123 V126 -6.317659865067078e-21

R123_127 V123 V127 192.62423982313896
L123_127 V123 V127 -6.578045408928109e-12
C123_127 V123 V127 2.8593467536564526e-21

R123_128 V123 V128 484.74404511455646
L123_128 V123 V128 -2.624282645063776e-12
C123_128 V123 V128 -1.0577513226953784e-20

R123_129 V123 V129 17850.356833118178
L123_129 V123 V129 -8.9461106390026e-13
C123_129 V123 V129 -3.543757228555038e-20

R123_130 V123 V130 1259.1444788827166
L123_130 V123 V130 7.840254330987638e-13
C123_130 V123 V130 -8.997167449516444e-21

R123_131 V123 V131 53426.02681851288
L123_131 V123 V131 9.557012693169594e-13
C123_131 V123 V131 2.904872309627292e-20

R123_132 V123 V132 -785.0030541019709
L123_132 V123 V132 7.898617446936314e-12
C123_132 V123 V132 6.396205803243851e-21

R123_133 V123 V133 -30082.466389791498
L123_133 V123 V133 2.8862563800118807e-12
C123_133 V123 V133 4.221017180873511e-20

R123_134 V123 V134 -907.6786398852043
L123_134 V123 V134 4.248443380324692e-12
C123_134 V123 V134 -7.296566335680128e-21

R123_135 V123 V135 286.51728816128605
L123_135 V123 V135 -4.010230285156114e-12
C123_135 V123 V135 -3.143130363533467e-20

R123_136 V123 V136 987.9291875764353
L123_136 V123 V136 1.6572243337877748e-10
C123_136 V123 V136 -2.3678054958474267e-21

R123_137 V123 V137 -1310.8582985367564
L123_137 V123 V137 3.969047358971919e-12
C123_137 V123 V137 -2.680274382691353e-21

R123_138 V123 V138 -219.51341395293488
L123_138 V123 V138 7.087995440413472e-13
C123_138 V123 V138 -6.674899004353521e-20

R123_139 V123 V139 147.24293760396432
L123_139 V123 V139 -2.9026859494577755e-12
C123_139 V123 V139 -4.74586291939435e-21

R123_140 V123 V140 -1134.23433768689
L123_140 V123 V140 5.200278737957857e-12
C123_140 V123 V140 -1.0107762354035283e-20

R123_141 V123 V141 -360.524955522741
L123_141 V123 V141 1.2793944371772193e-11
C123_141 V123 V141 -2.6815218699375285e-20

R123_142 V123 V142 4464.794702783155
L123_142 V123 V142 9.753551502819581e-13
C123_142 V123 V142 -9.806277938153695e-20

R123_143 V123 V143 -708.0628611207745
L123_143 V123 V143 3.6196167539915443e-12
C123_143 V123 V143 -1.9902581533055837e-20

R123_144 V123 V144 1356.1187973309131
L123_144 V123 V144 -5.162047774187861e-12
C123_144 V123 V144 -6.772728052853908e-21

R124_124 V124 0 -731.645282055768
L124_124 V124 0 -9.49431546690314e-13
C124_124 V124 0 4.2152878734831714e-19

R124_125 V124 V125 -739.5015813946059
L124_125 V124 V125 1.5602170090647828e-12
C124_125 V124 V125 -3.997706508495596e-20

R124_126 V124 V126 858.0276868290481
L124_126 V124 V126 1.511651826794729e-11
C124_126 V124 V126 1.0824054858188181e-20

R124_127 V124 V127 -1656.0333685049995
L124_127 V124 V127 4.733074102830253e-12
C124_127 V124 V127 -3.543152644422214e-20

R124_128 V124 V128 1788.415269227211
L124_128 V124 V128 1.0008484959943404e-12
C124_128 V124 V128 1.07315077028915e-20

R124_129 V124 V129 -365.1516144491053
L124_129 V124 V129 -1.6111224235144354e-12
C124_129 V124 V129 -5.829081046021014e-20

R124_130 V124 V130 342.80736637626114
L124_130 V124 V130 1.556181964509238e-12
C124_130 V124 V130 -6.246800266110664e-20

R124_131 V124 V131 381.03374652503715
L124_131 V124 V131 1.1949300371153356e-12
C124_131 V124 V131 7.077416053572675e-20

R124_132 V124 V132 4597.205619970507
L124_132 V124 V132 -1.509145161770435e-11
C124_132 V124 V132 -7.915609621173425e-20

R124_133 V124 V133 2726.918187798434
L124_133 V124 V133 1.4561440575323206e-12
C124_133 V124 V133 1.6000771352328594e-19

R124_134 V124 V134 -4800878.427604393
L124_134 V124 V134 1.7032042704734447e-11
C124_134 V124 V134 -8.010465145091256e-21

R124_135 V124 V135 -1681.1687973634841
L124_135 V124 V135 8.546977568028119e-11
C124_135 V124 V135 -5.589778340423226e-20

R124_136 V124 V136 1848.1972420544566
L124_136 V124 V136 1.7964561235746955e-12
C124_136 V124 V136 -3.8920074567028504e-20

R124_137 V124 V137 -947.4474381262668
L124_137 V124 V137 6.921649882080057e-12
C124_137 V124 V137 -9.618299689752694e-20

R124_138 V124 V138 384.7394732794946
L124_138 V124 V138 2.040601600929174e-12
C124_138 V124 V138 -7.292121872610188e-20

R124_139 V124 V139 -1320.426951809007
L124_139 V124 V139 2.4610116772862072e-12
C124_139 V124 V139 2.2153544491061282e-20

R124_140 V124 V140 1623.191353665085
L124_140 V124 V140 2.1278559951345276e-12
C124_140 V124 V140 -6.563261325230364e-20

R124_141 V124 V141 -997.9883754476865
L124_141 V124 V141 -1.5655983816786968e-12
C124_141 V124 V141 1.4819210975347138e-20

R124_142 V124 V142 363.212034862074
L124_142 V124 V142 2.091922049632291e-12
C124_142 V124 V142 -1.0845334781159558e-19

R124_143 V124 V143 856.1615284603146
L124_143 V124 V143 2.0771185159053686e-11
C124_143 V124 V143 -3.7088620860485293e-20

R124_144 V124 V144 -10169.936284341566
L124_144 V124 V144 -5.465596231499398e-12
C124_144 V124 V144 4.69352117398209e-20

R125_125 V125 0 -63.07448898599216
L125_125 V125 0 1.887463571240719e-13
C125_125 V125 0 8.996429909930275e-19

R125_126 V125 V126 -295.27225678770606
L125_126 V125 V126 -1.8242843239913704e-12
C125_126 V125 V126 -2.4117717923968242e-20

R125_127 V125 V127 222.40618163823595
L125_127 V125 V127 -2.7682164005860615e-12
C125_127 V125 V127 1.651564568900151e-20

R125_128 V125 V128 1538.082809335135
L125_128 V125 V128 -3.4258598136637547e-12
C125_128 V125 V128 -1.105280499483454e-20

R125_129 V125 V129 822.2421105467473
L125_129 V125 V129 1.3626573170152432e-11
C125_129 V125 V129 7.448904304299156e-20

R125_130 V125 V130 -1173.5325854631894
L125_130 V125 V130 -1.4538120692013345e-12
C125_130 V125 V130 -9.101717864327113e-20

R125_131 V125 V131 -12606.202834340398
L125_131 V125 V131 -1.2392219064042334e-12
C125_131 V125 V131 2.6527593504516684e-21

R125_132 V125 V132 -2122.2960512177374
L125_132 V125 V132 -3.658030141605545e-12
C125_132 V125 V132 4.7771567897741394e-21

R125_133 V125 V133 581.948296609956
L125_133 V125 V133 -1.5141029599656075e-12
C125_133 V125 V133 6.264337940557601e-20

R125_134 V125 V134 1442.4684248991693
L125_134 V125 V134 -1.6749394268753394e-12
C125_134 V125 V134 -7.3112760915307e-20

R125_135 V125 V135 372.9196279848694
L125_135 V125 V135 -8.112938724006405e-12
C125_135 V125 V135 -3.6237119103846306e-20

R125_136 V125 V136 1437.944627757593
L125_136 V125 V136 -2.971224462387204e-12
C125_136 V125 V136 1.615762203237005e-20

R125_137 V125 V137 238.04115893739737
L125_137 V125 V137 -5.715210574999313e-13
C125_137 V125 V137 3.3019797852588957e-20

R125_138 V125 V138 -557.9710912187131
L125_138 V125 V138 -9.018141612569963e-13
C125_138 V125 V138 3.117764122109091e-20

R125_139 V125 V139 169.16429748613612
L125_139 V125 V139 -1.967054565977971e-12
C125_139 V125 V139 2.4204737534037072e-20

R125_140 V125 V140 -32040.964142212244
L125_140 V125 V140 -1.2443615314918607e-12
C125_140 V125 V140 -1.655000628287912e-20

R125_141 V125 V141 -3402.872973427739
L125_141 V125 V141 -1.1635692057439923e-11
C125_141 V125 V141 -2.0027787887640964e-20

R125_142 V125 V142 -1007.6254493256301
L125_142 V125 V142 -1.9128547906629034e-12
C125_142 V125 V142 1.3134163825757502e-20

R125_143 V125 V143 -401.5738506901901
L125_143 V125 V143 4.265140706783049e-12
C125_143 V125 V143 -9.614718337250722e-20

R125_144 V125 V144 -1503.284502985704
L125_144 V125 V144 2.1395778712953687e-12
C125_144 V125 V144 -8.397399755128659e-20

R126_126 V126 0 27.29368067534396
L126_126 V126 0 4.165547661387291e-13
C126_126 V126 0 5.428511928406385e-19

R126_127 V126 V127 -32.59624027168583
L126_127 V126 V127 3.9890181561937416e-13
C126_127 V126 V127 -1.5702786638904164e-21

R126_128 V126 V128 -425.6761265438653
L126_128 V126 V128 -2.3791433847573903e-11
C126_128 V126 V128 1.9372573304145185e-21

R126_129 V126 V129 -85.08643225883377
L126_129 V126 V129 8.101419432361309e-13
C126_129 V126 V129 6.150346377157639e-20

R126_130 V126 V130 118.61006220135486
L126_130 V126 V130 -5.210232997094329e-13
C126_130 V126 V130 9.611553471991226e-20

R126_131 V126 V131 92.069255892473
L126_131 V126 V131 -2.421602278280391e-12
C126_131 V126 V131 -9.868317757665144e-20

R126_132 V126 V132 127.12749361977306
L126_132 V126 V132 -1.4948463217768745e-12
C126_132 V126 V132 -6.638325726014627e-21

R126_133 V126 V133 418.66872487248355
L126_133 V126 V133 -1.9661679415471877e-11
C126_133 V126 V133 -1.464053849882863e-19

R126_134 V126 V134 167.6754051826866
L126_134 V126 V134 -1.966498797912174e-12
C126_134 V126 V134 -1.3145849576632898e-20

R126_135 V126 V135 -47.04499691923191
L126_135 V126 V135 7.15129751513924e-13
C126_135 V126 V135 -2.1320227259594904e-20

R126_136 V126 V136 -4340.047935134725
L126_136 V126 V136 -6.717300272785253e-12
C126_136 V126 V136 9.694412562511365e-21

R126_137 V126 V137 -4928.068772959778
L126_137 V126 V137 -2.899010446278322e-12
C126_137 V126 V137 8.322312825750948e-20

R126_138 V126 V138 28.61713993509375
L126_138 V126 V138 -3.0743615519401176e-13
C126_138 V126 V138 7.794026084813414e-20

R126_139 V126 V139 -25.46868615679002
L126_139 V126 V139 2.955649239530087e-13
C126_139 V126 V139 -6.219805878288273e-20

R126_140 V126 V140 94.8832493813672
L126_140 V126 V140 -7.242028916005675e-13
C126_140 V126 V140 5.189164891746346e-20

R126_141 V126 V141 131.68740670505744
L126_141 V126 V141 -1.6135735408377289e-12
C126_141 V126 V141 -5.067285145729403e-22

R126_142 V126 V142 95.19728959962559
L126_142 V126 V142 -6.914626188656589e-13
C126_142 V126 V142 2.1918519382024403e-21

R126_143 V126 V143 78.20073277366508
L126_143 V126 V143 -7.612755513993222e-13
C126_143 V126 V143 -5.456784539037098e-20

R126_144 V126 V144 -173.14114102463537
L126_144 V126 V144 1.115358813317931e-12
C126_144 V126 V144 -4.65573241119391e-20

R127_127 V127 0 -32.639449414646826
L127_127 V127 0 -1.0519378346224136e-12
C127_127 V127 0 1.1666378117394718e-19

R127_128 V127 V128 739.9974752792004
L127_128 V127 V128 1.111253312632329e-11
C127_128 V127 V128 9.188283992716971e-21

R127_129 V127 V129 107.92872225008253
L127_129 V127 V129 -1.4604630145831065e-12
C127_129 V127 V129 -2.4688488969406213e-20

R127_130 V127 V130 -145.27978214963267
L127_130 V127 V130 8.20018627307269e-13
C127_130 V127 V130 1.6320754640933066e-20

R127_131 V127 V131 -118.83526687618084
L127_131 V127 V131 -9.37948839659876e-12
C127_131 V127 V131 4.344619522150854e-20

R127_132 V127 V132 -171.7348367684339
L127_132 V127 V132 1.9757078550236757e-12
C127_132 V127 V132 -1.035166373071114e-20

R127_133 V127 V133 -681.2174988610813
L127_133 V127 V133 -2.5013490510023538e-12
C127_133 V127 V133 -5.189953142765945e-21

R127_134 V127 V134 -244.66133569536393
L127_134 V127 V134 5.053463252786668e-12
C127_134 V127 V134 2.4322526071227678e-21

R127_135 V127 V135 62.458665543814625
L127_135 V127 V135 -7.656069352242205e-13
C127_135 V127 V135 8.879042686054195e-21

R127_136 V127 V136 28061.903857730063
L127_136 V127 V136 3.045842662761844e-11
C127_136 V127 V136 -1.4073533238556996e-20

R127_137 V127 V137 774.9557640133544
L127_137 V127 V137 -1.5350458250448295e-11
C127_137 V127 V137 -1.016384610775315e-20

R127_138 V127 V138 -38.42149035367946
L127_138 V127 V138 4.5374172949463775e-13
C127_138 V127 V138 -4.754705954899382e-20

R127_139 V127 V139 33.73977938008258
L127_139 V127 V139 -3.17893678658721e-13
C127_139 V127 V139 -1.6224590142105875e-20

R127_140 V127 V140 -126.99741197391579
L127_140 V127 V140 9.045104301198843e-13
C127_140 V127 V140 1.1063468612817687e-20

R127_141 V127 V141 -194.70043478606604
L127_141 V127 V141 1.9003931596663054e-12
C127_141 V127 V141 -1.5365334679321093e-21

R127_142 V127 V142 -120.0138499930882
L127_142 V127 V142 1.2842458147235852e-12
C127_142 V127 V142 -3.072232919540055e-20

R127_143 V127 V143 -99.94215177920879
L127_143 V127 V143 9.192061418080078e-13
C127_143 V127 V143 -3.1459121940679098e-21

R127_144 V127 V144 243.79538796874553
L127_144 V127 V144 -1.5656491597227025e-12
C127_144 V127 V144 1.8955988591940698e-20

R128_128 V128 0 -400.96530140612003
L128_128 V128 0 7.711111025131399e-13
C128_128 V128 0 1.9486834139562096e-20

R128_129 V128 V129 430.03383014026934
L128_129 V128 V129 1.843623674648577e-10
C128_129 V128 V129 -3.5212283079464465e-20

R128_130 V128 V130 -431.66033641446404
L128_130 V128 V130 -3.5524928955939045e-12
C128_130 V128 V130 -9.846469558683515e-20

R128_131 V128 V131 -434.21489700132327
L128_131 V128 V131 -6.714951430410302e-12
C128_131 V128 V131 -2.8731807258854933e-21

R128_132 V128 V132 -2253.4040666986934
L128_132 V128 V132 -5.486485983290737e-12
C128_132 V128 V132 -7.710144554554478e-20

R128_133 V128 V133 -3122.7224815754253
L128_133 V128 V133 -4.462234512938569e-12
C128_133 V128 V133 7.973283663780802e-20

R128_134 V128 V134 -3261.5250802691307
L128_134 V128 V134 2.1191621271386e-11
C128_134 V128 V134 1.3038120129604887e-20

R128_135 V128 V135 885.9370142187904
L128_135 V128 V135 2.3470996796385845e-10
C128_135 V128 V135 -1.7206937878130547e-20

R128_136 V128 V136 101748.25077331763
L128_136 V128 V136 -1.7791272944798071e-12
C128_136 V128 V136 1.1583341423177655e-19

R128_137 V128 V137 2696.097574101508
L128_137 V128 V137 -3.9901347335064805e-11
C128_137 V128 V137 -2.4693613826174733e-20

R128_138 V128 V138 -302.1312132975736
L128_138 V128 V138 9.41570775657918e-12
C128_138 V128 V138 4.943987571385973e-20

R128_139 V128 V139 545.610192720835
L128_139 V128 V139 -3.285406139257189e-11
C128_139 V128 V139 4.213025890189354e-20

R128_140 V128 V140 -2280.800476515678
L128_140 V128 V140 -1.5341406783802188e-12
C128_140 V128 V140 5.666544771075716e-20

R128_141 V128 V141 -48714.03768547344
L128_141 V128 V141 1.1359014959271158e-12
C128_141 V128 V141 2.1602228953107208e-20

R128_142 V128 V142 -436.90899254009446
L128_142 V128 V142 -1.0951886571335135e-11
C128_142 V128 V142 -3.9422548416284886e-20

R128_143 V128 V143 -867.7005939489338
L128_143 V128 V143 -1.1329255481032973e-11
C128_143 V128 V143 9.60008556059495e-21

R128_144 V128 V144 5396.1061118196085
L128_144 V128 V144 4.376008419885926e-12
C128_144 V128 V144 -4.98441379021583e-20

R129_129 V129 0 -57.232808846057445
L129_129 V129 0 -4.4258436338135803e-13
C129_129 V129 0 -3.735064793515701e-19

R129_130 V129 V130 2061.5613972381852
L129_130 V129 V130 6.329050249806787e-13
C129_130 V129 V130 -4.207184303482462e-20

R129_131 V129 V131 -1888.513857801613
L129_131 V129 V131 8.617725653287569e-13
C129_131 V129 V131 6.962619485470388e-20

R129_132 V129 V132 -456.5326350651985
L129_132 V129 V132 9.220457159551069e-12
C129_132 V129 V132 -5.778431783361906e-20

R129_133 V129 V133 44881.896154897935
L129_133 V129 V133 4.76377188267751e-12
C129_133 V129 V133 5.834506656542165e-20

R129_134 V129 V134 -620.3847869904956
L129_134 V129 V134 9.22895834448926e-12
C129_134 V129 V134 6.616393406796912e-20

R129_135 V129 V135 160.8483935047809
L129_135 V129 V135 -1.8875423828535076e-12
C129_135 V129 V135 7.894383814762894e-22

R129_136 V129 V136 845.0073554423867
L129_136 V129 V136 5.198275544070534e-12
C129_136 V129 V136 1.8792233164113106e-20

R129_137 V129 V137 -2802.8877607356662
L129_137 V129 V137 -5.204903799331075e-12
C129_137 V129 V137 -5.78842322709171e-20

R129_138 V129 V138 -123.30828427103619
L129_138 V129 V138 6.058449986596765e-13
C129_138 V129 V138 -8.221547712763672e-20

R129_139 V129 V139 83.52141482325268
L129_139 V129 V139 -1.11857226974459e-12
C129_139 V129 V139 1.8734029965117407e-20

R129_140 V129 V140 -483.2199057218082
L129_140 V129 V140 1.8030792252578372e-12
C129_140 V129 V140 -1.166843454562842e-20

R129_141 V129 V141 -259.63175895198685
L129_141 V129 V141 -3.152367819149252e-11
C129_141 V129 V141 1.0584000192754433e-20

R129_142 V129 V142 -2961.006569923779
L129_142 V129 V142 8.26885735106389e-13
C129_142 V129 V142 -1.2013815258179712e-19

R129_143 V129 V143 -337.8194766674509
L129_143 V129 V143 1.2863540278223776e-12
C129_143 V129 V143 6.34226925160801e-20

R129_144 V129 V144 754.2654914406452
L129_144 V129 V144 -6.167146955188008e-12
C129_144 V129 V144 6.986870312446653e-20

R130_130 V130 0 77.27021724334291
L130_130 V130 0 4.1830526366245266e-13
C130_130 V130 0 1.3255335817270924e-20

R130_131 V130 V131 -1345.9329519447842
L130_131 V130 V131 -8.323532544055787e-13
C130_131 V130 V131 1.338998705211174e-19

R130_132 V130 V132 654.0805838183107
L130_132 V130 V132 -1.926344174403047e-12
C130_132 V130 V132 -6.320022359707667e-20

R130_133 V130 V133 -4595.713637589134
L130_133 V130 V133 -9.228029620831917e-12
C130_133 V130 V133 3.024535409627094e-19

R130_134 V130 V134 779.9507274925455
L130_134 V130 V134 -2.0678290753417435e-12
C130_134 V130 V134 8.501470003536997e-21

R130_135 V130 V135 -219.59040162808287
L130_135 V130 V135 1.272219718432026e-12
C130_135 V130 V135 -8.041986777808193e-20

R130_136 V130 V136 -763.9183162228201
L130_136 V130 V136 -7.477203795726095e-12
C130_136 V130 V136 9.976667855350771e-20

R130_137 V130 V137 2631.3151872089707
L130_137 V130 V137 -2.490609794316176e-12
C130_137 V130 V137 -1.4302399055323313e-19

R130_138 V130 V138 201.95344506587813
L130_138 V130 V138 -3.693088182312481e-13
C130_138 V130 V138 1.868822605276162e-20

R130_139 V130 V139 -112.72141867725533
L130_139 V130 V139 5.567408138235815e-13
C130_139 V130 V139 1.5119127941160998e-19

R130_140 V130 V140 914.9299541373002
L130_140 V130 V140 -1.0140461496057492e-12
C130_140 V130 V140 -4.49926657257407e-20

R130_141 V130 V141 292.27101949438486
L130_141 V130 V141 3.0755250172019385e-11
C130_141 V130 V141 2.3959846753983947e-20

R130_142 V130 V142 -999.9533677800538
L130_142 V130 V142 -5.542258955061541e-13
C130_142 V130 V142 -6.161581662004559e-20

R130_143 V130 V143 553.5837643894309
L130_143 V130 V143 -1.2427694407563652e-12
C130_143 V130 V143 2.0490861822853694e-20

R130_144 V130 V144 -1238.3928705317135
L130_144 V130 V144 1.8432485101919336e-12
C130_144 V130 V144 -2.216633355501331e-20

R131_131 V131 0 75.95542348243275
L131_131 V131 0 1.6158267444075837e-12
C131_131 V131 0 -3.2019205453005523e-19

R131_132 V131 V132 484.96707475485766
L131_132 V131 V132 -2.1679668460975624e-11
C131_132 V131 V132 1.697078013211631e-20

R131_133 V131 V133 7637.2941182549885
L131_133 V131 V133 -1.917619212601137e-12
C131_133 V131 V133 -7.327211372147443e-20

R131_134 V131 V134 577.8036055568894
L131_134 V131 V134 -3.6294196761886043e-12
C131_134 V131 V134 -4.666631942746191e-20

R131_135 V131 V135 -177.61690540115953
L131_135 V131 V135 -2.221562281012573e-11
C131_135 V131 V135 3.6071763293133365e-20

R131_136 V131 V136 -881.6504823072044
L131_136 V131 V136 -4.687915798237944e-12
C131_136 V131 V136 3.010731112612948e-20

R131_137 V131 V137 1144.5716917969553
L131_137 V131 V137 -5.498085289644519e-12
C131_137 V131 V137 8.033042746048146e-20

R131_138 V131 V138 133.22589015049218
L131_138 V131 V138 -9.58431072373093e-13
C131_138 V131 V138 1.7529946383483748e-19

R131_139 V131 V139 -91.84216925764134
L131_139 V131 V139 -5.395437973557472e-12
C131_139 V131 V139 -5.3456112943947306e-20

R131_140 V131 V140 514.6078757728951
L131_140 V131 V140 -3.3664979404122467e-12
C131_140 V131 V140 3.5324534555699155e-20

R131_141 V131 V141 265.1700052442488
L131_141 V131 V141 3.8906545904183845e-12
C131_141 V131 V141 2.9373825936789736e-20

R131_142 V131 V142 11939.731851605224
L131_142 V131 V142 -1.0058883888630734e-12
C131_142 V131 V142 1.1835647604308005e-19

R131_143 V131 V143 398.4707286020956
L131_143 V131 V143 -3.986716765100038e-12
C131_143 V131 V143 -3.470742238589942e-21

R131_144 V131 V144 -748.2529729573895
L131_144 V131 V144 8.475015338013543e-12
C131_144 V131 V144 -6.229872976080987e-20

R132_132 V132 0 130.25736098481332
L132_132 V132 0 8.624631701149479e-13
C132_132 V132 0 2.4073655720262743e-19

R132_133 V132 V133 1962.0998797036914
L132_133 V132 V133 -8.580011619288175e-10
C132_133 V132 V133 6.508254170734862e-22

R132_134 V132 V134 871.4048564126374
L132_134 V132 V134 -1.3705140503757822e-11
C132_134 V132 V134 3.816447800448922e-20

R132_135 V132 V135 -247.0168994211225
L132_135 V132 V135 3.8827045485475026e-12
C132_135 V132 V135 -3.7640844806990006e-20

R132_136 V132 V136 97492.73225784344
L132_136 V132 V136 1.0999794061180315e-11
C132_136 V132 V136 1.1807613563398355e-19

R132_137 V132 V137 22326.333904769304
L132_137 V132 V137 -4.749600672748081e-12
C132_137 V132 V137 -1.624862659778909e-20

R132_138 V132 V138 150.25849807440483
L132_138 V132 V138 -1.413340953930948e-12
C132_138 V132 V138 -2.3320638464659767e-21

R132_139 V132 V139 -134.71036391622062
L132_139 V132 V139 1.3613180105436865e-12
C132_139 V132 V139 2.208595031239238e-20

R132_140 V132 V140 510.2247676011979
L132_140 V132 V140 -2.7737358883879476e-12
C132_140 V132 V140 4.082638079085486e-20

R132_141 V132 V141 638.3325687967678
L132_141 V132 V141 -1.4998092020178535e-11
C132_141 V132 V141 6.47512443724684e-21

R132_142 V132 V142 518.8423566426493
L132_142 V132 V142 -2.8188127695230576e-12
C132_142 V132 V142 -6.551360840383928e-20

R132_143 V132 V143 419.60948460809783
L132_143 V132 V143 -4.465371378131969e-12
C132_143 V132 V143 -1.300662019860926e-21

R132_144 V132 V144 -890.774472897497
L132_144 V132 V144 3.96490731524933e-12
C132_144 V132 V144 -4.3292985833818976e-20

R133_133 V133 0 559.0390941746206
L133_133 V133 0 8.488177271326878e-13
C133_133 V133 0 1.017276503199156e-18

R133_134 V133 V134 1564.396815465782
L133_134 V133 V134 -3.1936098235677914e-11
C133_134 V133 V134 4.62041753204351e-20

R133_135 V133 V135 -938.5767639047244
L133_135 V133 V135 -6.333077504865537e-12
C133_135 V133 V135 2.898659046589549e-20

R133_136 V133 V136 -10202.902817809812
L133_136 V133 V136 -3.6035072253466726e-12
C133_136 V133 V136 -1.8958921884841038e-20

R133_137 V133 V137 863.9269479890849
L133_137 V133 V137 -2.0256329342625096e-10
C133_137 V133 V137 3.0601280409545955e-19

R133_138 V133 V138 544.6393489399667
L133_138 V133 V138 -3.075372043401129e-12
C133_138 V133 V138 -1.889246417024577e-20

R133_139 V133 V139 -533.3979348422513
L133_139 V133 V139 -1.570910607743436e-12
C133_139 V133 V139 -1.688283388319119e-19

R133_140 V133 V140 1566.9063344056399
L133_140 V133 V140 -9.707256095387263e-12
C133_140 V133 V140 6.900693687391928e-20

R133_141 V133 V141 1114.8166614796253
L133_141 V133 V141 6.597724437813904e-12
C133_141 V133 V141 -2.933036126477653e-20

R133_142 V133 V142 -25505.54954246339
L133_142 V133 V142 -5.363198150891265e-12
C133_142 V133 V142 2.832765669485856e-20

R133_143 V133 V143 4019.6208344369547
L133_143 V133 V143 -4.994313438480868e-11
C133_143 V133 V143 -6.794024624924869e-20

R133_144 V133 V144 -1730.0394695752077
L133_144 V133 V144 8.890787319479125e-11
C133_144 V133 V144 -6.592024892709994e-20

R134_134 V134 0 145.9367275710814
L134_134 V134 0 4.7303877513992e-13
C134_134 V134 0 4.482503921533006e-19

R134_135 V134 V135 -343.4353239591457
L134_135 V134 V135 3.995618406508145e-12
C134_135 V134 V135 3.3735584790193375e-20

R134_136 V134 V136 16324.356661293434
L134_136 V134 V136 -5.935615160367535e-10
C134_136 V134 V136 -7.167927454490991e-21

R134_137 V134 V137 1575.8286634956498
L134_137 V134 V137 -4.752155499586019e-12
C134_137 V134 V137 3.9599445943161255e-20

R134_138 V134 V138 191.93271366505817
L134_138 V134 V138 -1.8433251470393853e-12
C134_138 V134 V138 3.3450345318642084e-20

R134_139 V134 V139 -192.0158274954777
L134_139 V134 V139 3.639565790972891e-12
C134_139 V134 V139 -1.4792363914159728e-20

R134_140 V134 V140 624.8708435847152
L134_140 V134 V140 -2.7599912442993593e-12
C134_140 V134 V140 -8.477949114014401e-21

R134_141 V134 V141 829.5166810877085
L134_141 V134 V141 -5.561403982452126e-12
C134_141 V134 V141 8.475445343139759e-22

R134_142 V134 V142 675.5029836317019
L134_142 V134 V142 -4.383299418138308e-12
C134_142 V134 V142 6.397919644644339e-20

R134_143 V134 V143 617.9219399467173
L134_143 V134 V143 -4.506932133916033e-12
C134_143 V134 V143 -4.5418032702456654e-20

R134_144 V134 V144 -977.9013209932237
L134_144 V134 V144 5.1574256668952617e-11
C134_144 V134 V144 -6.482944353880622e-20

R135_135 V135 0 -49.736587537121835
L135_135 V135 0 -3.8398245782140906e-12
C135_135 V135 0 3.2894122603240724e-19

R135_136 V135 V136 9087.061139980604
L135_136 V135 V136 1.3014790489643166e-11
C135_136 V135 V136 1.5110257021624694e-20

R135_137 V135 V137 1590.0191355012892
L135_137 V135 V137 -3.8975159083857903e-10
C135_137 V135 V137 -4.1181134152114624e-20

R135_138 V135 V138 -55.68464162857914
L135_138 V135 V138 6.627590651570651e-13
C135_138 V135 V138 2.5867644928798227e-21

R135_139 V135 V139 48.72002376572903
L135_139 V135 V139 -5.741085889859002e-13
C135_139 V135 V139 6.907842185872682e-20

R135_140 V135 V140 -184.97503522532355
L135_140 V135 V140 1.5280393633818832e-12
C135_140 V135 V140 -6.272661306070537e-22

R135_141 V135 V141 -266.0182619858349
L135_141 V135 V141 3.4715232313643203e-12
C135_141 V135 V141 -9.77080315228006e-21

R135_142 V135 V142 -179.20085180816312
L135_142 V135 V142 1.7877698790270691e-12
C135_142 V135 V142 -5.71462538940976e-20

R135_143 V135 V143 -147.12266869016526
L135_143 V135 V143 1.6029672279894534e-12
C135_143 V135 V143 3.3802593572897445e-22

R135_144 V135 V144 349.58598254054107
L135_144 V135 V144 -2.3969912655629264e-12
C135_144 V135 V144 9.460105609617907e-23

R136_136 V136 0 -2436.468333102485
L136_136 V136 0 9.481564201447606e-13
C136_136 V136 0 -1.7791418555541253e-19

R136_137 V136 V137 2081.1945526241593
L136_137 V136 V137 -9.431139185700036e-12
C136_137 V136 V137 -1.9125180012414236e-20

R136_138 V136 V138 -1035.0684300135597
L136_138 V136 V138 -2.818465185353978e-12
C136_138 V136 V138 -6.260516162551285e-20

R136_139 V136 V139 10471.122536499372
L136_139 V136 V139 -1.0080751449373467e-11
C136_139 V136 V139 -3.5127168193478375e-20

R136_140 V136 V140 -40359.23477560839
L136_140 V136 V140 -1.8138956906534905e-12
C136_140 V136 V140 -8.313379482180849e-20

R136_141 V136 V141 2820.7662279850474
L136_141 V136 V141 2.9710678076879e-12
C136_141 V136 V141 -2.352563890656111e-20

R136_142 V136 V142 -804.4718896071046
L136_142 V136 V142 -5.16643137776083e-12
C136_142 V136 V142 2.5179621404957144e-20

R136_143 V136 V143 -2286.8639778287893
L136_143 V136 V143 -1.2298317886628067e-11
C136_143 V136 V143 -1.7689419555119356e-22

R136_144 V136 V144 -16242.852345486208
L136_144 V136 V144 2.731688381927541e-12
C136_144 V136 V144 1.1627627805582582e-19

R137_137 V137 0 -106.02633453040055
L137_137 V137 0 2.5111708314849802e-12
C137_137 V137 0 -8.1204194082672835e-19

R137_138 V137 V138 1302.4850867169018
L137_138 V137 V138 -1.393110526760292e-12
C137_138 V137 V138 -2.123440863893389e-21

R137_139 V137 V139 567.0149597843243
L137_139 V137 V139 1.0423093050015485e-10
C137_139 V137 V139 9.08960986491445e-20

R137_140 V137 V140 2067.3395910302447
L137_140 V137 V140 -1.9046646766275093e-12
C137_140 V137 V140 -6.819459284614422e-20

R137_141 V137 V141 -9953.85851651637
L137_141 V137 V141 -4.215820750066674e-12
C137_141 V137 V141 -1.198071025047849e-20

R137_142 V137 V142 2637.002488380925
L137_142 V137 V142 -3.5325201736348605e-12
C137_142 V137 V142 -4.4232686534868226e-20

R137_143 V137 V143 -1454.2702504166687
L137_143 V137 V143 2.768713450499181e-12
C137_143 V137 V143 8.586738825282009e-20

R137_144 V137 V144 -1712.7035447761612
L137_144 V137 V144 1.8590458739497414e-12
C137_144 V137 V144 9.794648415235502e-20

R138_138 V138 0 29.745731490946017
L138_138 V138 0 3.6062031637932426e-13
C138_138 V138 0 5.819520743534201e-19

R138_139 V138 V139 -29.933510892502998
L138_139 V138 V139 3.197146693970391e-13
C138_139 V138 V139 -1.9220278884129203e-20

R138_140 V138 V140 121.40800770923536
L138_140 V138 V140 -5.982795937162521e-13
C138_140 V138 V140 -5.697951260091013e-20

R138_141 V138 V141 128.7728647502174
L138_141 V138 V141 -1.5598451559574783e-12
C138_141 V138 V141 -5.834660570524967e-20

R138_142 V138 V142 142.80183237653648
L138_142 V138 V142 -4.3992348458208757e-13
C138_142 V138 V142 -1.0386916470945673e-19

R138_143 V138 V143 99.26404086643305
L138_143 V138 V143 -8.157663734701766e-13
C138_143 V138 V143 1.575345707484835e-20

R138_144 V138 V144 -209.34380711447182
L138_144 V138 V144 8.739315390882233e-13
C138_144 V138 V144 6.25589329699507e-20

R139_139 V139 0 -24.70247327617
L139_139 V139 0 -8.78460913589763e-13
C139_139 V139 0 -2.7626761155045066e-20

R139_140 V139 V140 -99.86757411432804
L139_140 V139 V140 7.249835870597121e-13
C139_140 V139 V140 1.1703196236699935e-20

R139_141 V139 V141 -151.89855356343594
L139_141 V139 V141 1.255981174420621e-12
C139_141 V139 V141 -2.173471876977917e-21

R139_142 V139 V142 -93.33818690506523
L139_142 V139 V142 8.501017999844819e-13
C139_142 V139 V142 2.6342959681933233e-20

R139_143 V139 V143 -77.80905186998608
L139_143 V139 V143 7.422799106987648e-13
C139_143 V139 V143 -7.725999392746573e-20

R139_144 V139 V144 191.47792532110532
L139_144 V139 V144 -1.20392594748779e-12
C139_144 V139 V144 1.7553085899308565e-20

R140_140 V140 0 80.77037311601622
L140_140 V140 0 3.6908033018294263e-13
C140_140 V140 0 -2.839591107212548e-19

R140_141 V140 V141 442.9730039990277
L140_141 V140 V141 4.933641066898563e-12
C140_141 V140 V141 2.67636976718027e-20

R140_142 V140 V142 587.629821357127
L140_142 V140 V142 -1.4621165673757334e-12
C140_142 V140 V142 1.7075343559385672e-20

R140_143 V140 V143 344.2258959236817
L140_143 V140 V143 -2.103082032291315e-12
C140_143 V140 V143 1.7272543763962415e-20

R140_144 V140 V144 -621.3725192771402
L140_144 V140 V144 1.4631675103274672e-12
C140_144 V140 V144 3.3944502056837235e-20

R141_141 V141 0 370.3244678131836
L141_141 V141 0 -3.783500036417908e-12
C141_141 V141 0 3.056143576720609e-19

R141_142 V141 V142 271.95497987524374
L141_142 V141 V142 -2.66008124371028e-11
C141_142 V141 V142 -1.2692636256434318e-20

R141_143 V141 V143 368.67839692257513
L141_143 V141 V143 -1.2428989130326132e-11
C141_143 V141 V143 7.95391280080075e-21

R141_144 V141 V144 -863.3867491885983
L141_144 V141 V144 2.3842747707728683e-11
C141_144 V141 V144 -8.997395722334272e-21

R142_142 V142 0 56.99740471363452
L142_142 V142 0 3.6938967335627976e-13
C142_142 V142 0 2.550323157656514e-19

R142_143 V142 V143 395.86211237395406
L142_143 V142 V143 -1.6693095498198837e-12
C142_143 V142 V143 3.525790380154136e-20

R142_144 V142 V144 -859.1004343882959
L142_144 V142 V144 2.3500048616185198e-12
C142_144 V142 V144 2.4227897350025297e-21

R143_143 V143 0 65.6509181439905
L143_143 V143 0 7.517633994698873e-13
C143_143 V143 0 7.375687752077353e-19

R143_144 V143 V144 -659.1751284661063
L143_144 V143 V144 3.693503070205084e-12
C143_144 V143 V144 2.483854408238265e-21

R144_144 V144 0 -417.01554884665404
L144_144 V144 0 4.227167477077889e-12
C144_144 V144 0 1.235121313725904e-18

ISRC1_p1 0 V1  ac 6.346106463412155e-04*Ip1
ISRC1_p2 0 V1  ac 7.592674059024366e-05*Ip2
ISRC1_p3 0 V1  ac 1.100664147328153e-04*Ip3
ISRC1_p4 0 V1  ac 9.804084227331987e-05*Ip4

ISRC2_p1 0 V2  ac -1.275305890652397e-03*Ip1
ISRC2_p2 0 V2  ac 1.202874550473938e-03*Ip2
ISRC2_p3 0 V2  ac 1.959211508249852e-05*Ip3
ISRC2_p4 0 V2  ac 6.364076900024252e-05*Ip4

ISRC3_p1 0 V3  ac -1.304257337842080e-03*Ip1
ISRC3_p2 0 V3  ac -1.206250199988911e-03*Ip2
ISRC3_p3 0 V3  ac 2.526262024587809e-05*Ip3
ISRC3_p4 0 V3  ac -3.615441361394585e-04*Ip4

ISRC4_p1 0 V4  ac 1.110911742403385e-04*Ip1
ISRC4_p2 0 V4  ac 3.728878201374582e-05*Ip2
ISRC4_p3 0 V4  ac 5.466885091878189e-06*Ip3
ISRC4_p4 0 V4  ac 6.640204954207361e-03*Ip4

ISRC5_p1 0 V5  ac 6.743460732342449e-03*Ip1
ISRC5_p2 0 V5  ac 1.074536917181697e-03*Ip2
ISRC5_p3 0 V5  ac 8.642325052228133e-04*Ip3
ISRC5_p4 0 V5  ac 1.050391553673756e-03*Ip4

ISRC6_p1 0 V6  ac -1.537862538609469e-04*Ip1
ISRC6_p2 0 V6  ac 9.149431900296504e-03*Ip2
ISRC6_p3 0 V6  ac 1.414353189952099e-03*Ip3
ISRC6_p4 0 V6  ac 2.195135293225690e-03*Ip4

ISRC7_p1 0 V7  ac 2.787107199654842e-04*Ip1
ISRC7_p2 0 V7  ac -2.316464577597189e-03*Ip2
ISRC7_p3 0 V7  ac 4.032874966431459e-03*Ip3
ISRC7_p4 0 V7  ac 3.282022794234710e-04*Ip4

ISRC8_p1 0 V8  ac 2.320940118525939e-03*Ip1
ISRC8_p2 0 V8  ac 1.207446414350427e-03*Ip2
ISRC8_p3 0 V8  ac 1.595848213114707e-03*Ip3
ISRC8_p4 0 V8  ac 1.301486842096976e-02*Ip4

ISRC9_p1 0 V9  ac 2.965154378616991e-02*Ip1
ISRC9_p2 0 V9  ac 5.287684862158463e-03*Ip2
ISRC9_p3 0 V9  ac 7.486634618171250e-03*Ip3
ISRC9_p4 0 V9  ac 5.412467421761420e-03*Ip4

ISRC10_p1 0 V10  ac 9.975305582160940e-04*Ip1
ISRC10_p2 0 V10  ac 2.229375272502028e-02*Ip2
ISRC10_p3 0 V10  ac 2.830946861691208e-03*Ip3
ISRC10_p4 0 V10  ac 6.610407498910029e-03*Ip4

ISRC11_p1 0 V11  ac 8.818033552330637e-03*Ip1
ISRC11_p2 0 V11  ac -1.751789725563776e-02*Ip2
ISRC11_p3 0 V11  ac 4.108987713136609e-03*Ip3
ISRC11_p4 0 V11  ac 1.762948923339443e-03*Ip4

ISRC12_p1 0 V12  ac -4.318971470622608e-03*Ip1
ISRC12_p2 0 V12  ac -7.958549216422264e-03*Ip2
ISRC12_p3 0 V12  ac -2.405895762543746e-02*Ip3
ISRC12_p4 0 V12  ac 4.231076755660474e-02*Ip4

ISRC13_p1 0 V13  ac 2.914732835388200e-03*Ip1
ISRC13_p2 0 V13  ac 2.150854297432134e-03*Ip2
ISRC13_p3 0 V13  ac -7.744746461805463e-03*Ip3
ISRC13_p4 0 V13  ac -1.893583895175155e-02*Ip4

ISRC14_p1 0 V14  ac 8.649777724797063e-03*Ip1
ISRC14_p2 0 V14  ac 1.353824386312290e-02*Ip2
ISRC14_p3 0 V14  ac 3.150645817034577e-02*Ip3
ISRC14_p4 0 V14  ac 2.906644119593309e-02*Ip4

ISRC15_p1 0 V15  ac 9.041031201663422e-04*Ip1
ISRC15_p2 0 V15  ac -2.485963612920159e-04*Ip2
ISRC15_p3 0 V15  ac 1.322768928667090e-02*Ip3
ISRC15_p4 0 V15  ac 2.100744355413053e-02*Ip4

ISRC16_p1 0 V16  ac 9.992196397322784e-04*Ip1
ISRC16_p2 0 V16  ac 4.730526446118883e-03*Ip2
ISRC16_p3 0 V16  ac 4.641329949397410e-03*Ip3
ISRC16_p4 0 V16  ac 2.226279790373395e-02*Ip4

ISRC17_p1 0 V17  ac 1.991370518982710e-02*Ip1
ISRC17_p2 0 V17  ac 1.048430863111751e-02*Ip2
ISRC17_p3 0 V17  ac 1.258103341888880e-02*Ip3
ISRC17_p4 0 V17  ac 7.786582371754731e-03*Ip4

ISRC18_p1 0 V18  ac 2.989933299097533e-03*Ip1
ISRC18_p2 0 V18  ac 9.738624567410354e-03*Ip2
ISRC18_p3 0 V18  ac 8.600827392616801e-04*Ip3
ISRC18_p4 0 V18  ac -2.659265899017694e-03*Ip4

ISRC19_p1 0 V19  ac 1.402481180585170e-02*Ip1
ISRC19_p2 0 V19  ac -9.580875845916004e-04*Ip2
ISRC19_p3 0 V19  ac 3.246073021201043e-03*Ip3
ISRC19_p4 0 V19  ac 4.586094866247754e-03*Ip4

ISRC20_p1 0 V20  ac -2.675390794811799e-03*Ip1
ISRC20_p2 0 V20  ac -1.656764886876315e-03*Ip2
ISRC20_p3 0 V20  ac -2.812223952121029e-03*Ip3
ISRC20_p4 0 V20  ac -8.137444175390054e-03*Ip4

ISRC21_p1 0 V21  ac 7.900200553567568e-02*Ip1
ISRC21_p2 0 V21  ac 9.505750466625391e-03*Ip2
ISRC21_p3 0 V21  ac 1.191358026283119e-02*Ip3
ISRC21_p4 0 V21  ac 6.816548309257890e-03*Ip4

ISRC22_p1 0 V22  ac -1.146142664262965e-02*Ip1
ISRC22_p2 0 V22  ac 7.576751763997121e-02*Ip2
ISRC22_p3 0 V22  ac 8.693788141496911e-03*Ip3
ISRC22_p4 0 V22  ac 8.089292324472081e-03*Ip4

ISRC23_p1 0 V23  ac -1.083758565549345e-02*Ip1
ISRC23_p2 0 V23  ac -1.427067189839449e-02*Ip2
ISRC23_p3 0 V23  ac 8.131110901602316e-02*Ip3
ISRC23_p4 0 V23  ac -1.606511631788440e-03*Ip4

ISRC24_p1 0 V24  ac -6.836052403876650e-03*Ip1
ISRC24_p2 0 V24  ac -1.151700350296665e-02*Ip2
ISRC24_p3 0 V24  ac -6.564768001465768e-03*Ip3
ISRC24_p4 0 V24  ac 6.108923751892247e-02*Ip4

ISRC25_p1 0 V25  ac 3.519775238645972e-02*Ip1
ISRC25_p2 0 V25  ac -2.732140707386713e-03*Ip2
ISRC25_p3 0 V25  ac -7.434316581940417e-03*Ip3
ISRC25_p4 0 V25  ac -3.337844849974045e-03*Ip4

ISRC26_p1 0 V26  ac -3.727440782982116e-03*Ip1
ISRC26_p2 0 V26  ac 4.033829782695830e-02*Ip2
ISRC26_p3 0 V26  ac -4.903126625398302e-03*Ip3
ISRC26_p4 0 V26  ac -5.211121754744218e-03*Ip4

ISRC27_p1 0 V27  ac 1.193767612179376e-04*Ip1
ISRC27_p2 0 V27  ac 8.028182528241872e-03*Ip2
ISRC27_p3 0 V27  ac 2.203545513371015e-02*Ip3
ISRC27_p4 0 V27  ac -5.361801686161956e-03*Ip4

ISRC28_p1 0 V28  ac 3.010248660111186e-04*Ip1
ISRC28_p2 0 V28  ac 5.066074477169142e-03*Ip2
ISRC28_p3 0 V28  ac 5.829226268677232e-03*Ip3
ISRC28_p4 0 V28  ac 3.924995420787877e-02*Ip4

ISRC29_p1 0 V29  ac 3.499269520234437e-02*Ip1
ISRC29_p2 0 V29  ac -7.728875645331933e-04*Ip2
ISRC29_p3 0 V29  ac -4.416370510730337e-03*Ip3
ISRC29_p4 0 V29  ac -3.401384426574232e-03*Ip4

ISRC30_p1 0 V30  ac -5.364831527585583e-03*Ip1
ISRC30_p2 0 V30  ac 3.068270053413872e-02*Ip2
ISRC30_p3 0 V30  ac -2.338424947961174e-03*Ip3
ISRC30_p4 0 V30  ac -2.020578206679665e-04*Ip4

ISRC31_p1 0 V31  ac -9.643038190517147e-03*Ip1
ISRC31_p2 0 V31  ac -1.205529644405060e-02*Ip2
ISRC31_p3 0 V31  ac 2.608104444626582e-02*Ip3
ISRC31_p4 0 V31  ac -4.927180250174206e-03*Ip4

ISRC32_p1 0 V32  ac -3.466932315628427e-03*Ip1
ISRC32_p2 0 V32  ac -5.863979955056444e-03*Ip2
ISRC32_p3 0 V32  ac -4.091889243741318e-03*Ip3
ISRC32_p4 0 V32  ac 2.348331413681459e-02*Ip4

ISRC33_p1 0 V33  ac 1.933675915148123e-03*Ip1
ISRC33_p2 0 V33  ac 6.213927148997303e-03*Ip2
ISRC33_p3 0 V33  ac 1.322501588744237e-02*Ip3
ISRC33_p4 0 V33  ac 3.577113763644577e-03*Ip4

ISRC34_p1 0 V34  ac -1.048176760179002e-03*Ip1
ISRC34_p2 0 V34  ac 1.431852336231152e-03*Ip2
ISRC34_p3 0 V34  ac -1.283895086078936e-03*Ip3
ISRC34_p4 0 V34  ac 1.578474511797673e-03*Ip4

ISRC35_p1 0 V35  ac 1.407045960348299e-03*Ip1
ISRC35_p2 0 V35  ac -1.595324180473933e-03*Ip2
ISRC35_p3 0 V35  ac -8.559691582698443e-03*Ip3
ISRC35_p4 0 V35  ac 7.737644877577284e-03*Ip4

ISRC36_p1 0 V36  ac 2.213842092088088e-03*Ip1
ISRC36_p2 0 V36  ac 1.606003230246826e-03*Ip2
ISRC36_p3 0 V36  ac 1.569050493253182e-03*Ip3
ISRC36_p4 0 V36  ac 8.763609005594966e-03*Ip4

ISRC37_p1 0 V37  ac 1.049735546790006e-02*Ip1
ISRC37_p2 0 V37  ac -6.684194164581400e-04*Ip2
ISRC37_p3 0 V37  ac -6.666551338619187e-04*Ip3
ISRC37_p4 0 V37  ac 5.956226445335781e-04*Ip4

ISRC38_p1 0 V38  ac -1.407187331990688e-03*Ip1
ISRC38_p2 0 V38  ac 1.017156832346207e-02*Ip2
ISRC38_p3 0 V38  ac 2.174902055324819e-03*Ip3
ISRC38_p4 0 V38  ac 2.808641197125347e-03*Ip4

ISRC39_p1 0 V39  ac -1.086698066173301e-03*Ip1
ISRC39_p2 0 V39  ac 1.458717068540285e-03*Ip2
ISRC39_p3 0 V39  ac 8.302430987138471e-03*Ip3
ISRC39_p4 0 V39  ac 1.906204914203072e-03*Ip4

ISRC40_p1 0 V40  ac -4.575409546930745e-05*Ip1
ISRC40_p2 0 V40  ac -3.322594930673124e-03*Ip2
ISRC40_p3 0 V40  ac -1.568653435679795e-03*Ip3
ISRC40_p4 0 V40  ac 1.520637019225258e-03*Ip4

ISRC41_p1 0 V41  ac 6.324641924772928e-03*Ip1
ISRC41_p2 0 V41  ac -5.018707518794296e-03*Ip2
ISRC41_p3 0 V41  ac -4.279988000371204e-03*Ip3
ISRC41_p4 0 V41  ac -4.261928790591415e-03*Ip4

ISRC42_p1 0 V42  ac -6.246191288598855e-03*Ip1
ISRC42_p2 0 V42  ac 5.266795785155909e-03*Ip2
ISRC42_p3 0 V42  ac -5.989920215850017e-03*Ip3
ISRC42_p4 0 V42  ac -7.449632076858133e-03*Ip4

ISRC43_p1 0 V43  ac -1.997013831285873e-03*Ip1
ISRC43_p2 0 V43  ac -9.440409333119034e-03*Ip2
ISRC43_p3 0 V43  ac 7.839142411458675e-03*Ip3
ISRC43_p4 0 V43  ac 1.399815942723882e-03*Ip4

ISRC44_p1 0 V44  ac -2.660668310471603e-03*Ip1
ISRC44_p2 0 V44  ac -2.485570012589662e-03*Ip2
ISRC44_p3 0 V44  ac -6.418514288677280e-03*Ip3
ISRC44_p4 0 V44  ac 1.550788141624861e-02*Ip4

ISRC45_p1 0 V45  ac -2.274064214225990e-03*Ip1
ISRC45_p2 0 V45  ac -1.529519659587875e-03*Ip2
ISRC45_p3 0 V45  ac -7.511078268440212e-03*Ip3
ISRC45_p4 0 V45  ac -8.986034273292968e-03*Ip4

ISRC46_p1 0 V46  ac -4.831231851979878e-03*Ip1
ISRC46_p2 0 V46  ac 1.068992628321842e-03*Ip2
ISRC46_p3 0 V46  ac 1.076209894896850e-02*Ip3
ISRC46_p4 0 V46  ac -1.195627505148670e-02*Ip4

ISRC47_p1 0 V47  ac 1.353795420265234e-03*Ip1
ISRC47_p2 0 V47  ac -8.391454213601228e-03*Ip2
ISRC47_p3 0 V47  ac 7.447136263212467e-03*Ip3
ISRC47_p4 0 V47  ac 3.464497216989849e-03*Ip4

ISRC48_p1 0 V48  ac 9.758245927584296e-05*Ip1
ISRC48_p2 0 V48  ac -2.665250710830668e-03*Ip2
ISRC48_p3 0 V48  ac -3.329999207423905e-03*Ip3
ISRC48_p4 0 V48  ac -9.717784983339334e-03*Ip4

ISRC49_p1 0 V49  ac -8.076577271225152e-04*Ip1
ISRC49_p2 0 V49  ac -5.764631343569090e-04*Ip2
ISRC49_p3 0 V49  ac -8.163374450410599e-03*Ip3
ISRC49_p4 0 V49  ac 9.039798430344257e-03*Ip4

ISRC50_p1 0 V50  ac -1.128552230531831e-04*Ip1
ISRC50_p2 0 V50  ac -5.204655384638101e-03*Ip2
ISRC50_p3 0 V50  ac -5.235537915862471e-03*Ip3
ISRC50_p4 0 V50  ac -1.358848809140783e-02*Ip4

ISRC51_p1 0 V51  ac -1.315011857976928e-03*Ip1
ISRC51_p2 0 V51  ac 5.278526471016343e-04*Ip2
ISRC51_p3 0 V51  ac -2.027850101857681e-03*Ip3
ISRC51_p4 0 V51  ac 5.719325882244172e-03*Ip4

ISRC52_p1 0 V52  ac -1.270328470110405e-03*Ip1
ISRC52_p2 0 V52  ac -1.668444353359911e-03*Ip2
ISRC52_p3 0 V52  ac 3.917974122099733e-04*Ip3
ISRC52_p4 0 V52  ac -1.369110652939482e-02*Ip4

ISRC53_p1 0 V53  ac -7.530666599068639e-03*Ip1
ISRC53_p2 0 V53  ac -3.055299715578457e-03*Ip2
ISRC53_p3 0 V53  ac 4.033625208729985e-03*Ip3
ISRC53_p4 0 V53  ac -4.947839613922373e-03*Ip4

ISRC54_p1 0 V54  ac 5.376721403715146e-03*Ip1
ISRC54_p2 0 V54  ac 1.620826710117128e-03*Ip2
ISRC54_p3 0 V54  ac 9.343135626067161e-03*Ip3
ISRC54_p4 0 V54  ac -1.040391298753681e-03*Ip4

ISRC55_p1 0 V55  ac 2.491039181786035e-03*Ip1
ISRC55_p2 0 V55  ac -4.316661069262689e-03*Ip2
ISRC55_p3 0 V55  ac -1.499671619417231e-02*Ip3
ISRC55_p4 0 V55  ac -1.361174485294494e-02*Ip4

ISRC56_p1 0 V56  ac 1.909968355130813e-03*Ip1
ISRC56_p2 0 V56  ac -1.749303580679016e-03*Ip2
ISRC56_p3 0 V56  ac 1.369915262245224e-03*Ip3
ISRC56_p4 0 V56  ac -2.565564116276514e-03*Ip4

ISRC57_p1 0 V57  ac 1.267165599960369e-02*Ip1
ISRC57_p2 0 V57  ac 2.863179139218962e-03*Ip2
ISRC57_p3 0 V57  ac 2.956538476922818e-03*Ip3
ISRC57_p4 0 V57  ac 7.516989781621669e-03*Ip4

ISRC58_p1 0 V58  ac 4.879750948880766e-04*Ip1
ISRC58_p2 0 V58  ac 5.434376864277056e-03*Ip2
ISRC58_p3 0 V58  ac 6.326027445618964e-03*Ip3
ISRC58_p4 0 V58  ac 9.047100428825840e-03*Ip4

ISRC59_p1 0 V59  ac -1.072272065520433e-03*Ip1
ISRC59_p2 0 V59  ac -1.674109743332485e-04*Ip2
ISRC59_p3 0 V59  ac 5.204095602148031e-03*Ip3
ISRC59_p4 0 V59  ac 3.427957297828252e-03*Ip4

ISRC60_p1 0 V60  ac -6.716065409500528e-04*Ip1
ISRC60_p2 0 V60  ac -1.779350410697259e-03*Ip2
ISRC60_p3 0 V60  ac -4.209472988692553e-03*Ip3
ISRC60_p4 0 V60  ac 1.111718799325368e-02*Ip4

ISRC61_p1 0 V61  ac -5.825948799868762e-03*Ip1
ISRC61_p2 0 V61  ac 2.112194593676166e-03*Ip2
ISRC61_p3 0 V61  ac -3.009337004920750e-03*Ip3
ISRC61_p4 0 V61  ac -1.693749273536392e-03*Ip4

ISRC62_p1 0 V62  ac -3.388113340993143e-03*Ip1
ISRC62_p2 0 V62  ac -9.002188224471942e-03*Ip2
ISRC62_p3 0 V62  ac 2.985088321153592e-03*Ip3
ISRC62_p4 0 V62  ac 4.933649645693559e-03*Ip4

ISRC63_p1 0 V63  ac -5.528437715447159e-03*Ip1
ISRC63_p2 0 V63  ac 2.424062360065161e-03*Ip2
ISRC63_p3 0 V63  ac 6.088251466377038e-03*Ip3
ISRC63_p4 0 V63  ac 1.291066981532625e-04*Ip4

ISRC64_p1 0 V64  ac 9.530266858520662e-04*Ip1
ISRC64_p2 0 V64  ac 2.023225406454935e-03*Ip2
ISRC64_p3 0 V64  ac 7.281619181966106e-04*Ip3
ISRC64_p4 0 V64  ac 2.607469687436367e-02*Ip4

ISRC65_p1 0 V65  ac 1.586359905596358e-02*Ip1
ISRC65_p2 0 V65  ac -2.570159214966885e-03*Ip2
ISRC65_p3 0 V65  ac -7.123292363159313e-03*Ip3
ISRC65_p4 0 V65  ac 9.184094888432942e-05*Ip4

ISRC66_p1 0 V66  ac 1.279222278183897e-02*Ip1
ISRC66_p2 0 V66  ac 8.723201597053306e-03*Ip2
ISRC66_p3 0 V66  ac 1.153805676514909e-02*Ip3
ISRC66_p4 0 V66  ac 1.536401842911712e-02*Ip4

ISRC67_p1 0 V67  ac 1.192241650967459e-02*Ip1
ISRC67_p2 0 V67  ac -7.360936810427599e-03*Ip2
ISRC67_p3 0 V67  ac 3.656030147013498e-03*Ip3
ISRC67_p4 0 V67  ac 5.059658455592233e-03*Ip4

ISRC68_p1 0 V68  ac -4.511442623065477e-03*Ip1
ISRC68_p2 0 V68  ac -5.814369453342782e-03*Ip2
ISRC68_p3 0 V68  ac 6.199450113101962e-04*Ip3
ISRC68_p4 0 V68  ac -1.798135874101468e-02*Ip4

ISRC69_p1 0 V69  ac 3.900860179727549e-03*Ip1
ISRC69_p2 0 V69  ac -3.800193364471405e-03*Ip2
ISRC69_p3 0 V69  ac 2.899805701214004e-03*Ip3
ISRC69_p4 0 V69  ac 7.444821376327288e-03*Ip4

ISRC70_p1 0 V70  ac -1.797871005490095e-02*Ip1
ISRC70_p2 0 V70  ac -8.335319047511803e-03*Ip2
ISRC70_p3 0 V70  ac -4.801712039753787e-04*Ip3
ISRC70_p4 0 V70  ac 5.130378253366752e-03*Ip4

ISRC71_p1 0 V71  ac -4.626569659350281e-03*Ip1
ISRC71_p2 0 V71  ac 1.950763489265903e-02*Ip2
ISRC71_p3 0 V71  ac -1.639103045355010e-03*Ip3
ISRC71_p4 0 V71  ac 1.356853863647158e-03*Ip4

ISRC72_p1 0 V72  ac -4.746399639988754e-03*Ip1
ISRC72_p2 0 V72  ac -7.871698811405163e-03*Ip2
ISRC72_p3 0 V72  ac 1.179894188166736e-02*Ip3
ISRC72_p4 0 V72  ac 6.554767157681684e-03*Ip4

ISRC73_p1 0 V73  ac -1.408726436224106e-04*Ip1
ISRC73_p2 0 V73  ac 4.006127159807733e-04*Ip2
ISRC73_p3 0 V73  ac -2.698972795326769e-03*Ip3
ISRC73_p4 0 V73  ac 4.359947535059886e-03*Ip4

ISRC74_p1 0 V74  ac 9.974354191985863e-05*Ip1
ISRC74_p2 0 V74  ac 1.934499587146157e-03*Ip2
ISRC74_p3 0 V74  ac -4.444936747573328e-03*Ip3
ISRC74_p4 0 V74  ac 3.196632094906631e-05*Ip4

ISRC75_p1 0 V75  ac 8.086069110414667e-03*Ip1
ISRC75_p2 0 V75  ac 2.861150925797630e-03*Ip2
ISRC75_p3 0 V75  ac -1.020147482530409e-03*Ip3
ISRC75_p4 0 V75  ac 2.460260362016569e-03*Ip4

ISRC76_p1 0 V76  ac -3.136370674058806e-03*Ip1
ISRC76_p2 0 V76  ac 2.140303011436383e-03*Ip2
ISRC76_p3 0 V76  ac 1.642461471757356e-03*Ip3
ISRC76_p4 0 V76  ac -2.811105470664783e-03*Ip4

ISRC77_p1 0 V77  ac -3.102114090849042e-03*Ip1
ISRC77_p2 0 V77  ac 4.539706886892221e-03*Ip2
ISRC77_p3 0 V77  ac -3.266611386607619e-03*Ip3
ISRC77_p4 0 V77  ac -1.682340536022993e-03*Ip4

ISRC78_p1 0 V78  ac -5.500309188008278e-03*Ip1
ISRC78_p2 0 V78  ac 3.645251361754489e-04*Ip2
ISRC78_p3 0 V78  ac -1.513610731400753e-03*Ip3
ISRC78_p4 0 V78  ac -5.174996872876207e-03*Ip4

ISRC79_p1 0 V79  ac -6.472521663605781e-04*Ip1
ISRC79_p2 0 V79  ac -1.544067143958829e-03*Ip2
ISRC79_p3 0 V79  ac -3.243614101814482e-03*Ip3
ISRC79_p4 0 V79  ac -1.166217408242488e-03*Ip4

ISRC80_p1 0 V80  ac 5.242723270134053e-04*Ip1
ISRC80_p2 0 V80  ac 8.250365682500233e-03*Ip2
ISRC80_p3 0 V80  ac 8.438696892001256e-04*Ip3
ISRC80_p4 0 V80  ac 2.898555832567650e-03*Ip4

ISRC81_p1 0 V81  ac -9.050064902309427e-04*Ip1
ISRC81_p2 0 V81  ac 1.114015962956693e-03*Ip2
ISRC81_p3 0 V81  ac 2.058949452453598e-03*Ip3
ISRC81_p4 0 V81  ac 7.970752844730157e-03*Ip4

ISRC82_p1 0 V82  ac -1.778325163484467e-03*Ip1
ISRC82_p2 0 V82  ac 2.470867096029108e-03*Ip2
ISRC82_p3 0 V82  ac -4.554674378273517e-03*Ip3
ISRC82_p4 0 V82  ac 3.365988117595225e-04*Ip4

ISRC83_p1 0 V83  ac -1.172110526177762e-03*Ip1
ISRC83_p2 0 V83  ac 4.512782485409501e-03*Ip2
ISRC83_p3 0 V83  ac 6.556299890350756e-06*Ip3
ISRC83_p4 0 V83  ac -6.382949921531413e-04*Ip4

ISRC84_p1 0 V84  ac 6.965333394744981e-04*Ip1
ISRC84_p2 0 V84  ac 6.029265519806254e-03*Ip2
ISRC84_p3 0 V84  ac 7.085823103334453e-03*Ip3
ISRC84_p4 0 V84  ac -1.653321673452158e-03*Ip4

ISRC85_p1 0 V85  ac -7.393430351475031e-03*Ip1
ISRC85_p2 0 V85  ac 2.770745612920664e-04*Ip2
ISRC85_p3 0 V85  ac 3.827911694640923e-03*Ip3
ISRC85_p4 0 V85  ac 7.043190364653214e-03*Ip4

ISRC86_p1 0 V86  ac -4.834600325943211e-03*Ip1
ISRC86_p2 0 V86  ac -7.210929999218544e-03*Ip2
ISRC86_p3 0 V86  ac -2.570369090992396e-03*Ip3
ISRC86_p4 0 V86  ac 1.596799643522864e-02*Ip4

ISRC87_p1 0 V87  ac 1.639274895166965e-03*Ip1
ISRC87_p2 0 V87  ac 1.694630917696926e-03*Ip2
ISRC87_p3 0 V87  ac -8.214019213997038e-03*Ip3
ISRC87_p4 0 V87  ac -3.643206295791067e-03*Ip4

ISRC88_p1 0 V88  ac 1.273668665799432e-04*Ip1
ISRC88_p2 0 V88  ac -3.817852173249642e-03*Ip2
ISRC88_p3 0 V88  ac -1.954991135919028e-03*Ip3
ISRC88_p4 0 V88  ac -6.506700252870971e-03*Ip4

ISRC89_p1 0 V89  ac 7.295067025886404e-03*Ip1
ISRC89_p2 0 V89  ac 1.963231430110190e-04*Ip2
ISRC89_p3 0 V89  ac 1.784236587433312e-03*Ip3
ISRC89_p4 0 V89  ac -1.121889924195504e-03*Ip4

ISRC90_p1 0 V90  ac -1.171810664883530e-03*Ip1
ISRC90_p2 0 V90  ac 4.486712646037810e-04*Ip2
ISRC90_p3 0 V90  ac -3.861963264175038e-03*Ip3
ISRC90_p4 0 V90  ac 2.851688308081966e-03*Ip4

ISRC91_p1 0 V91  ac -3.118924159780281e-03*Ip1
ISRC91_p2 0 V91  ac -2.600545537240776e-03*Ip2
ISRC91_p3 0 V91  ac 4.727380822120719e-03*Ip3
ISRC91_p4 0 V91  ac -1.240026442435307e-03*Ip4

ISRC92_p1 0 V92  ac 3.148192348582590e-04*Ip1
ISRC92_p2 0 V92  ac 9.430618816540735e-04*Ip2
ISRC92_p3 0 V92  ac -5.245285164035843e-03*Ip3
ISRC92_p4 0 V92  ac 5.533049966170791e-03*Ip4

ISRC93_p1 0 V93  ac -2.117927387980365e-02*Ip1
ISRC93_p2 0 V93  ac 3.423908258029789e-03*Ip2
ISRC93_p3 0 V93  ac 2.152142944967626e-03*Ip3
ISRC93_p4 0 V93  ac 2.517612886030656e-03*Ip4

ISRC94_p1 0 V94  ac -7.384616881916622e-03*Ip1
ISRC94_p2 0 V94  ac 1.209120992174927e-03*Ip2
ISRC94_p3 0 V94  ac -1.411047309813515e-03*Ip3
ISRC94_p4 0 V94  ac -3.410800762288906e-03*Ip4

ISRC95_p1 0 V95  ac -1.477493842825339e-03*Ip1
ISRC95_p2 0 V95  ac 7.953774915104673e-03*Ip2
ISRC95_p3 0 V95  ac 3.120819196924550e-03*Ip3
ISRC95_p4 0 V95  ac 7.884847209801468e-04*Ip4

ISRC96_p1 0 V96  ac 3.852033154375753e-03*Ip1
ISRC96_p2 0 V96  ac 9.212838139054983e-04*Ip2
ISRC96_p3 0 V96  ac 1.475260001194145e-02*Ip3
ISRC96_p4 0 V96  ac 7.450697559579278e-04*Ip4

ISRC97_p1 0 V97  ac -1.104443728978292e-02*Ip1
ISRC97_p2 0 V97  ac -7.986175864918047e-03*Ip2
ISRC97_p3 0 V97  ac 6.061719858711083e-03*Ip3
ISRC97_p4 0 V97  ac 8.678418880698013e-04*Ip4

ISRC98_p1 0 V98  ac -1.332324413921675e-02*Ip1
ISRC98_p2 0 V98  ac 2.672154906104989e-03*Ip2
ISRC98_p3 0 V98  ac 5.835491044417039e-04*Ip3
ISRC98_p4 0 V98  ac -4.071227463307991e-03*Ip4

ISRC99_p1 0 V99  ac -6.852119081119081e-03*Ip1
ISRC99_p2 0 V99  ac 5.356838571212312e-03*Ip2
ISRC99_p3 0 V99  ac -4.427421031621993e-03*Ip3
ISRC99_p4 0 V99  ac -2.354408832712312e-03*Ip4

ISRC100_p1 0 V100  ac 3.666903188651501e-03*Ip1
ISRC100_p2 0 V100  ac 7.044406275531569e-05*Ip2
ISRC100_p3 0 V100  ac 8.267127980598140e-03*Ip3
ISRC100_p4 0 V100  ac -1.242565560792767e-02*Ip4

ISRC101_p1 0 V101  ac -7.895838174250399e-03*Ip1
ISRC101_p2 0 V101  ac -3.852769943010937e-03*Ip2
ISRC101_p3 0 V101  ac 1.175749956429380e-03*Ip3
ISRC101_p4 0 V101  ac -6.833666388873662e-04*Ip4

ISRC102_p1 0 V102  ac -5.001905720831757e-03*Ip1
ISRC102_p2 0 V102  ac 7.615789786343760e-03*Ip2
ISRC102_p3 0 V102  ac -1.518808320272783e-02*Ip3
ISRC102_p4 0 V102  ac -9.738473735011934e-03*Ip4

ISRC103_p1 0 V103  ac -1.710401773318942e-03*Ip1
ISRC103_p2 0 V103  ac -9.809158988214937e-03*Ip2
ISRC103_p3 0 V103  ac -4.426456889558856e-03*Ip3
ISRC103_p4 0 V103  ac -2.695475704600838e-03*Ip4

ISRC104_p1 0 V104  ac -2.736565633752142e-05*Ip1
ISRC104_p2 0 V104  ac 2.297595757455079e-03*Ip2
ISRC104_p3 0 V104  ac 1.191655171400520e-03*Ip3
ISRC104_p4 0 V104  ac 1.225256452920634e-02*Ip4

ISRC105_p1 0 V105  ac 9.594756020429963e-03*Ip1
ISRC105_p2 0 V105  ac 9.954000521859276e-03*Ip2
ISRC105_p3 0 V105  ac 7.295712150569758e-03*Ip3
ISRC105_p4 0 V105  ac -7.900830096723783e-03*Ip4

ISRC106_p1 0 V106  ac 9.327564779386855e-03*Ip1
ISRC106_p2 0 V106  ac -3.453431865016474e-04*Ip2
ISRC106_p3 0 V106  ac 6.148653551475385e-03*Ip3
ISRC106_p4 0 V106  ac 5.477183912819458e-03*Ip4

ISRC107_p1 0 V107  ac -3.532827724538975e-03*Ip1
ISRC107_p2 0 V107  ac -3.061948690011276e-05*Ip2
ISRC107_p3 0 V107  ac 3.691864214329156e-03*Ip3
ISRC107_p4 0 V107  ac -1.645884629806138e-03*Ip4

ISRC108_p1 0 V108  ac -1.972563144291352e-03*Ip1
ISRC108_p2 0 V108  ac 1.391946112819302e-02*Ip2
ISRC108_p3 0 V108  ac 1.166103711750789e-02*Ip3
ISRC108_p4 0 V108  ac -7.075753672756239e-03*Ip4

ISRC109_p1 0 V109  ac -4.752489178355556e-03*Ip1
ISRC109_p2 0 V109  ac -1.086165417537380e-04*Ip2
ISRC109_p3 0 V109  ac -3.966212958258216e-03*Ip3
ISRC109_p4 0 V109  ac 2.532796503968637e-02*Ip4

ISRC110_p1 0 V110  ac 1.381227677641326e-03*Ip1
ISRC110_p2 0 V110  ac 8.077587103289785e-03*Ip2
ISRC110_p3 0 V110  ac -1.227346242536562e-02*Ip3
ISRC110_p4 0 V110  ac -4.621666790731322e-04*Ip4

ISRC111_p1 0 V111  ac 5.011832926578092e-03*Ip1
ISRC111_p2 0 V111  ac -7.356623493012281e-03*Ip2
ISRC111_p3 0 V111  ac -3.352720715299541e-04*Ip3
ISRC111_p4 0 V111  ac -2.282596986742242e-03*Ip4

ISRC112_p1 0 V112  ac 2.179718812752370e-03*Ip1
ISRC112_p2 0 V112  ac 7.606796928063222e-03*Ip2
ISRC112_p3 0 V112  ac -7.709575355168167e-03*Ip3
ISRC112_p4 0 V112  ac 5.527361791952841e-04*Ip4

ISRC113_p1 0 V113  ac 6.000195415157086e-03*Ip1
ISRC113_p2 0 V113  ac 7.263097860189795e-03*Ip2
ISRC113_p3 0 V113  ac 7.045016326804056e-03*Ip3
ISRC113_p4 0 V113  ac -1.536334166531749e-02*Ip4

ISRC114_p1 0 V114  ac -3.448043120003624e-03*Ip1
ISRC114_p2 0 V114  ac -1.654565471452592e-03*Ip2
ISRC114_p3 0 V114  ac 1.311781455502847e-02*Ip3
ISRC114_p4 0 V114  ac 1.580752913073906e-03*Ip4

ISRC115_p1 0 V115  ac -7.432600717936885e-03*Ip1
ISRC115_p2 0 V115  ac 1.466905698991494e-02*Ip2
ISRC115_p3 0 V115  ac -5.447079733475513e-03*Ip3
ISRC115_p4 0 V115  ac 2.907222902259507e-03*Ip4

ISRC116_p1 0 V116  ac -3.294207437120392e-03*Ip1
ISRC116_p2 0 V116  ac 9.296744007862516e-04*Ip2
ISRC116_p3 0 V116  ac 1.316697979649944e-02*Ip3
ISRC116_p4 0 V116  ac 1.511981669632378e-03*Ip4

ISRC117_p1 0 V117  ac -1.008277186238438e-02*Ip1
ISRC117_p2 0 V117  ac -4.159504540313699e-03*Ip2
ISRC117_p3 0 V117  ac 4.039902850680092e-03*Ip3
ISRC117_p4 0 V117  ac 1.053931955759978e-02*Ip4

ISRC118_p1 0 V118  ac 8.310808966793641e-03*Ip1
ISRC118_p2 0 V118  ac 3.695848789909233e-03*Ip2
ISRC118_p3 0 V118  ac -8.045187819829687e-03*Ip3
ISRC118_p4 0 V118  ac 6.212341211878387e-03*Ip4

ISRC119_p1 0 V119  ac 1.157396164389935e-02*Ip1
ISRC119_p2 0 V119  ac 7.793864030888750e-04*Ip2
ISRC119_p3 0 V119  ac -2.806493126208042e-03*Ip3
ISRC119_p4 0 V119  ac -5.478757891465721e-03*Ip4

ISRC120_p1 0 V120  ac -9.399928098590317e-03*Ip1
ISRC120_p2 0 V120  ac -9.383156819497140e-04*Ip2
ISRC120_p3 0 V120  ac -2.841289584824904e-03*Ip3
ISRC120_p4 0 V120  ac -9.644297751592333e-03*Ip4

ISRC121_p1 0 V121  ac 6.973266424962036e-03*Ip1
ISRC121_p2 0 V121  ac 4.679605569630897e-04*Ip2
ISRC121_p3 0 V121  ac -5.926367081411161e-03*Ip3
ISRC121_p4 0 V121  ac 2.056489921289263e-03*Ip4

ISRC122_p1 0 V122  ac 7.444069759469345e-03*Ip1
ISRC122_p2 0 V122  ac 1.152901498832748e-02*Ip2
ISRC122_p3 0 V122  ac 1.703951198537643e-03*Ip3
ISRC122_p4 0 V122  ac 2.722183135326872e-03*Ip4

ISRC123_p1 0 V123  ac -2.898803656346932e-03*Ip1
ISRC123_p2 0 V123  ac -3.403439820304659e-03*Ip2
ISRC123_p3 0 V123  ac 7.825764068833046e-04*Ip3
ISRC123_p4 0 V123  ac 1.944545263147081e-04*Ip4

ISRC124_p1 0 V124  ac 1.169489822020017e-03*Ip1
ISRC124_p2 0 V124  ac 1.452536770039820e-03*Ip2
ISRC124_p3 0 V124  ac -5.943937938148350e-03*Ip3
ISRC124_p4 0 V124  ac -1.438558693809106e-02*Ip4

ISRC125_p1 0 V125  ac -1.574430361350370e-02*Ip1
ISRC125_p2 0 V125  ac 3.299343445670577e-03*Ip2
ISRC125_p3 0 V125  ac 1.008817029506263e-03*Ip3
ISRC125_p4 0 V125  ac 5.853942663290103e-03*Ip4

ISRC126_p1 0 V126  ac -6.563412516697788e-03*Ip1
ISRC126_p2 0 V126  ac -6.114543639451758e-03*Ip2
ISRC126_p3 0 V126  ac 3.838454254361517e-03*Ip3
ISRC126_p4 0 V126  ac -2.640542271695792e-03*Ip4

ISRC127_p1 0 V127  ac -2.500214855138326e-03*Ip1
ISRC127_p2 0 V127  ac 5.147229561216031e-03*Ip2
ISRC127_p3 0 V127  ac -6.264375015465108e-03*Ip3
ISRC127_p4 0 V127  ac -8.584530063463330e-03*Ip4

ISRC128_p1 0 V128  ac -3.904808242866301e-03*Ip1
ISRC128_p2 0 V128  ac -1.386802758053344e-03*Ip2
ISRC128_p3 0 V128  ac -4.936300131828784e-03*Ip3
ISRC128_p4 0 V128  ac -2.831809547365511e-03*Ip4

ISRC129_p1 0 V129  ac -5.117233089399107e-03*Ip1
ISRC129_p2 0 V129  ac 1.526894796730689e-03*Ip2
ISRC129_p3 0 V129  ac -7.289986851222383e-03*Ip3
ISRC129_p4 0 V129  ac -6.330807820952292e-03*Ip4

ISRC130_p1 0 V130  ac -2.364870696619276e-03*Ip1
ISRC130_p2 0 V130  ac 3.397663456203753e-03*Ip2
ISRC130_p3 0 V130  ac -1.026918446806047e-02*Ip3
ISRC130_p4 0 V130  ac -6.246209810759353e-04*Ip4

ISRC131_p1 0 V131  ac -3.614831628136720e-03*Ip1
ISRC131_p2 0 V131  ac 5.122497425628946e-04*Ip2
ISRC131_p3 0 V131  ac -3.862787805881542e-03*Ip3
ISRC131_p4 0 V131  ac 2.122636736412996e-03*Ip4

ISRC132_p1 0 V132  ac 8.781075936361223e-04*Ip1
ISRC132_p2 0 V132  ac -2.113162567853712e-03*Ip2
ISRC132_p3 0 V132  ac 3.196561090854507e-04*Ip3
ISRC132_p4 0 V132  ac 3.650977316633442e-03*Ip4

ISRC133_p1 0 V133  ac 3.240692405894743e-03*Ip1
ISRC133_p2 0 V133  ac -1.320649694302663e-03*Ip2
ISRC133_p3 0 V133  ac 3.764902031656979e-03*Ip3
ISRC133_p4 0 V133  ac -1.022047218521783e-03*Ip4

ISRC134_p1 0 V134  ac 1.299557373257865e-02*Ip1
ISRC134_p2 0 V134  ac -1.199699215588814e-04*Ip2
ISRC134_p3 0 V134  ac -1.102118172567805e-02*Ip3
ISRC134_p4 0 V134  ac -6.582343919146034e-04*Ip4

ISRC135_p1 0 V135  ac 2.710016143834529e-03*Ip1
ISRC135_p2 0 V135  ac -2.784756927489527e-03*Ip2
ISRC135_p3 0 V135  ac 2.094128490592779e-03*Ip3
ISRC135_p4 0 V135  ac -4.350827751155229e-03*Ip4

ISRC136_p1 0 V136  ac -2.235374724720000e-03*Ip1
ISRC136_p2 0 V136  ac -4.085805514367681e-04*Ip2
ISRC136_p3 0 V136  ac -4.221852679971540e-04*Ip3
ISRC136_p4 0 V136  ac -2.693932168828197e-03*Ip4

ISRC137_p1 0 V137  ac -1.161446328698614e-02*Ip1
ISRC137_p2 0 V137  ac 1.766365790343214e-03*Ip2
ISRC137_p3 0 V137  ac -9.459391300391772e-03*Ip3
ISRC137_p4 0 V137  ac -1.367544566960272e-02*Ip4

ISRC138_p1 0 V138  ac 3.312210690588179e-04*Ip1
ISRC138_p2 0 V138  ac -1.246698840889468e-02*Ip2
ISRC138_p3 0 V138  ac -5.669675579892195e-03*Ip3
ISRC138_p4 0 V138  ac -1.247503591727212e-02*Ip4

ISRC139_p1 0 V139  ac -1.312627831663283e-02*Ip1
ISRC139_p2 0 V139  ac 1.223651590186538e-02*Ip2
ISRC139_p3 0 V139  ac 4.111108649677790e-03*Ip3
ISRC139_p4 0 V139  ac 3.825224023842333e-03*Ip4

ISRC140_p1 0 V140  ac 7.547943818020987e-03*Ip1
ISRC140_p2 0 V140  ac 7.967225905283763e-03*Ip2
ISRC140_p3 0 V140  ac 5.219962793316524e-03*Ip3
ISRC140_p4 0 V140  ac 6.817620454113468e-03*Ip4

ISRC141_p1 0 V141  ac -5.588090231627570e-03*Ip1
ISRC141_p2 0 V141  ac -2.595346674111618e-03*Ip2
ISRC141_p3 0 V141  ac -4.805606464368197e-03*Ip3
ISRC141_p4 0 V141  ac 5.119140217969091e-04*Ip4

ISRC142_p1 0 V142  ac 1.006705391060052e-02*Ip1
ISRC142_p2 0 V142  ac 6.922426863419029e-03*Ip2
ISRC142_p3 0 V142  ac 1.440748176176290e-02*Ip3
ISRC142_p4 0 V142  ac -4.520554812414901e-03*Ip4

ISRC143_p1 0 V143  ac 2.086322751841429e-03*Ip1
ISRC143_p2 0 V143  ac 9.738112370383054e-04*Ip2
ISRC143_p3 0 V143  ac 8.710365012514094e-04*Ip3
ISRC143_p4 0 V143  ac -4.724276813945843e-03*Ip4

ISRC144_p1 0 V144  ac 1.114021717758165e-02*Ip1
ISRC144_p2 0 V144  ac -9.764262503083364e-03*Ip2
ISRC144_p3 0 V144  ac 4.616438761935150e-03*Ip3
ISRC144_p4 0 V144  ac -1.312957291002842e-02*Ip4


.ends subckt equivalent_circuit

.end

