* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 node_ref
X_11 node_1 node_ref yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 node_ref yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 node_ref yp33
X_34 node_3 node_4 yp34
X_44 node_4 node_ref yp44
.ends


* Y'11
.subckt yp11 node_1 node_ref
* Branch 0
Rabr0 node_1 netRa0 465.3590496994122
Lbr0 netRa0 netL0 1.0535927569713485e-12
Rbbr0 netL0 node_ref 3419.170790757784
Cbr0 netL0 node_ref 6.802531243650122e-19

* Branch 1
Rabr1 node_1 netRa1 78.14116472376968
Lbr1 netRa1 netL1  1.3219148027074502e-13
Rbbr1 netL1 node_ref 333.6040827306789
Cbr1 netL1 node_ref  4.657809257395912e-18

* Branch 2
Rabr2 node_1 netRa2  18053.815557757902
Lbr2 netRa2 netL2 6.515442612087674e-11
Rbbr2 netL2 node_ref  310385.7429602686
Cbr2 netL2 node_ref 1.156324040106853e-20

* Branch 3
Rabr3 node_1 netRa3  1623.3620446699088
Lbr3 netRa3 netL3 2.36858486398064e-12
Rbbr3 netL3 node_ref  5906.826978499476
Cbr3 netL3 node_ref 2.445840783404925e-19

* Branch 4
Rabr4 node_1 netRa4  19.581655304066693
Lbr4 netRa4 netL4 1.3825295800916076e-13
Rbbr4 netL4 node_ref  1179.8068774603723
Cbr4 netL4 node_ref 5.426132852258792e-18

* Branch 5
Rabr5 node_1 netRa5 630.4506311309683
Lbr5 netRa5 netL5 2.0413388890010182e-12
Rbbr5 netL5 node_ref 9592.721564292142
Cbr5 netL5 node_ref 3.4495963802903313e-19

* Branch 6
Rabr6 node_1 netRa6 221.1898149394218
Lbr6 netRa6 netL6 1.4830156552455697e-12
Rbbr6 netL6 node_ref 14631.97850367413
Cbr6 netL6 node_ref 4.847340063792159e-19

* Branch 7
Rabr7 node_1 netRa7 32642.417619454816
Lbr7 netRa7 netL7 5.111294910101473e-11
Rbbr7 netL7 node_ref 143753.85579243323
Cbr7 netL7 node_ref 1.0916411455822865e-20

* Branch 8
Rabr8 node_1 netRa8 558.4566506955852
Lbr8 netRa8 netL8  3.827956750077595e-13
Rbbr8 netL8 node_ref 918.7678847714785
Cbr8 netL8 node_ref  7.317273900273909e-19

* Branch 9
Rabr9 node_1 netRa9  10990.712259826938
Lbr9 netRa9 netL9 2.5406465712456204e-12
Rbbr9 netL9 node_ref  11820.052020040788
Cbr9 netL9 node_ref 1.9491914723442453e-20

* Branch 10
Rabr10 node_1 netRa10 803890.1083318385
Lbr10 netRa10 netL10  3.4252845431400583e-10
Rbbr10 netL10 node_ref 1015303.1126398303
Cbr10 netL10 node_ref  4.1941428276042376e-22

* Branch 11
Rabr11 node_1 netRa11  788.9155049066959
Lbr11 netRa11 netL11 3.651745155623721e-12
Rbbr11 netL11 node_ref  24826.473706082976
Cbr11 netL11 node_ref 1.824745669782806e-19

* Branch 12
Rabr12 node_1 netRa12 103.38680034091067
Lbr12 netRa12 netL12 2.3150502575375388e-12
Rbbr12 netL12 node_ref 90597.8696169187
Cbr12 netL12 node_ref 2.885063378808514e-19

* Branch 13
Rabr13 node_1 netRa13 12.20824003472247
Lbr13 netRa13 netL13 1.1599667513668128e-13
Rbbr13 netL13 node_ref 1975.6100586608272
Cbr13 netL13 node_ref 5.603642594393949e-18

* Branch 14
Rabr14 node_1 netRa14 842.0831866748524
Lbr14 netRa14 netL14 9.722840537266248e-13
Rbbr14 netL14 node_ref 2641.74279288616
Cbr14 netL14 node_ref 4.429147642408437e-19

* Branch 15
Rabr15 node_1 netRa15  8.26267721579585
Lbr15 netRa15 netL15  1.4772371412347928e-14
Rbbr15 netL15 node_ref  102.81567745828492
Cbr15 netL15 node_ref  3.9179281502971683e-17

* Branch 16
Rabr16 node_1 netRa16  274.87284187788606
Lbr16 netRa16 netL16  4.357188101093571e-12
Rbbr16 netL16 node_ref  119388.63481255948
Cbr16 netL16 node_ref  1.4391181131667356e-19

* Branch 17
Rabr17 node_1 netRa17 1124.928715423784
Lbr17 netRa17 netL17 1.0343206962553166e-12
Rbbr17 netL17 node_ref 2684.7069972239133
Cbr17 netL17 node_ref 3.460016386826557e-19

* Branch 18
Rabr18 node_1 netRa18 842.9209060219782
Lbr18 netRa18 netL18  1.0234319651247775e-12
Rbbr18 netL18 node_ref 2845.9080269412034
Cbr18 netL18 node_ref  4.187697351219914e-19

* Branch 19
Rabr19 node_1 netRa19 362936.280741566
Lbr19 netRa19 netL19 1.9852301454367583e-10
Rbbr19 netL19 node_ref 543955.9525525789
Cbr19 netL19 node_ref 1.0060314344016708e-21

* Branch 20
Rabr20 node_1 netRa20  425.1937499250724
Lbr20 netRa20 netL20 5.562519011631224e-12
Rbbr20 netL20 node_ref  116491.71679044554
Cbr20 netL20 node_ref 1.0715663793836882e-19

* Branch 21
Rabr21 node_1 netRa21 1.8225771401012247
Lbr21 netRa21 netL21 2.692225460845098e-12
Rbbr21 netL21 node_ref  1014073.5784445624
Cbr21 netL21 node_ref 2.1639589801258422e-19

* Branch 22
Rabr22 node_1 netRa22  3.263449486113174
Lbr22 netRa22 netL22 1.1532283695219184e-13
Rbbr22 netL22 node_ref  4768.733671935622
Cbr22 netL22 node_ref 4.9138051304811e-18

* Branch 23
Rabr23 node_1 netRa23 98.10504060041033
Lbr23 netRa23 netL23  1.5185133741790936e-13
Rbbr23 netL23 node_ref 474.07252779279884
Cbr23 netL23 node_ref  2.920515512409872e-18

* Branch 24
Rabr24 node_1 netRa24  1038.6043932901548
Lbr24 netRa24 netL24 2.0762566563976822e-12
Rbbr24 netL24 node_ref  8442.816570698466
Cbr24 netL24 node_ref 2.332946229193833e-19

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 565.3184456620916
Lbr0 netRa0 netL0 1.1291878313412533e-12
Rbbr0 netL0 node_2 3349.3207912130088
Cbr0 netL0 node_2 6.107000646126544e-19

* Branch 1
Rabr1 node_1 netRa1  2798.4465923124008
Lbr1 netRa1 netL1  2.2558042332518356e-12
Rbbr1 netL1 node_2  5159.757560713924
Cbr1 netL1 node_2  1.6312147317755216e-19

* Branch 2
Rabr2 node_1 netRa2  1868092.94764946
Lbr2 netRa2 netL2 8.897094488742557e-10
Rbbr2 netL2 node_2  2397429.9962005904
Cbr2 netL2 node_2 1.9851217464340905e-22

* Branch 3
Rabr3 node_1 netRa3 7724707.10493273
Lbr3 netRa3 netL3 5.957333013190807e-10
Rbbr3 netL3 node_2 7782247.59615922
Cbr3 netL3 node_2 9.915002074007648e-24

* Branch 4
Rabr4 node_1 netRa4  17.701654474268363
Lbr4 netRa4 netL4  8.585257349416879e-13
Rbbr4 netL4 node_2  186078.0501984501
Cbr4 netL4 node_2  8.884619670286928e-19

* Branch 5
Rabr5 node_1 netRa5  171611.07697561168
Lbr5 netRa5 netL5 1.1079315104385917e-10
Rbbr5 netL5 node_2  266107.2478980396
Cbr5 netL5 node_2 2.415748708993497e-21

* Branch 6
Rabr6 node_1 netRa6 18849.332278744936
Lbr6 netRa6 netL6  8.993318324713527e-11
Rbbr6 netL6 node_2 584695.0225715635
Cbr6 netL6 node_2  7.854402962089361e-21

* Branch 7
Rabr7 node_1 netRa7 806250.3164874004
Lbr7 netRa7 netL7  1.1316227105521114e-09
Rbbr7 netL7 node_2 3002144.2990635335
Cbr7 netL7 node_2  4.666053567212349e-22

* Branch 8
Rabr8 node_1 netRa8  581052.0099498214
Lbr8 netRa8 netL8 6.452719639206344e-11
Rbbr8 netL8 node_2  591053.1743275005
Cbr8 netL8 node_2 1.8729472772607427e-22

* Branch 9
Rabr9 node_1 netRa9 83.46103487609531
Lbr9 netRa9 netL9 8.792673791781152e-13
Rbbr9 netL9 node_2 15557.155403982748
Cbr9 netL9 node_2 7.984146953490269e-19

* Branch 10
Rabr10 node_1 netRa10 25967705.353225134
Lbr10 netRa10 netL10  4.022631207121687e-09
Rbbr10 netL10 node_2 26870705.97873812
Cbr10 netL10 node_2  5.76371696681098e-24

* Branch 11
Rabr11 node_1 netRa11  115233.97822260883
Lbr11 netRa11 netL11  1.8451864510957146e-10
Rbbr11 netL11 node_2  547802.8696809304
Cbr11 netL11 node_2  2.9452232222876746e-21

* Branch 12
Rabr12 node_1 netRa12 1009847.660903161
Lbr12 netRa12 netL12 3.556861975612034e-10
Rbbr12 netL12 node_2 1197626.4832951382
Cbr12 netL12 node_2 2.947608989048322e-22

* Branch 13
Rabr13 node_1 netRa13 39.118371276354
Lbr13 netRa13 netL13  8.456004641721166e-13
Rbbr13 netL13 node_2 21172.057729432145
Cbr13 netL13 node_2  7.720396997797725e-19

* Branch 14
Rabr14 node_1 netRa14 33683.49459213949
Lbr14 netRa14 netL14 5.852752231925972e-11
Rbbr14 netL14 node_2 197820.337569444
Cbr14 netL14 node_2 8.961660367070948e-21

* Branch 15
Rabr15 node_1 netRa15  65.74546330304061
Lbr15 netRa15 netL15 2.1173652431683889e-13
Rbbr15 netL15 node_2  606.9975738355852
Cbr15 netL15 node_2 2.6503765540801095e-18

* Branch 16
Rabr16 node_1 netRa16 8130060.753178986
Lbr16 netRa16 netL16  1.293992602754745e-09
Rbbr16 netL16 node_2 8457498.420169717
Cbr16 netL16 node_2  1.8804366696168042e-23

* Branch 17
Rabr17 node_1 netRa17  725186.8026396815
Lbr17 netRa17 netL17 1.1060068276134998e-10
Rbbr17 netL17 node_2  752524.7198856114
Cbr17 netL17 node_2 2.023271863040074e-22

* Branch 18
Rabr18 node_1 netRa18 171.58803057562227
Lbr18 netRa18 netL18 7.787714871792324e-13
Rbbr18 netL18 node_2 6413.954274531287
Cbr18 netL18 node_2 7.610099091511814e-19

* Branch 19
Rabr19 node_1 netRa19 10027871.338044755
Lbr19 netRa19 netL19  2.455072402010571e-09
Rbbr19 netL19 node_2 11029190.01843211
Cbr19 netL19 node_2  2.219344736294675e-23

* Branch 20
Rabr20 node_1 netRa20 47801.51185253626
Lbr20 netRa20 netL20  1.1872787323258382e-10
Rbbr20 netL20 node_2 536277.7115515383
Cbr20 netL20 node_2  4.589650662477695e-21

* Branch 21
Rabr21 node_1 netRa21  45921.049905922904
Lbr21 netRa21 netL21 8.788016298335461e-11
Rbbr21 netL21 node_2  331733.92458000267
Cbr21 netL21 node_2 5.711638578521806e-21

* Branch 22
Rabr22 node_1 netRa22  102.64977421684704
Lbr22 netRa22 netL22  8.913120462946025e-13
Rbbr22 netL22 node_2  15697.537857713005
Cbr22 netL22 node_2  6.320500968432652e-19

* Branch 23
Rabr23 node_1 netRa23 52302.512499907956
Lbr23 netRa23 netL23  4.250317183595329e-12
Rbbr23 netL23 node_2 52916.36829383442
Cbr23 netL23 node_2  1.5262568490255976e-21

* Branch 24
Rabr24 node_1 netRa24  1852.9921212517875
Lbr24 netRa24 netL24  2.489342683077404e-11
Rbbr24 netL24 node_2  674891.4273090736
Cbr24 netL24 node_2  2.2126643264632092e-20

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 452.254862529488
Lbr0 netRa0 netL0 9.033503678841172e-13
Rbbr0 netL0 node_3 2679.4567174644963
Cbr0 netL0 node_3 7.633749624420183e-19

* Branch 1
Rabr1 node_1 netRa1  2238.7580853609916
Lbr1 netRa1 netL1  1.8046428072568314e-12
Rbbr1 netL1 node_3  4127.804905468089
Cbr1 netL1 node_3  2.0390175241761034e-19

* Branch 2
Rabr2 node_1 netRa2  1494472.5704617177
Lbr2 netRa2 netL2 7.117668382189893e-10
Rbbr2 netL2 node_3  1917941.8580084923
Cbr2 netL2 node_3 2.4814054050811585e-22

* Branch 3
Rabr3 node_1 netRa3 6179785.527150136
Lbr3 netRa3 netL3 4.765872585842643e-10
Rbbr3 netL3 node_3 6225817.891566737
Cbr3 netL3 node_3 1.2393689397841176e-23

* Branch 4
Rabr4 node_1 netRa4  14.161358288591625
Lbr4 netRa4 netL4  6.868205942288705e-13
Rbbr4 netL4 node_3  148861.20260526586
Cbr4 netL4 node_3  1.1105774475010846e-18

* Branch 5
Rabr5 node_1 netRa5  137288.30020399016
Lbr5 netRa5 netL5 8.863430171660088e-11
Rbbr5 netL5 node_3  212885.17176211547
Cbr5 netL5 node_3 3.019699635263966e-21

* Branch 6
Rabr6 node_1 netRa6 15079.369081858262
Lbr6 netRa6 netL6  7.19465203264736e-11
Rbbr6 netL6 node_3 467758.39225618466
Cbr6 netL6 node_3  9.818011045871765e-21

* Branch 7
Rabr7 node_1 netRa7 645001.5910415638
Lbr7 netRa7 netL7  9.053009430975665e-10
Rbbr7 netL7 node_3 2401723.898284056
Cbr7 netL7 node_3  5.832552183428765e-22

* Branch 8
Rabr8 node_1 netRa8  464843.0535505105
Lbr8 netRa8 netL8 5.1621846013586355e-11
Rbbr8 netL8 node_3  472843.9877634971
Cbr8 netL8 node_3 2.341173687023611e-22

* Branch 9
Rabr9 node_1 netRa9 66.76880494581424
Lbr9 netRa9 netL9 7.03413951775661e-13
Rbbr9 netL9 node_3 12445.73117527794
Cbr9 netL9 node_3 9.980183052826583e-19

* Branch 10
Rabr10 node_1 netRa10 20773421.704153534
Lbr10 netRa10 netL10  3.2180446540102308e-09
Rbbr10 netL10 node_3 21495820.94695395
Cbr10 netL10 node_3  7.205018005353678e-24

* Branch 11
Rabr11 node_1 netRa11  92187.76287732941
Lbr11 netRa11 netL11  1.4761484954439377e-10
Rbbr11 netL11 node_3  438240.36800648115
Cbr11 netL11 node_3  3.681520199783549e-21

* Branch 12
Rabr12 node_1 netRa12 807887.7600959836
Lbr12 netRa12 netL12 2.845504314587136e-10
Rbbr12 netL12 node_3 958110.5805221625
Cbr12 netL12 node_3 3.6844502081088883e-22

* Branch 13
Rabr13 node_1 netRa13 31.294712639161734
Lbr13 netRa13 netL13  6.76480330756411e-13
Rbbr13 netL13 node_3 16937.63803801074
Cbr13 netL13 node_3  9.6504968086634e-19

* Branch 14
Rabr14 node_1 netRa14 26947.21182679576
Lbr14 netRa14 netL14 4.682210546303704e-11
Rbbr14 netL14 node_3 158255.1136047566
Cbr14 netL14 node_3 1.1202002197713253e-20

* Branch 15
Rabr15 node_1 netRa15  52.5961858777642
Lbr15 netRa15 netL15 1.6938904162108628e-13
Rbbr15 netL15 node_3  485.5979524712106
Cbr15 netL15 node_3 3.3129754960377035e-18

* Branch 16
Rabr16 node_1 netRa16 6503629.442874395
Lbr16 netRa16 netL16  1.035162587987019e-09
Rbbr16 netL16 node_3 6765580.512603145
Cbr16 netL16 node_3  2.3507710585681957e-23

* Branch 17
Rabr17 node_1 netRa17  580147.8920820685
Lbr17 netRa17 netL17 8.848053040551065e-11
Rbbr17 netL17 node_3  602018.2764071036
Cbr17 netL17 node_3 2.5291024230739794e-22

* Branch 18
Rabr18 node_1 netRa18 137.27046989941582
Lbr18 netRa18 netL18 6.23017313053251e-13
Rbbr18 netL18 node_3 5131.163738664318
Cbr18 netL18 node_3 9.51262191132007e-19

* Branch 19
Rabr19 node_1 netRa19 8022013.862322145
Lbr19 netRa19 netL19  1.9640253279607016e-09
Rbbr19 netL19 node_3 8823070.496143522
Cbr19 netL19 node_3  2.774321327686526e-23

* Branch 20
Rabr20 node_1 netRa20 38240.989103754284
Lbr20 netRa20 netL20  9.498231071105714e-11
Rbbr20 netL20 node_3 429024.279860405
Cbr20 netL20 node_3  5.73706859304262e-21

* Branch 21
Rabr21 node_1 netRa21  36736.73747086625
Lbr21 netRa21 netL21 7.030406264492435e-11
Rbbr21 netL21 node_3  265387.23011200037
Cbr21 netL21 node_3 7.139558692539796e-21

* Branch 22
Rabr22 node_1 netRa22  82.1198143349312
Lbr22 netRa22 netL22  7.130497095507288e-13
Rbbr22 netL22 node_3  12558.033874304567
Cbr22 netL22 node_3  7.900625425120072e-19

* Branch 23
Rabr23 node_1 netRa23 41841.57390785672
Lbr23 netRa23 netL23  3.400236039313734e-12
Rbbr23 netL23 node_3 42332.65853064579
Cbr23 netL23 node_3  1.9078506029164446e-21

* Branch 24
Rabr24 node_1 netRa24  1482.3956622558703
Lbr24 netRa24 netL24  1.991476726491402e-11
Rbbr24 netL24 node_3  539913.823299124
Cbr24 netL24 node_3  2.7658268243624383e-20

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 508.78668700326176
Lbr0 netRa0 netL0 1.0162691352386342e-12
Rbbr0 netL0 node_4 3014.3887990755557
Cbr0 netL0 node_4 6.785555499480596e-19

* Branch 1
Rabr1 node_1 netRa1  2518.603838329864
Lbr1 netRa1 netL1  2.0302239908707417e-12
Rbbr1 netL1 node_4  4643.782418478498
Cbr1 netL1 node_4  1.8124593105870242e-19

* Branch 2
Rabr2 node_1 netRa2  1681270.4490885255
Lbr2 netRa2 netL2 8.007353516911834e-10
Rbbr2 netL2 node_4  2157673.781870917
Cbr2 netL2 node_4 2.205712970941372e-22

* Branch 3
Rabr3 node_1 netRa3 6952386.251949257
Lbr3 netRa3 netL3 5.361655772343879e-10
Rbbr3 netL3 node_4 7004172.660435655
Cbr3 netL3 node_4 1.1016310980201708e-23

* Branch 4
Rabr4 node_1 netRa4  15.931494351366737
Lbr4 netRa4 netL4  7.726731595649137e-13
Rbbr4 netL4 node_4  167470.05261305178
Cbr4 netL4 node_4  9.871799656310793e-19

* Branch 5
Rabr5 node_1 netRa5  154449.8544833236
Lbr5 netRa5 netL5 9.971376894688715e-11
Rbbr5 netL5 node_4  239496.35722151332
Cbr5 netL5 node_4 2.6841672822287003e-21

* Branch 6
Rabr6 node_1 netRa6 16964.32385036715
Lbr6 netRa6 netL6  8.093980603579611e-11
Rbbr6 netL6 node_4 526226.8908967449
Cbr6 netL6 node_4  8.72712279748986e-21

* Branch 7
Rabr7 node_1 netRa7 725622.995120041
Lbr7 netRa7 netL7  1.0184609666451618e-09
Rbbr7 netL7 node_4 2701935.8473583534
Cbr7 netL7 node_4  5.184511498517828e-22

* Branch 8
Rabr8 node_1 netRa8  522942.25402593496
Lbr8 netRa8 netL8 5.807422455470927e-11
Rbbr8 netL8 node_4  531943.3020647692
Cbr8 netL8 node_4 2.0810794098654821e-22

* Branch 9
Rabr9 node_1 netRa9 75.11495226173666
Lbr9 netRa9 netL9 7.913406691004769e-13
Rbbr9 netL9 node_4 14001.436389354107
Cbr9 netL9 node_4 8.871274055496859e-19

* Branch 10
Rabr10 node_1 netRa10 23370962.240110207
Lbr10 netRa10 netL10  3.620365954470082e-09
Rbbr10 netL10 node_4 24183660.892652012
Cbr10 netL10 node_4  6.404111924292728e-24

* Branch 11
Rabr11 node_1 netRa11  103710.32593668677
Lbr11 netRa11 netL11  1.660664945056263e-10
Rbbr11 netL11 node_4  493021.9442405779
Cbr11 netL11 node_4  3.272476894686753e-21

* Branch 12
Rabr12 node_1 netRa12 908861.8227571636
Lbr12 netRa12 netL12 3.2011729829499184e-10
Rbbr12 netL12 node_4 1077862.6672474765
Cbr12 netL12 node_4 3.275125652888308e-22

* Branch 13
Rabr13 node_1 netRa13 35.206547645298166
Lbr13 netRa13 netL13  7.610404260486583e-13
Rbbr13 netL13 node_4 19054.8468205753
Cbr13 netL13 node_4  8.578218782590139e-19

* Branch 14
Rabr14 node_1 netRa14 30314.92669308051
Lbr14 netRa14 netL14 5.267465424965948e-11
Rbbr14 netL14 node_4 178038.51508979764
Cbr14 netL14 node_4 9.957439454383384e-21

* Branch 15
Rabr15 node_1 netRa15  59.170895814087636
Lbr15 netRa15 netL15 1.905627132228037e-13
Rbbr15 netL15 node_4  546.2972741244225
Cbr15 netL15 node_4 2.944865062558032e-18

* Branch 16
Rabr16 node_1 netRa16 7317250.29876917
Lbr16 netRa16 netL16  1.164607213706955e-09
Rbbr16 netL16 node_4 7611943.34397322
Cbr16 netL16 node_4  2.0892896693130357e-23

* Branch 17
Rabr17 node_1 netRa17  652647.3064064401
Lbr17 netRa17 netL17 9.953898960822332e-11
Rbbr17 netL17 node_4  677251.4127395508
Cbr17 netL17 node_4 2.248183953928113e-22

* Branch 18
Rabr18 node_1 netRa18 154.42938350738962
Lbr18 netRa18 netL18 7.008943533088141e-13
Rbbr18 netL18 node_4 5772.553146982343
Cbr18 netL18 node_4 8.455665013829686e-19

* Branch 19
Rabr19 node_1 netRa19 9024990.079379758
Lbr19 netRa19 netL19  2.2095478794445178e-09
Rbbr19 netL19 node_4 9926172.192495458
Cbr19 netL19 node_4  2.46596957566184e-23

* Branch 20
Rabr20 node_1 netRa20 43021.176473437634
Lbr20 netRa20 netL20  1.0685496783240038e-10
Rbbr20 netL20 node_4 482650.65424211277
Cbr20 netL20 node_4  5.099620357073807e-21

* Branch 21
Rabr21 node_1 netRa21  41328.92599012883
Lbr21 netRa21 netL21 7.90920810342737e-11
Rbbr21 netL21 node_4  298560.20490454964
Cbr21 netL21 node_4 6.346269704390805e-21

* Branch 22
Rabr22 node_1 netRa22  92.38490482229848
Lbr22 netRa22 netL22  8.021808908026702e-13
Rbbr22 netL22 node_4  14127.767269205162
Cbr22 netL22 node_4  7.02277831460328e-19

* Branch 23
Rabr23 node_1 netRa23 47072.20989443224
Lbr23 netRa23 netL23  3.825282175380209e-12
Rbbr23 netL23 node_4 47624.67976064109
Cbr23 netL23 node_4  1.6958431737222404e-21

* Branch 24
Rabr24 node_1 netRa24  1667.7066277704953
Lbr24 netRa24 netL24  2.2404092726991972e-11
Rbbr24 netL24 node_4  607397.2493348238
Cbr24 netL24 node_4  2.4585148650498324e-20

.ends


* Y'22
.subckt yp22 node_2 node_ref
* Branch 0
Rabr0 node_2 netRa0  440.18783349292937
Lbr0 netRa0 netL0  2.0257106439116213e-12
Rbbr0 netL0 node_ref  12318.95316035401
Cbr0 netL0 node_ref  3.9491296554680645e-19

* Branch 1
Rabr1 node_2 netRa1  36.18401201559627
Lbr1 netRa1 netL1  1.9068768674589719e-13
Rbbr1 netL1 node_ref  1763.2213924140387
Cbr1 netL1 node_ref  4.130103117776678e-18

* Branch 2
Rabr2 node_2 netRa2  60500.57049056161
Lbr2 netRa2 netL2  1.1371500093511289e-10
Rbbr2 netL2 node_ref  328466.0956929684
Cbr2 netL2 node_ref  5.738780442180008e-21

* Branch 3
Rabr3 node_2 netRa3  897.3637513905778
Lbr3 netRa3 netL3 1.2073563884102585e-11
Rbbr3 netL3 node_ref  187181.89699780935
Cbr3 netL3 node_ref 6.58496748951499e-20

* Branch 4
Rabr4 node_2 netRa4  1.7285648681059023
Lbr4 netRa4 netL4 1.0874065437730325e-13
Rbbr4 netL4 node_ref  4680.601431655105
Cbr4 netL4 node_ref 7.012633102788394e-18

* Branch 5
Rabr5 node_2 netRa5 3834.1552380487806
Lbr5 netRa5 netL5  3.199608297131588e-11
Rbbr5 netL5 node_ref 339477.7107802046
Cbr5 netL5 node_ref  2.329042410120042e-20

* Branch 6
Rabr6 node_2 netRa6  3779.759838505421
Lbr6 netRa6 netL6 2.267427715549704e-11
Rbbr6 netL6 node_ref  181440.11078362685
Cbr6 netL6 node_ref 3.152015112601641e-20

* Branch 7
Rabr7 node_2 netRa7  1137808.6997073893
Lbr7 netRa7 netL7 7.114691949144688e-10
Rbbr7 netL7 node_ref  1753541.4928296371
Cbr7 netL7 node_ref 3.562802151596418e-22

* Branch 8
Rabr8 node_2 netRa8  1011.9185892200868
Lbr8 netRa8 netL8 1.1782875909460213e-12
Rbbr8 netL8 node_ref  2871.0093285853736
Cbr8 netL8 node_ref 3.925174937073315e-19

* Branch 9
Rabr9 node_2 netRa9 106446.58131351073
Lbr9 netRa9 netL9 2.94830386664819e-11
Rbbr9 netL9 node_ref 118062.78614029007
Cbr9 netL9 node_ref 2.3553998865951004e-21

* Branch 10
Rabr10 node_2 netRa10  1660811.1720622082
Lbr10 netRa10 netL10  8.982780918968519e-10
Rbbr10 netL10 node_ref  2365551.375358388
Cbr10 netL10 node_ref  2.2881776825087312e-22

* Branch 11
Rabr11 node_2 netRa11  31349.806760957454
Lbr11 netRa11 netL11 9.973509184139513e-11
Rbbr11 netL11 node_ref  485588.42035904265
Cbr11 netL11 node_ref 6.454984867715862e-21

* Branch 12
Rabr12 node_2 netRa12  11843.920711895338
Lbr12 netRa12 netL12  4.0284209893289845e-11
Rbbr12 netL12 node_ref  221313.49535852554
Cbr12 netL12 node_ref  1.5710494977556728e-20

* Branch 13
Rabr13 node_2 netRa13  2.0718425112849475
Lbr13 netRa13 netL13 1.0349789933627387e-13
Rbbr13 netL13 node_ref  4531.645815044048
Cbr13 netL13 node_ref 6.316519934196353e-18

* Branch 14
Rabr14 node_2 netRa14  1636659.634887984
Lbr14 netRa14 netL14 3.788428227307873e-10
Rbbr14 netL14 node_ref  1775015.6983208675
Cbr14 netL14 node_ref 1.3006199682296691e-22

* Branch 15
Rabr15 node_2 netRa15  0.42428220135429734
Lbr15 netRa15 netL15  1.1585953470691502e-14
Rbbr15 netL15 node_ref 66.64953890569122
Cbr15 netL15 node_ref  5.466568973988867e-17

* Branch 16
Rabr16 node_2 netRa16  220771.34187620037
Lbr16 netRa16 netL16  4.1661141749438575e-10
Rbbr16 netL16 node_ref  1483284.3721981396
Cbr16 netL16 node_ref  1.2840563222736563e-21

* Branch 17
Rabr17 node_2 netRa17 233823.01829479952
Lbr17 netRa17 netL17  6.160181121173909e-11
Rbbr17 netL17 node_ref 260093.44019806923
Cbr17 netL17 node_ref  1.0099771849596121e-21

* Branch 18
Rabr18 node_2 netRa18 1952.946134878048
Lbr18 netRa18 netL18  6.599543044654041e-12
Rbbr18 netL18 node_ref 36758.252020385415
Cbr18 netL18 node_ref  8.736826399425266e-20

* Branch 19
Rabr19 node_2 netRa19 3535555.8808041643
Lbr19 netRa19 netL19 1.1717694231578305e-09
Rbbr19 netL19 node_ref 4182824.076673481
Cbr19 netL19 node_ref 7.92561332972382e-23

* Branch 20
Rabr20 node_2 netRa20 157119.39317379048
Lbr20 netRa20 netL20  1.0046931652867288e-10
Rbbr20 netL20 node_ref 264256.57920862356
Cbr20 netL20 node_ref  2.414124353787986e-21

* Branch 21
Rabr21 node_2 netRa21  18868037.368667074
Lbr21 netRa21 netL21 6.714730172490403e-10
Rbbr21 netL21 node_ref  18909047.375857674
Cbr21 netL21 node_ref 1.8817039676341987e-24

* Branch 22
Rabr22 node_2 netRa22 0.7179351635411342
Lbr22 netRa22 netL22 1.1160864516501584e-13
Rbbr22 netL22 node_ref  24773.402707195117
Cbr22 netL22 node_ref 5.080954485714095e-18

* Branch 23
Rabr23 node_2 netRa23  9792.339431237766
Lbr23 netRa23 netL23  9.586179515482856e-13
Rbbr23 netL23 node_ref  9961.416214062727
Cbr23 netL23 node_ref  9.901248702221964e-21

* Branch 24
Rabr24 node_2 netRa24 9652.598114379312
Lbr24 netRa24 netL24  2.1868081623301938e-11
Rbbr24 netL24 node_ref 97857.57931065583
Cbr24 netL24 node_ref  2.2765763620637947e-20

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 395.7228754330737
Lbr0 netRa0 netL0 7.904314928937305e-13
Rbbr0 netL0 node_3 2344.524756208284
Cbr0 netL0 node_3 8.724286832852998e-19

* Branch 1
Rabr1 node_2 netRa1  1958.9155693179905
Lbr1 netRa1 netL1  1.5790640251926527e-12
Rbbr1 netL1 node_3  3611.8329162376403
Cbr1 netL1 node_3  2.3303030331609623e-19

* Branch 2
Rabr2 node_2 netRa2  1307656.7798530895
Lbr2 netRa2 netL2 6.227950505074677e-10
Rbbr2 netL2 node_3  1678193.1993315585
Cbr2 netL2 node_3 2.8359122226987322e-22

* Branch 3
Rabr3 node_2 netRa3 5407459.406045928
Lbr3 netRa3 netL3 4.170196865408143e-10
Rbbr3 netL3 node_3 5447737.756365688
Cbr3 netL3 node_3 1.4163646857917306e-23

* Branch 4
Rabr4 node_2 netRa4  12.391148283760398
Lbr4 netRa4 netL4  6.009680336807378e-13
Rbbr4 netL4 node_3  130255.00634764571
Cbr4 netL4 node_3  1.2692313413141574e-18

* Branch 5
Rabr5 node_2 netRa5  120127.85820748762
Lbr5 netRa5 netL5 7.755526611553081e-11
Rbbr5 netL5 node_3  186275.22343834434
Cbr5 netL5 node_3 3.451066498213454e-21

* Branch 6
Rabr6 node_2 netRa6 13194.493775266508
Lbr6 netRa6 netL6  6.295324233627373e-11
Rbbr6 netL6 node_3 409287.7723315674
Cbr6 netL6 node_3  1.1220575400742e-20

* Branch 7
Rabr7 node_2 netRa7 564376.030925027
Lbr7 netRa7 netL7  7.92137298810995e-10
Rbbr7 netL7 node_3 2101505.052171803
Cbr7 netL7 node_3  6.665780215791926e-22

* Branch 8
Rabr8 node_2 netRa8  406732.76714367786
Lbr8 netRa8 netL8 4.5168839264953136e-11
Rbbr8 netL8 node_3  413733.58331487497
Cbr8 netL8 node_3 2.675674663630597e-22

* Branch 9
Rabr9 node_2 netRa9 58.42273176467365
Lbr9 netRa9 netL9 6.154871833706237e-13
Rbbr9 netL9 node_3 10890.007871367907
Cbr9 netL9 node_3 1.1405923873815813e-18

* Branch 10
Rabr10 node_2 netRa10 18177342.8469882
Lbr10 netRa10 netL10  2.8158376427102853e-09
Rbbr10 netL10 node_3 18809443.16801886
Cbr10 netL10 node_3  8.233914480223114e-24

* Branch 11
Rabr11 node_2 netRa11  80663.85074858849
Lbr11 netRa11 netL11  1.291630419178014e-10
Rbbr11 netL11 node_3  383461.7797056161
Cbr11 netL11 node_3  4.207460474208194e-21

* Branch 12
Rabr12 node_2 netRa12 706894.2461978458
Lbr12 netRa12 netL12 2.489804966417441e-10
Rbbr12 netL12 node_3 838339.4245885041
Cbr12 netL12 node_3 4.210862941627179e-22

* Branch 13
Rabr13 node_2 netRa13 27.38285940757869
Lbr13 netRa13 netL13  5.919203182567388e-13
Rbbr13 netL13 node_3 14820.440316128193
Cbr13 netL13 node_3  1.1029138692678816e-18

* Branch 14
Rabr14 node_2 netRa14 23578.532615953078
Lbr14 netRa14 netL14 4.096930085155444e-11
Rbbr14 netL14 node_3 138474.09273126512
Cbr14 netL14 node_3 1.2802348593398031e-20

* Branch 15
Rabr15 node_2 netRa15  46.021764917416526
Lbr15 netRa15 netL15 1.4821557587400724e-13
Rbbr15 netL15 node_3  424.89852047908744
Cbr15 netL15 node_3 3.786252824356571e-18

* Branch 16
Rabr16 node_2 netRa16 5691010.054131387
Lbr16 netRa16 netL16  9.057923374960781e-10
Rbbr16 netL16 node_3 5920216.471007599
Cbr16 netL16 node_3  2.686360765671023e-23

* Branch 17
Rabr17 node_2 netRa17  507628.2724491482
Lbr17 netRa17 netL17 7.74203512191131e-11
Rbbr17 netL17 node_3  526764.8456194011
Cbr17 netL17 node_3 2.890411292418735e-22

* Branch 18
Rabr18 node_2 netRa18 120.11162714448747
Lbr18 netRa18 netL18 5.451401282145451e-13
Rbbr18 netL18 node_3 4489.769223765927
Cbr18 netL18 node_3 1.0871568459633502e-18

* Branch 19
Rabr19 node_2 netRa19 7019395.105568854
Lbr19 netRa19 netL19  1.7185357781013893e-09
Rbbr19 netL19 node_3 7720317.490252877
Cbr19 netL19 node_3  3.170564288840564e-23

* Branch 20
Rabr20 node_2 netRa20 33460.81986808859
Lbr20 netRa20 netL20  8.310961356965314e-11
Rbbr20 netL20 node_3 375397.4121619812
Cbr20 netL20 node_3  6.55664545587564e-21

* Branch 21
Rabr21 node_2 netRa21  32144.72018595644
Lbr21 netRa21 netL21 6.151615022362634e-11
Rbbr21 netL21 node_3  232214.0572207498
Cbr21 netL21 node_3 8.159481242303913e-21

* Branch 22
Rabr22 node_2 netRa22  71.85479558589158
Lbr22 netRa22 netL22  6.239183820525139e-13
Rbbr22 netL22 node_3  10988.282615190143
Cbr22 netL22 node_3  9.029287897899093e-19

* Branch 23
Rabr23 node_2 netRa23 36611.7525725535
Lbr23 netRa23 netL23  2.9752223336456446e-12
Rbbr23 netL23 node_3 37041.451788223356
Cbr23 netL23 node_3  2.1803678692417456e-21

* Branch 24
Rabr24 node_2 netRa24  1297.08392334097
Lbr24 netRa24 netL24  1.742540152675766e-11
Rbbr24 netL24 node_3  472428.4094620146
Cbr24 netL24 node_3  3.160948691928956e-20

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 339.1910249504919
Lbr0 netRa0 netL0 6.775127246813013e-13
Rbbr0 netL0 node_4 2009.5927754694155
Cbr0 netL0 node_4 1.01783345894121e-18

* Branch 1
Rabr1 node_2 netRa1  1679.0713647849905
Lbr1 netRa1 netL1  1.353483657770896e-12
Rbbr1 netL1 node_4  3095.857333880094
Cbr1 netL1 node_4  2.7186853433963785e-19

* Branch 2
Rabr2 node_2 netRa2  1120852.2377281701
Lbr2 netRa2 netL2 5.338251828568357e-10
Rbbr2 netL2 node_4  1438454.8879834444
Cbr2 netL2 node_4 3.3085507986437155e-22

* Branch 3
Rabr3 node_2 netRa3 4634929.707818214
Lbr3 netRa3 netL3 3.5744410344224695e-10
Rbbr3 netL3 node_4 4669454.013302447
Cbr3 netL3 node_4 1.6524444808152513e-23

* Branch 4
Rabr4 node_2 netRa4  10.620989988773522
Lbr4 netRa4 netL4  5.151154609226296e-13
Rbbr4 netL4 node_4  111646.94577264998
Cbr4 netL4 node_4  1.480769887858611e-18

* Branch 5
Rabr5 node_2 netRa5  102966.43018721818
Lbr5 netRa5 netL5 6.647587953017029e-11
Rbbr5 netL5 node_4  159664.23228283814
Cbr5 netL5 node_4 4.026258525798773e-21

* Branch 6
Rabr6 node_2 netRa6 11309.597538073069
Lbr6 netRa6 netL6  5.395994458430222e-11
Rbbr6 netL6 node_4 350817.4922531263
Cbr6 netL6 node_4  1.3090663866366125e-20

* Branch 7
Rabr7 node_2 netRa7 483751.21424966614
Lbr7 netRa7 netL7  6.789743596779798e-10
Rbbr7 netL7 node_4 1801287.6626362794
Cbr7 netL7 node_4  7.776743216621798e-22

* Branch 8
Rabr8 node_2 netRa8  348628.75038747804
Lbr8 netRa8 netL8 3.871620118484713e-11
Rbbr8 netL8 node_4  354629.4550439576
Cbr8 netL8 node_4 3.121612899341386e-22

* Branch 9
Rabr9 node_2 netRa9 50.07661729410075
Lbr9 netRa9 netL9 5.275604638780006e-13
Rbbr9 netL9 node_4 9334.295427316581
Cbr9 netL9 node_4 1.3306910693749436e-18

* Branch 10
Rabr10 node_2 netRa10 15580499.696818648
Lbr10 netRa10 netL10  2.4135678187668344e-09
Rbbr10 netL10 node_4 16122299.470703954
Cbr10 netL10 node_4  9.606301639087272e-24

* Branch 11
Rabr11 node_2 netRa11  69140.44056378515
Lbr11 netRa11 netL11  1.1071108931559147e-10
Rbbr11 netL11 node_4  328681.1125411363
Cbr11 netL11 node_4  4.908706266249837e-21

* Branch 12
Rabr12 node_2 netRa12 605909.377819562
Lbr12 netRa12 netL12 2.1341176436952952e-10
Rbbr12 netL12 node_4 718576.5740979448
Cbr12 netL12 node_4 4.912671679871142e-22

* Branch 13
Rabr13 node_2 netRa13 23.47103666661165
Lbr13 netRa13 netL13  5.073602752913396e-13
Rbbr13 netL13 node_4 12703.228832046369
Cbr13 netL13 node_4  1.2867328386129878e-18

* Branch 14
Rabr14 node_2 netRa14 20210.087390617675
Lbr14 netRa14 netL14 3.51164352859917e-11
Rbbr14 netL14 node_4 118691.79721049868
Cbr14 netL14 node_4 1.4936124785373548e-20

* Branch 15
Rabr15 node_2 netRa15  39.4472006593484
Lbr15 netRa15 netL15 1.2704180787381894e-13
Rbbr15 netL15 node_4  364.198375898689
Cbr15 netL15 node_4 4.417298771012099e-18

* Branch 16
Rabr16 node_2 netRa16 4877976.095637949
Lbr16 netRa16 netL16  7.76389794017217e-10
Rbbr16 netL16 node_4 5074438.206991164
Cbr16 netL16 node_4  3.1341141792111317e-23

* Branch 17
Rabr17 node_2 netRa17  435095.67304095393
Lbr17 netRa17 netL17 6.635920878813455e-11
Rbbr17 netL17 node_4  451498.44776396395
Cbr17 netL17 node_4 3.3723081778305943e-22

* Branch 18
Rabr18 node_2 netRa18 102.9529405673915
Lbr18 netRa18 netL18 4.67263005421131e-13
Rbbr18 netL18 node_4 3848.369786772258
Cbr18 netL18 node_4 1.2683494749912018e-18

* Branch 19
Rabr19 node_2 netRa19 6016509.345521548
Lbr19 netRa19 netL19  1.4730159646802592e-09
Rbbr19 netL19 node_4 6617299.45337607
Cbr19 netL19 node_4  3.699090050095652e-23

* Branch 20
Rabr20 node_2 netRa20 28680.589454122222
Lbr20 netRa20 netL20  7.123670298476983e-11
Rbbr20 netL20 node_4 321769.35442255746
Cbr20 netL20 node_4  7.649434656789711e-21

* Branch 21
Rabr21 node_2 netRa21  27552.60545687094
Lbr21 netRa21 netL21 5.272809098464529e-11
Rbbr21 netL21 node_4  199040.43710851905
Cbr21 netL21 node_4 9.519400851639413e-21

* Branch 22
Rabr22 node_2 netRa22  61.58986277225151
Lbr22 netRa22 netL22  5.347872161947751e-13
Rbbr22 netL22 node_4  9418.522583827988
Cbr22 netL22 node_4  1.053416850987761e-18

* Branch 23
Rabr23 node_2 netRa23 31381.407071909936
Lbr23 netRa23 netL23  2.5501859614556862e-12
Rbbr23 netL23 node_4 31749.720467435494
Cbr23 netL23 node_4  2.543773247231517e-21

* Branch 24
Rabr24 node_2 netRa24  1111.8028931157103
Lbr24 netRa24 netL24  1.4936061125504272e-11
Rbbr24 netL24 node_4  404932.07435545523
Cbr24 netL24 node_4  3.6877724968960895e-20

.ends


* Y'33
.subckt yp33 node_3 node_ref
* Branch 0
Rabr0 node_3 netRa0  645.4971255792519
Lbr0 netRa0 netL0  1.5747615938397319e-12
Rbbr0 netL0 node_ref  5412.900219240011
Cbr0 netL0 node_ref  4.640003860947413e-19

* Branch 1
Rabr1 node_3 netRa1  174.083594260938
Lbr1 netRa1 netL1  2.8394519223227844e-13
Rbbr1 netL1 node_ref  803.9548920816143
Cbr1 netL1 node_ref  2.218575796971884e-18

* Branch 2
Rabr2 node_3 netRa2  1482569.1322433155
Lbr2 netRa2 netL2  4.3422383214595164e-10
Rbbr2 netL2 node_ref  1641628.115297933
Cbr2 netL2 node_ref  1.7849200063545392e-22

* Branch 3
Rabr3 node_3 netRa3 21192.615638784802
Lbr3 netRa3 netL3 2.0917122595488706e-11
Rbbr3 netL3 node_ref 47210.39190741267
Cbr3 netL3 node_ref 2.1047804114196334e-20

* Branch 4
Rabr4 node_3 netRa4  4.887633964391439
Lbr4 netRa4 netL4 1.2252395232172819e-13
Rbbr4 netL4 node_ref  2954.063110171491
Cbr4 netL4 node_ref 6.2157469120128884e-18

* Branch 5
Rabr5 node_3 netRa5 18549.2928077763
Lbr5 netRa5 netL5 3.611096993057943e-11
Rbbr5 netL5 node_ref 113042.04374000849
Cbr5 netL5 node_ref 1.7447230604516023e-20

* Branch 6
Rabr6 node_3 netRa6 40485.64392037922
Lbr6 netRa6 netL6  7.596623339509036e-11
Rbbr6 netL6 node_ref 232829.72668709705
Cbr6 netL6 node_ref  7.937510944876781e-21

* Branch 7
Rabr7 node_3 netRa7 4902271.407473896
Lbr7 netRa7 netL7  3.6333020493172212e-09
Rbbr7 netL7 node_ref 8628631.235758683
Cbr7 netL7 node_ref  8.580506922482819e-23

* Branch 8
Rabr8 node_3 netRa8 5373.871684409021
Lbr8 netRa8 netL8  6.528512933774881e-12
Rbbr8 netL8 node_ref 16105.840269081593
Cbr8 netL8 node_ref  7.289975578419429e-20

* Branch 9
Rabr9 node_3 netRa9  15275051.530689776
Lbr9 netRa9 netL9 7.759386310090133e-10
Rbbr9 netL9 node_ref  15330855.945883859
Cbr9 netL9 node_ref 3.3110096195546786e-24

* Branch 10
Rabr10 node_3 netRa10 675768566.9935782
Lbr10 netRa10 netL10  7.718105011435312e-08
Rbbr10 netL10 node_ref 688543231.5013634
Cbr10 netL10 node_ref  1.658484805872133e-25

* Branch 11
Rabr11 node_3 netRa11 119417.13995187839
Lbr11 netRa11 netL11  3.499651957908825e-10
Rbbr11 netL11 node_ref 1589395.240519359
Cbr11 netL11 node_ref  1.8187859614971738e-21

* Branch 12
Rabr12 node_3 netRa12  242064.03533510264
Lbr12 netRa12 netL12  2.3140102487063806e-10
Rbbr12 netL12 node_ref  574918.1281425629
Cbr12 netL12 node_ref  1.6729936220067845e-21

* Branch 13
Rabr13 node_3 netRa13  2.326481288794787
Lbr13 netRa13 netL13 1.1710402311773368e-13
Rbbr13 netL13 node_ref  5149.680452224358
Cbr13 netL13 node_ref 5.582644159713205e-18

* Branch 14
Rabr14 node_3 netRa14  45447.722205303486
Lbr14 netRa14 netL14 1.9476989025526022e-11
Rbbr14 netL14 node_ref  58587.705987354864
Cbr14 netL14 node_ref 7.279138771495933e-21

* Branch 15
Rabr15 node_3 netRa15  1.7972140113213586
Lbr15 netRa15 netL15  1.674081579908367e-14
Rbbr15 netL15 node_ref 128.76849734102035
Cbr15 netL15 node_ref  3.8118307293345036e-17

* Branch 16
Rabr16 node_3 netRa16 45599.57905211703
Lbr16 netRa16 netL16 5.017491328798671e-11
Rbbr16 netL16 node_ref 133917.36117464284
Cbr16 netL16 node_ref 8.260920334396147e-21

* Branch 17
Rabr17 node_3 netRa17  633572.3165689758
Lbr17 netRa17 netL17  8.13631900100307e-11
Rbbr17 netL17 node_ref  650559.0717714496
Cbr17 netL17 node_ref  1.97680176156884e-22

* Branch 18
Rabr18 node_3 netRa18  9666.208344223138
Lbr18 netRa18 netL18 9.005277761472031e-12
Rbbr18 netL18 node_ref  23247.80953500808
Cbr18 netL18 node_ref 3.950470202133758e-20

* Branch 19
Rabr19 node_3 netRa19  4365562.274915578
Lbr19 netRa19 netL19  1.4259478656641397e-09
Rbbr19 netL19 node_ref  5141850.597515443
Cbr19 netL19 node_ref  6.354191874160293e-23

* Branch 20
Rabr20 node_3 netRa20  322139.1873054985
Lbr20 netRa20 netL20 1.665536370345292e-10
Rbbr20 netL20 node_ref  465808.02130670013
Cbr20 netL20 node_ref 1.1078479077197043e-21

* Branch 21
Rabr21 node_3 netRa21 63116.528836429716
Lbr21 netRa21 netL21  6.07664718929575e-11
Rbbr21 netL21 node_ref 163034.19905007145
Cbr21 netL21 node_ref  5.87569485803929e-21

* Branch 22
Rabr22 node_3 netRa22 2.195563684081517
Lbr22 netRa22 netL22 1.2396125379603616e-13
Rbbr22 netL22 node_ref 65559.34359494748
Cbr22 netL22 node_ref 4.5743569436789524e-18

* Branch 23
Rabr23 node_3 netRa23  1372.819700898355
Lbr23 netRa23 netL23  6.796343745026638e-13
Rbbr23 netL23 node_ref  1998.086953244281
Cbr23 netL23 node_ref  2.574830239296998e-19

* Branch 24
Rabr24 node_3 netRa24 3692.6063836438934
Lbr24 netRa24 netL24  2.4556597284798925e-11
Rbbr24 netL24 node_ref 285368.0692532492
Cbr24 netL24 node_ref  2.2200855845606926e-20

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 621.8501936996532
Lbr0 netRa0 netL0 1.2421065536502092e-12
Rbbr0 netL0 node_4 3684.252957067631
Cbr0 netL0 node_4 5.551819242611099e-19

* Branch 1
Rabr1 node_3 netRa1  3078.292170277253
Lbr1 netRa1 netL1  2.481385132994093e-12
Rbbr1 netL1 node_4  5675.734445493021
Cbr1 netL1 node_4  1.482922023692054e-19

* Branch 2
Rabr2 node_3 netRa2  2054906.067694486
Lbr2 netRa2 netL2 9.786817277796095e-10
Rbbr2 netL2 node_4  2637177.32475402
Cbr2 netL2 node_4 1.8046522718831825e-22

* Branch 3
Rabr3 node_3 netRa3 8497205.730950043
Lbr3 netRa3 netL3 6.553077967181445e-10
Rbbr3 netL3 node_4 8560500.288410451
Cbr3 netL3 node_4 9.013595246671652e-24

* Branch 4
Rabr4 node_3 netRa4  19.47182628865752
Lbr4 netRa4 netL4  9.443783158359591e-13
Rbbr4 netL4 node_4  204685.6341736599
Cbr4 netL4 node_4  8.076926908616597e-19

* Branch 5
Rabr5 node_3 netRa5  188771.93307878645
Lbr5 netRa5 netL5 1.2187240190419712e-10
Rbbr5 netL5 node_4  292717.7496857921
Cbr5 netL5 node_4 2.196138624849146e-21

* Branch 6
Rabr6 node_3 netRa6 20734.167555997556
Lbr6 netRa6 netL6  9.892651982255423e-11
Rbbr6 netL6 node_4 643167.4825213051
Cbr6 netL6 node_4  7.140367229347556e-21

* Branch 7
Rabr7 node_3 netRa7 886874.60165284
Lbr7 netRa7 netL7  1.2447867749294485e-09
Rbbr7 netL7 node_4 3302366.9646469713
Cbr7 netL7 node_4  4.24186596316225e-22

* Branch 8
Rabr8 node_3 netRa8  639152.132618862
Lbr8 netRa8 netL8 7.0979646348415e-11
Rbbr8 netL8 node_4  650153.4171021653
Cbr8 netL8 node_4 1.7026996698899454e-22

* Branch 9
Rabr9 node_3 netRa9 91.80714579833665
Lbr9 netRa9 netL9 9.671941400039135e-13
Rbbr9 netL9 node_4 17112.870205132804
Cbr9 netL9 node_4 7.258315235489175e-19

* Branch 10
Rabr10 node_3 netRa10 28564358.37623192
Lbr10 netRa10 netL10  4.424880694856891e-09
Rbbr10 netL10 node_4 29557657.02978081
Cbr10 netL10 node_4  5.239769300702537e-24

* Branch 11
Rabr11 node_3 netRa11  126757.2779433239
Lbr11 netRa11 netL11  2.0297026283735479e-10
Rbbr11 netL11 node_4  602582.2681361982
Cbr11 netL11 node_4  2.6774784123606283e-21

* Branch 12
Rabr12 node_3 netRa12 1110835.8734155193
Lbr12 netRa12 netL12 3.912553239012902e-10
Rbbr12 netL12 node_4 1317392.4712353067
Cbr12 netL12 node_4 2.679632887403644e-22

* Branch 13
Rabr13 node_3 netRa13 43.03021086405141
Lbr13 netRa13 netL13  9.301604928882806e-13
Rbbr13 netL13 node_4 23289.261722997497
Cbr13 netL13 node_4  7.018542857098872e-19

* Branch 14
Rabr14 node_3 netRa14 37052.09684935743
Lbr14 netRa14 netL14 6.438037544005411e-11
Rbbr14 netL14 node_4 217601.93890173838
Cbr14 netL14 node_4 8.146936473762455e-21

* Branch 15
Rabr15 node_3 netRa15  72.31995938123761
Lbr15 netRa15 netL15 2.329102192940437e-13
Rbbr15 netL15 node_4  667.6976507102723
Cbr15 netL15 node_4 2.4094331342604176e-18

* Branch 16
Rabr16 node_3 netRa16 8942907.784173658
Lbr16 netRa16 netL16  1.423381237361842e-09
Rbbr16 netL16 node_4 9303090.242982265
Cbr16 netL16 node_4  1.709534545483593e-23

* Branch 17
Rabr17 node_3 netRa17  797705.5045307777
Lbr17 netRa17 netL17 1.2166082741699166e-10
Rbbr17 netL17 node_4  827777.2504140352
Cbr17 netL17 node_4 1.8393390302515943e-22

* Branch 18
Rabr18 node_3 netRa18 188.74682146319418
Lbr18 netRa18 netL18 8.566487340650796e-13
Rbbr18 netL18 node_4 7055.351799103551
Cbr18 netL18 node_4 6.918271177359345e-19

* Branch 19
Rabr19 node_3 netRa19 11030453.617862228
Lbr19 netRa19 netL19  2.7005570561701907e-09
Rbbr19 netL19 node_4 12131906.195792936
Cbr19 netL19 node_4  2.0176404464127192e-23

* Branch 20
Rabr20 node_3 netRa20 52581.442688475094
Lbr20 netRa20 netL20  1.306008261272721e-10
Rbbr20 netL20 node_4 589908.8499941806
Cbr20 netL20 node_4  4.1724084452205924e-21

* Branch 21
Rabr21 node_3 netRa21  50513.10526495849
Lbr21 netRa21 netL21 9.666812495307434e-11
Rbbr21 netL21 node_4  364907.2216162248
Cbr21 netL21 node_4 5.192402227475868e-21

* Branch 22
Rabr22 node_3 netRa22  112.91468535274404
Lbr22 netRa22 netL22  9.804432828830487e-13
Rbbr22 netL22 node_4  17267.304282150966
Cbr22 netL22 node_4  5.74590983389154e-19

* Branch 23
Rabr23 node_3 netRa23 57532.66491342991
Lbr23 netRa23 netL23  4.675345881266502e-12
Rbbr23 netL23 node_4 58207.90656977247
Cbr23 netL23 node_4  1.3875100536328836e-21

* Branch 24
Rabr24 node_3 netRa24  2038.243905246125
Lbr24 netRa24 netL24  2.738277773503915e-11
Rbbr24 netL24 node_4  742400.1412282359
Cbr24 netL24 node_4  2.0115126949899506e-20

.ends


* Y'44
.subckt yp44 node_4 node_ref
* Branch 0
Rabr0 node_4 netRa0  1102.7174314914473
Lbr0 netRa0 netL0  2.098875299282033e-12
Rbbr0 netL0 node_ref  6028.1938060556
Cbr0 netL0 node_ref  3.229651793236128e-19

* Branch 1
Rabr1 node_4 netRa1  128.91469158254023
Lbr1 netRa1 netL1  2.879821470497374e-13
Rbbr1 netL1 node_ref  1035.1613121796595
Cbr1 netL1 node_ref  2.4443391083942165e-18

* Branch 2
Rabr2 node_4 netRa2  457711.36479514156
Lbr2 netRa2 netL2  2.864870794363542e-10
Rbbr2 netL2 node_ref  682092.2582635963
Cbr2 netL2 node_ref  9.185159575144648e-22

* Branch 3
Rabr3 node_4 netRa3 8826.275978203239
Lbr3 netRa3 netL3 1.9772976667998604e-11
Rbbr3 netL3 node_ref 65133.31391975542
Cbr3 netL3 node_ref 3.4927187729413364e-20

* Branch 4
Rabr4 node_4 netRa4  3.83334196939648
Lbr4 netRa4 netL4 1.1936858519329505e-13
Rbbr4 netL4 node_ref  3355.7567528331733
Cbr4 netL4 node_ref 6.383326275585674e-18

* Branch 5
Rabr5 node_4 netRa5 56080.739779401985
Lbr5 netRa5 netL5 7.085333723621807e-11
Rbbr5 netL5 node_ref 175854.3518947195
Cbr5 netL5 node_ref 7.245275085006837e-21

* Branch 6
Rabr6 node_4 netRa6 22916062.44169336
Lbr6 netRa6 netL6  1.1685087192341058e-09
Rbbr6 netL6 node_ref 22997660.30557469
Cbr6 netL6 node_ref  2.216295711815287e-24

* Branch 7
Rabr7 node_4 netRa7 5891932.996206046
Lbr7 netRa7 netL7 2.3631192550120505e-09
Rbbr7 netL7 node_ref 7205599.855077251
Cbr7 netL7 node_ref 5.569305393178077e-23

* Branch 8
Rabr8 node_4 netRa8 8990.840700883551
Lbr8 netRa8 netL8  5.782449177901758e-12
Rbbr8 netL8 node_ref 14103.792217877963
Cbr8 netL8 node_ref  4.4778370580838694e-20

* Branch 9
Rabr9 node_4 netRa9  49779.58744851105
Lbr9 netRa9 netL9  3.283665172844791e-11
Rbbr9 netL9 node_ref  80763.01497220485
Cbr9 netL9 node_ref  8.246007547950216e-21

* Branch 10
Rabr10 node_4 netRa10 1839415.796315828
Lbr10 netRa10 netL10 1.485688579676037e-09
Rbbr10 netL10 node_ref 3580689.417853119
Cbr10 netL10 node_ref 2.2582731637299715e-22

* Branch 11
Rabr11 node_4 netRa11 260431.7884967161
Lbr11 netRa11 netL11  2.647529580893581e-10
Rbbr11 netL11 node_ref 649646.0882220423
Cbr11 netL11 node_ref  1.5573944813983722e-21

* Branch 12
Rabr12 node_4 netRa12  154165.30812142402
Lbr12 netRa12 netL12  2.5819740273002084e-10
Rbbr12 netL12 node_ref  807876.282258126
Cbr12 netL12 node_ref  2.0955629578427543e-21

* Branch 13
Rabr13 node_4 netRa13  1.9312706680914309
Lbr13 netRa13 netL13 1.1380933379029785e-13
Rbbr13 netL13 node_ref  5459.031500142727
Cbr13 netL13 node_ref 5.7448204222965565e-18

* Branch 14
Rabr14 node_4 netRa14  26277.95124255818
Lbr14 netRa14 netL14 1.501806764562925e-11
Rbbr14 netL14 node_ref  39767.39388161815
Cbr14 netL14 node_ref 1.4277964620602917e-20

* Branch 15
Rabr15 node_4 netRa15  1.5454401139317444
Lbr15 netRa15 netL15  1.5609006946038716e-14
Rbbr15 netL15 node_ref 115.40232127033917
Cbr15 netL15 node_ref  4.085947740657046e-17

* Branch 16
Rabr16 node_4 netRa16 53326.26688238849
Lbr16 netRa16 netL16 5.132770484466524e-11
Rbbr16 netL16 node_ref 132303.97428218165
Cbr16 netL16 node_ref 7.309431170722226e-21

* Branch 17
Rabr17 node_4 netRa17  414061.9039672748
Lbr17 netRa17 netL17  6.267009157066112e-11
Rbbr17 netL17 node_ref  429486.59758094803
Cbr17 netL17 node_ref  3.5299942439154505e-22

* Branch 18
Rabr18 node_4 netRa18  9258.551769585467
Lbr18 netRa18 netL18 8.402190783393743e-12
Rbbr18 netL18 node_ref  21607.06228573364
Cbr18 netL18 node_ref 4.1419350255062474e-20

* Branch 19
Rabr19 node_4 netRa19  5998621.569234493
Lbr19 netRa19 netL19  1.6976569949114295e-09
Rbbr19 netL19 node_ref  6799356.616869362
Cbr19 netL19 node_ref  4.1632399577100113e-23

* Branch 20
Rabr20 node_4 netRa20  195683.10429445075
Lbr20 netRa20 netL20 1.4048737693834367e-10
Rbbr20 netL20 node_ref  363834.1596895626
Cbr20 netL20 node_ref 1.968056129365019e-21

* Branch 21
Rabr21 node_4 netRa21 48702.168242274034
Lbr21 netRa21 netL21  5.300767106802256e-11
Rbbr21 netL21 node_ref 147171.83053465013
Cbr21 netL21 node_ref  7.353578007691922e-21

* Branch 22
Rabr22 node_4 netRa22 2.1706330645657026
Lbr22 netRa22 netL22 1.2051657853393978e-13
Rbbr22 netL22 node_ref 58486.73373474656
Cbr22 netL22 node_ref 4.705086836804274e-18

* Branch 23
Rabr23 node_4 netRa23  1215.3394575808538
Lbr23 netRa23 netL23  5.747256968311221e-13
Rbbr23 netL23 node_ref  1719.5248840174806
Cbr23 netL23 node_ref  2.852947930774962e-19

* Branch 24
Rabr24 node_4 netRa24  37207.94099466646
Lbr24 netRa24 netL24  5.0388264567845253e-11
Rbbr24 netL24 node_ref  162016.85270406833
Cbr24 netL24 node_ref  8.444039750566744e-21

.ends


.end
