* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 1588.9471354629384
Lbr0 netRa0 netL0 -9.817714433440466e-13
Rbbr0 netL0 0 -1982.8686402966084
Cbr0 netL0 0 -2.1612796083657685e-19

* Branch 1
Rabr1 node_1 netRa1 -1633201904740.1648
Lbr1 netRa1 netL1 0.0016921536386547812
Rbbr1 netL1 0 3918434021680.556
Cbr1 netL1 0 2.6429672309260165e-28

* Branch 2
Rabr2 node_1 netRa2 -361694178.1264218
Lbr2 netRa2 netL2 -7.294398913048427e-07
Rbbr2 netL2 0 2400120367.0507655
Cbr2 netL2 0 -8.880211455989857e-25

* Branch 3
Rabr3 node_1 netRa3 49370283.28002451
Lbr3 netRa3 netL3 3.475009057249854e-08
Rbbr3 netL3 0 -82540034.51781523
Cbr3 netL3 0 8.815242689963665e-24

* Branch 4
Rabr4 node_1 netRa4 -58142426.08026196
Lbr4 netRa4 netL4 -4.150973695985141e-09
Rbbr4 netL4 0 58533994.52865965
Cbr4 netL4 0 -1.2265850011291457e-24

* Branch 5
Rabr5 node_1 netRa5 2602611.277077282
Lbr5 netRa5 netL5 -5.153613979475081e-10
Rbbr5 netL5 0 -2734365.7244887003
Cbr5 netL5 0 -7.108910668175893e-23

* Branch 6
Rabr6 node_1 netRa6 -983521182513.7047
Lbr6 netRa6 netL6 0.0002912237123668366
Rbbr6 netL6 0 1097009556925.9934
Cbr6 netL6 0 2.6939998639935374e-28

* Branch 7
Rabr7 node_1 netRa7 455.3894017638663
Lbr7 netRa7 netL7 1.6276557598842337e-13
Rbbr7 netL7 0 -549.1158103472468
Cbr7 netL7 0 7.59783598014151e-19

* Branch 8
Rabr8 node_1 netRa8 3157.408169467105
Lbr8 netRa8 netL8 -1.6182672088391108e-12
Rbbr8 netL8 0 -4245.062119699056
Cbr8 netL8 0 -1.1121986259310061e-19

* Branch 9
Rabr9 node_1 netRa9 -612.9611836183382
Lbr9 netRa9 netL9 9.193839965030269e-13
Rbbr9 netL9 0 2455.537590047057
Cbr9 netL9 0 5.396700512128527e-19

* Branch 10
Rabr10 node_1 netRa10 369899257793.33234
Lbr10 netRa10 netL10 0.0002802488106937338
Rbbr10 netL10 0 -693506839275.9337
Cbr10 netL10 0 1.0950286500808124e-27

* Branch 11
Rabr11 node_1 netRa11 21845.238475881295
Lbr11 netRa11 netL11 8.279999353547912e-12
Rbbr11 netL11 0 -26745.65922358917
Cbr11 netL11 0 1.4482518391248816e-20

* Branch 12
Rabr12 node_1 netRa12 3880542.2251560586
Lbr12 netRa12 netL12 -3.4891107274974124e-10
Rbbr12 netL12 0 -3928331.6940910406
Cbr12 netL12 0 -2.2788174296430714e-23

* Branch 13
Rabr13 node_1 netRa13 -15928.686223765568
Lbr13 netRa13 netL13 -7.6985075952408e-12
Rbbr13 netL13 0 21776.95470306085
Cbr13 netL13 0 -2.2796728856453218e-20

* Branch 14
Rabr14 node_1 netRa14 39088.42441807922
Lbr14 netRa14 netL14 -4.841285373356898e-12
Rbbr14 netL14 0 -39997.4129234861
Cbr14 netL14 0 -3.0559428174996653e-21

* Branch 15
Rabr15 node_1 netRa15 -31221265535087.36
Lbr15 netRa15 netL15 -0.007535304925834823
Rbbr15 netL15 0 34069794581270.973
Cbr15 netL15 0 -7.084756601178615e-30

* Branch 16
Rabr16 node_1 netRa16 -29.696551058486257
Lbr16 netRa16 netL16 6.259858740444013e-14
Rbbr16 netL16 0 156.3071011441061
Cbr16 netL16 0 8.066239712068329e-18

* Branch 17
Rabr17 node_1 netRa17 -203.16454198463583
Lbr17 netRa17 netL17 -2.9009576587927123e-13
Rbbr17 netL17 0 1181.1581485218164
Cbr17 netL17 0 -1.7007561256816824e-18

* Branch 18
Rabr18 node_1 netRa18 5.501373650005231
Lbr18 netRa18 netL18 1.1433962808467956e-14
Rbbr18 netL18 0 40.20977984146593
Cbr18 netL18 0 5.163445772919673e-17

* Branch 19
Rabr19 node_1 netRa19 1.822579184032874
Lbr19 netRa19 netL19 2.6922249728502162e-12
Rbbr19 netL19 0 1014073.4885401423
Cbr19 netL19 0 2.163959372351423e-19

* Branch 20
Rabr20 node_1 netRa20 -73079962.45817956
Lbr20 netRa20 netL20 -2.100626033862185e-07
Rbbr20 netL20 0 1183782236.1721566
Cbr20 netL20 0 -2.5328394107190068e-24

* Branch 21
Rabr21 node_1 netRa21 1181372.8036314999
Lbr21 netRa21 netL21 2.9011433334724367e-09
Rbbr21 netL21 0 -14430780.522471026
Cbr21 netL21 0 1.7944814271927736e-22

* Branch 22
Rabr22 node_1 netRa22 -1109367.3712610272
Lbr22 netRa22 netL22 -2.705537870193153e-09
Rbbr22 netL22 0 13394694.079396812
Cbr22 netL22 0 -1.922200040104301e-22

* Branch 23
Rabr23 node_1 netRa23 3.2027793493043126
Lbr23 netRa23 netL23 1.154540453502919e-13
Rbbr23 netL23 0 4714.170123604154
Cbr23 netL23 0 4.9081794268272136e-18

* Branch 24
Rabr24 node_1 netRa24 -33657.54316800791
Lbr24 netRa24 netL24 -7.1825221418671966e-12
Rbbr24 netL24 0 36530.25353394228
Cbr24 netL24 0 -6.068495908677487e-21

* Branch 25
Rd node_1 0 1838.4552192525334

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -14068.149650445048
Lbr0 netRa0 netL0 -9.304249579618183e-12
Rbbr0 netL0 node_2 24997.659050898168
Cbr0 netL0 node_2 -5.019096915760049e-20

* Branch 1
Rabr1 node_1 netRa1 74161128216701.23
Lbr1 netRa1 netL1 -0.01754992879364137
Rbbr1 netL1 node_2 -79576345867220.17
Cbr1 netL1 node_2 -2.9735165192569e-30

* Branch 2
Rabr2 node_1 netRa2 17.703186390687247
Lbr2 netRa2 netL2 8.58527087635816e-13
Rbbr2 netL2 node_2 186132.4107205688
Cbr2 netL2 node_2 8.884605551912848e-19

* Branch 3
Rabr3 node_1 netRa3 -28366730.503201198
Lbr3 netRa3 netL3 4.497374537988834e-08
Rbbr3 netL3 node_2 115501686.30723193
Cbr3 netL3 node_2 1.2786676546829933e-23

* Branch 4
Rabr4 node_1 netRa4 174805.75842981064
Lbr4 netRa4 netL4 -1.1775341259264413e-09
Rbbr4 netL4 node_2 -6983935.112174665
Cbr4 netL4 node_2 -6.301819943113748e-22

* Branch 5
Rabr5 node_1 netRa5 50000.73422308884
Lbr5 netRa5 netL5 4.6249281122844404e-10
Rbbr5 netL5 node_2 -44400388.00524919
Cbr5 netL5 node_2 1.6421465962687632e-21

* Branch 6
Rabr6 node_1 netRa6 -131429173144.07864
Lbr6 netRa6 netL6 0.00027183556453430044
Rbbr6 netL6 node_2 862968926300.3029
Cbr6 netL6 node_2 2.3649384220103957e-27

* Branch 7
Rabr7 node_1 netRa7 -1017.6890137952681
Lbr7 netRa7 netL7 -1.521591636062863e-12
Rbbr7 netL7 node_2 8857.247902218494
Cbr7 netL7 node_2 -4.2145300989612294e-19

* Branch 8
Rabr8 node_1 netRa8 221.32868605003583
Lbr8 netRa8 netL8 1.3181385621721387e-12
Rbbr8 netL8 node_2 -1920627.9347843896
Cbr8 netL8 node_2 5.328620375578251e-19

* Branch 9
Rabr9 node_1 netRa9 20923.02508435117
Lbr9 netRa9 netL9 5.971927172340492e-11
Rbbr9 netL9 node_2 -365051.63880755805
Cbr9 netL9 node_2 1.0437543973478607e-20

* Branch 10
Rabr10 node_1 netRa10 -1525539021140.5413
Lbr10 netRa10 netL10 0.002363025239165184
Rbbr10 netL10 node_2 7064680075999.612
Cbr10 netL10 node_2 2.182141384192073e-28

* Branch 11
Rabr11 node_1 netRa11 234649.27475185032
Lbr11 netRa11 netL11 3.208641654786782e-10
Rbbr11 netL11 node_2 -961315.0608041008
Cbr11 netL11 node_2 1.5418498304421234e-21

* Branch 12
Rabr12 node_1 netRa12 15234586.469832871
Lbr12 netRa12 netL12 6.504004468382865e-09
Rbbr12 netL12 node_2 -19573591.886478808
Cbr12 netL12 node_2 2.2276095109923616e-23

* Branch 13
Rabr13 node_1 netRa13 -194792.268415142
Lbr13 netRa13 netL13 -3.444197056520512e-10
Rbbr13 netL13 node_2 1226506.9840190297
Cbr13 netL13 node_2 -1.5960648402585048e-21

* Branch 14
Rabr14 node_1 netRa14 -8.491559702577234
Lbr14 netRa14 netL14 8.915870766421362e-13
Rbbr14 netL14 node_2 11728.438654436193
Cbr14 netL14 node_2 7.296273459363355e-19

* Branch 15
Rabr15 node_1 netRa15 -3893893009474.2563
Lbr15 netRa15 netL15 -0.00907729074228034
Rbbr15 netL15 node_2 37066545063931.68
Cbr15 netL15 node_2 -6.29530054039314e-29

* Branch 16
Rabr16 node_1 netRa16 -37.89971878077015
Lbr16 netRa16 netL16 2.9972175930931246e-13
Rbbr16 netL16 node_2 1117.90219414303
Cbr16 netL16 node_2 2.0093108970126667e-18

* Branch 17
Rabr17 node_1 netRa17 101383.81346960185
Lbr17 netRa17 netL17 -1.0624564101529589e-11
Rbbr17 netL17 node_2 -103213.4992572819
Cbr17 netL17 node_2 -9.942242687654117e-22

* Branch 18
Rabr18 node_1 netRa18 77.93561859167578
Lbr18 netRa18 netL18 1.644920510865221e-13
Rbbr18 netL18 node_2 569.7960725068245
Cbr18 netL18 node_2 3.589026697541792e-18

* Branch 19
Rabr19 node_1 netRa19 6011440547681.191
Lbr19 netRa19 netL19 -0.004384023081428588
Rbbr19 netL19 node_2 -11478488297700.549
Cbr19 netL19 node_2 -6.329290218467077e-29

* Branch 20
Rabr20 node_1 netRa20 -6375093887.946673
Lbr20 netRa20 netL20 1.2039358398543554e-05
Rbbr20 netL20 node_2 45410180928.06233
Cbr20 netL20 node_2 4.048826186302198e-26

* Branch 21
Rabr21 node_1 netRa21 31475904.729200304
Lbr21 netRa21 netL21 -1.757306259310119e-07
Rbbr21 netL21 node_2 -1579821020.463824
Cbr21 netL21 node_2 -3.1623791291660385e-24

* Branch 22
Rabr22 node_1 netRa22 -25540230.639993984
Lbr22 netRa22 netL22 1.655655698443955e-07
Rbbr22 netL22 node_2 1685477180.896122
Cbr22 netL22 node_2 3.372849595481827e-24

* Branch 23
Rabr23 node_1 netRa23 -15999196.735114664
Lbr23 netRa23 netL23 -1.7164764581317053e-08
Rbbr23 netL23 node_2 51198305.21284598
Cbr23 netL23 node_2 -2.2681556580926354e-23

* Branch 24
Rabr24 node_1 netRa24 934.5330243417428
Lbr24 netRa24 netL24 2.647763378631919e-12
Rbbr24 netL24 node_2 -27794.63053163269
Cbr24 netL24 node_2 2.0229557828985536e-19

* Branch 25
Rd node_1 node_2 53018.07495038988

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 -6634.796098705327
Lbr0 netRa0 netL0 -6.939696432593943e-12
Rbbr0 netL0 node_3 33585.53095734019
Cbr0 netL0 node_3 -1.2350471144298714e-19

* Branch 1
Rabr1 node_1 netRa1 -3262219237326.67
Lbr1 netRa1 netL1 -0.0020812310649534955
Rbbr1 netL1 node_3 4994164444862.352
Cbr1 netL1 node_3 -1.2778056393006496e-28

* Branch 2
Rabr2 node_1 netRa2 14.161990423481035
Lbr2 netRa2 netL2 6.868351767830944e-13
Rbbr2 netL2 node_3 148878.8445162447
Cbr2 netL2 node_3 1.1105538694664266e-18

* Branch 3
Rabr3 node_1 netRa3 340428.481667969
Lbr3 netRa3 netL3 5.710793673448848e-09
Rbbr3 netL3 node_3 -565783727.942474
Cbr3 netL3 node_3 1.333996792026076e-22

* Branch 4
Rabr4 node_1 netRa4 -87601.15140212339
Lbr4 netRa4 netL4 -3.633250518561993e-10
Rbbr4 netL4 node_3 3027978.8964890605
Cbr4 netL4 node_3 -2.034243993616767e-21

* Branch 5
Rabr5 node_1 netRa5 75882.11170268759
Lbr5 netRa5 netL5 1.8595489773673843e-10
Rbbr5 netL5 node_3 -855580.9152158172
Cbr5 netL5 node_3 3.726185039250213e-21

* Branch 6
Rabr6 node_1 netRa6 250514813987.49377
Lbr6 netRa6 netL6 7.104358256397065e-05
Rbbr6 netL6 node_3 -277130288426.3605
Cbr6 netL6 node_3 1.0252002503944488e-27

* Branch 7
Rabr7 node_1 netRa7 -536.1932716823479
Lbr7 netRa7 netL7 -1.2188407337668296e-12
Rbbr7 netL7 node_3 43697.50246710902
Cbr7 netL7 node_3 -5.871451523112196e-19

* Branch 8
Rabr8 node_1 netRa8 207.8752967761388
Lbr8 netRa8 netL8 1.0590994755410786e-12
Rbbr8 netL8 node_3 -51590.03651740198
Cbr8 netL8 node_3 6.605955986567188e-19

* Branch 9
Rabr9 node_1 netRa9 9792.17583433229
Lbr9 netRa9 netL9 3.678169037470664e-11
Rbbr9 netL9 node_3 -321745.2882138047
Cbr9 netL9 node_3 1.7429775031273007e-20

* Branch 10
Rabr10 node_1 netRa10 4062225290825.1953
Lbr10 netRa10 netL10 0.0015601180736573928
Rbbr10 netL10 node_3 -4974371150645.984
Cbr10 netL10 node_3 7.72983027535332e-29

* Branch 11
Rabr11 node_1 netRa11 202918.10165148586
Lbr11 netRa11 netL11 1.3557678171487514e-10
Rbbr11 netL11 node_3 -346767.3235861877
Cbr11 netL11 node_3 2.002526899438682e-21

* Branch 12
Rabr12 node_1 netRa12 274158616.8117368
Lbr12 netRa12 netL12 1.2950359487924128e-08
Rbbr12 netL12 node_3 -275096752.1700587
Cbr12 netL12 node_3 1.721069660169454e-25

* Branch 13
Rabr13 node_1 netRa13 -191001.62403041363
Lbr13 netRa13 netL13 -1.3869767480656638e-10
Rbbr13 netL13 node_3 351498.19060441415
Cbr13 netL13 node_3 -2.1514060935447054e-21

* Branch 14
Rabr14 node_1 netRa14 -3.3071472458348716
Lbr14 netRa14 netL14 7.182399474762128e-13
Rbbr14 netL14 node_3 9859.534291596981
Cbr14 netL14 node_3 9.060750306146038e-19

* Branch 15
Rabr15 node_1 netRa15 -22797390066483.086
Lbr15 netRa15 netL15 -0.010018427719696202
Rbbr15 netL15 node_3 29693746813296.91
Cbr15 netL15 node_3 -1.4802319622723527e-29

* Branch 16
Rabr16 node_1 netRa16 -47.20004994712304
Lbr16 netRa16 netL16 2.4768444461059807e-13
Rbbr16 netL16 node_3 827.3402062891598
Cbr16 netL16 node_3 2.373199459669667e-18

* Branch 17
Rabr17 node_1 netRa17 133590.05438124863
Lbr17 netRa17 netL17 -1.0722531962117394e-11
Rbbr17 netL17 node_3 -135011.27530533753
Cbr17 netL17 node_3 -5.849916570666743e-22

* Branch 18
Rabr18 node_1 netRa18 57.81826898293501
Lbr18 netRa18 netL18 1.3024432706129608e-13
Rbbr18 netL18 node_3 425.52498072320515
Cbr18 netL18 node_3 4.52916029138509e-18

* Branch 19
Rabr19 node_1 netRa19 -63135470602141.69
Lbr19 netRa19 netL19 0.006050420050107373
Rbbr19 netL19 node_3 64130234874100.14
Cbr19 netL19 node_3 1.4935903268841845e-30

* Branch 20
Rabr20 node_1 netRa20 -5313750290.551541
Lbr20 netRa20 netL20 -5.444464855534572e-06
Rbbr20 netL20 node_3 15298192343.408133
Cbr20 netL20 node_3 -6.797653785017998e-26

* Branch 21
Rabr21 node_1 netRa21 107102034.47261105
Lbr21 netRa21 netL21 1.1593292356099775e-07
Rbbr21 netL21 node_3 -333578213.84611666
Cbr21 netL21 node_3 3.320623016036402e-24

* Branch 22
Rabr22 node_1 netRa22 -103781370.06359683
Lbr22 netRa22 netL22 -1.1259848740766349e-07
Rbbr22 netL22 node_3 324413198.0670477
Cbr22 netL22 node_3 -3.424801308073757e-24

* Branch 23
Rabr23 node_1 netRa23 -32503781.31893773
Lbr23 netRa23 netL23 -2.8946987143068606e-08
Rbbr23 netL23 node_3 81098482.64854234
Cbr23 netL23 node_3 -1.1722154704936155e-23

* Branch 24
Rabr24 node_1 netRa24 784.4465678714035
Lbr24 netRa24 netL24 2.121404130192113e-12
Rbbr24 netL24 node_3 -20444.96614673414
Cbr24 netL24 node_3 2.5124884096771903e-19

* Branch 25
Rd node_1 node_3 28067.38486012204

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 -11945.450488360362
Lbr0 netRa0 netL0 -8.289714149038187e-12
Rbbr0 netL0 node_4 22635.72643677847
Cbr0 netL0 node_4 -6.084999257433421e-20

* Branch 1
Rabr1 node_1 netRa1 -14226047150632.889
Lbr1 netRa1 netL1 0.008667394310024083
Rbbr1 netL1 node_4 21110414657936.41
Cbr1 netL1 node_4 2.8853102447493664e-29

* Branch 2
Rabr2 node_1 netRa2 15.932781675283815
Lbr2 netRa2 netL2 7.72676371225417e-13
Rbbr2 netL2 node_4 167515.0423400257
Cbr2 netL2 node_4 9.871758510142482e-19

* Branch 3
Rabr3 node_1 netRa3 -7841892.308916217
Lbr3 netRa3 netL3 2.4902385878599057e-08
Rbbr3 netL3 node_4 98269207.7519519
Cbr3 netL3 node_4 2.816786109708501e-23

* Branch 4
Rabr4 node_1 netRa4 56606.32234373995
Lbr4 netRa4 netL4 -9.123193683553871e-10
Rbbr4 netL4 node_4 -8569311.896998512
Cbr4 netL4 node_4 -8.287487213945387e-22

* Branch 5
Rabr5 node_1 netRa5 60351.72285527484
Lbr5 netRa5 netL5 3.796227602851541e-10
Rbbr5 netL5 node_4 -7791337.3743757475
Cbr5 netL5 node_4 1.9873615095577053e-21

* Branch 6
Rabr6 node_1 netRa6 457432329695.82104
Lbr6 netRa6 netL6 0.00030673748470997963
Rbbr6 netL6 node_4 -729840738932.0848
Cbr6 netL6 node_4 9.228027828465363e-28

* Branch 7
Rabr7 node_1 netRa7 -888.3153145427641
Lbr7 netRa7 netL7 -1.3722535892850259e-12
Rbbr7 netL7 node_4 8575.132374369614
Cbr7 netL7 node_4 -4.732883151987216e-19

* Branch 8
Rabr8 node_1 netRa8 201.97303872220652
Lbr8 netRa8 netL8 1.1866247438386573e-12
Rbbr8 netL8 node_4 -515981.95799123775
Cbr8 netL8 node_4 5.91755721141327e-19

* Branch 9
Rabr9 node_1 netRa9 18278.483067136236
Lbr9 netRa9 netL9 5.291348083721626e-11
Rbbr9 netL9 node_4 -329008.7539520334
Cbr9 netL9 node_4 1.180201376498e-20

* Branch 10
Rabr10 node_1 netRa10 19055941425765.32
Lbr10 netRa10 netL10 0.0062710265426241295
Rbbr10 netL10 node_4 -22197075872625.598
Cbr10 netL10 node_4 1.4840667705721482e-29

* Branch 11
Rabr11 node_1 netRa11 228099.3136086958
Lbr11 netRa11 netL11 2.838522526329282e-10
Rbbr11 netL11 node_4 -808737.3113985913
Cbr11 netL11 node_4 1.6553885871165548e-21

* Branch 12
Rabr12 node_1 netRa12 17502670.53603567
Lbr12 netRa12 netL12 6.364603268286836e-09
Rbbr12 netL12 node_4 -21107855.07986207
Cbr12 netL12 node_4 1.7539301365016966e-23

* Branch 13
Rabr13 node_1 netRa13 -194753.80008857857
Lbr13 netRa13 netL13 -3.043697353037252e-10
Rbbr13 netL13 node_4 990735.2008086717
Cbr13 netL13 node_4 -1.7250146268515765e-21

* Branch 14
Rabr14 node_1 netRa14 -7.373365164719973
Lbr14 netRa14 netL14 8.026985624789454e-13
Rbbr14 netL14 node_4 10589.519049980136
Cbr14 netL14 node_4 8.1044665093117635e-19

* Branch 15
Rabr15 node_1 netRa15 -1573729302101.4668
Lbr15 netRa15 netL15 -0.012681441825264131
Rbbr15 netL15 node_4 162159902745005.72
Cbr15 netL15 node_4 -4.98621119199178e-29

* Branch 16
Rabr16 node_1 netRa16 -35.59668198727279
Lbr16 netRa16 netL16 2.7082609875927304e-13
Rbbr16 netL16 node_4 1000.665794975588
Cbr16 netL16 node_4 2.219848409020725e-18

* Branch 17
Rabr17 node_1 netRa17 96341.78273805525
Lbr17 netRa17 netL17 -9.817449264898737e-12
Rbbr17 netL17 node_4 -97986.7407663091
Cbr17 netL17 node_4 -1.0189299124116377e-21

* Branch 18
Rabr18 node_1 netRa18 69.51038183977009
Lbr18 netRa18 netL18 1.4791089852135747e-13
Rbbr18 netL18 node_4 508.3810309337321
Cbr18 netL18 node_4 3.9911921667493296e-18

* Branch 19
Rabr19 node_1 netRa19 2933898327951.681
Lbr19 netRa19 netL19 -0.0027730268790541195
Rbbr19 netL19 node_4 -7410621753774.555
Cbr19 netL19 node_4 -1.269144899424929e-28

* Branch 20
Rabr20 node_1 netRa20 17476239241.344147
Lbr20 netRa20 netL20 9.954083647943965e-06
Rbbr20 netL20 node_4 -27557040999.541203
Cbr20 netL20 node_4 2.083971438041229e-26

* Branch 21
Rabr21 node_1 netRa21 -223775974.10526636
Lbr21 netRa21 netL21 -1.7011151912398515e-07
Rbbr21 netL21 node_4 455545779.59205914
Cbr21 netL21 node_4 -1.6958702304283235e-24

* Branch 22
Rabr22 node_1 netRa22 207917843.75988835
Lbr22 netRa22 netL22 1.6150299000629666e-07
Rbbr22 netL22 node_4 -432945072.1508967
Cbr22 netL22 node_4 1.824819828527278e-24

* Branch 23
Rabr23 node_1 netRa23 -17728319.410902724
Lbr23 netRa23 netL23 -1.651268469678644e-08
Rbbr23 netL23 node_4 46810703.10384697
Cbr23 netL23 node_4 -2.1305992787971099e-23

* Branch 24
Rabr24 node_1 netRa24 844.0323713392289
Lbr24 netRa24 netL24 2.381462726625111e-12
Rbbr24 netL24 node_4 -24805.178893130374
Cbr24 netL24 node_4 2.2482278568179794e-19

* Branch 25
Rd node_1 node_4 44392.730014294175

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 -58958.67280722766
Lbr0 netRa0 netL0 1.6866021586814657e-11
Rbbr0 netL0 0 62708.867363470265
Cbr0 netL0 0 3.787196124189996e-21

* Branch 1
Rabr1 node_2 netRa1 483262372871.12787
Lbr1 netRa1 netL1 -0.0004079616543122876
Rbbr1 netL1 0 -932196418702.4386
Cbr1 netL1 0 -9.052521356657034e-28

* Branch 2
Rabr2 node_2 netRa2 -422287052.4156599
Lbr2 netRa2 netL2 -2.788030451573498e-07
Rbbr2 netL2 0 667956352.1280181
Cbr2 netL2 0 -1.0061347295226722e-24

* Branch 3
Rabr3 node_2 netRa3 1.7267074189558724
Lbr3 netRa3 netL3 1.0874517038766501e-13
Rbbr3 netL3 0 4678.116696041926
Cbr3 netL3 0 7.012339555589282e-18

* Branch 4
Rabr4 node_2 netRa4 11902.474111870413
Lbr4 netRa4 netL4 1.0821479399659834e-10
Rbbr4 netL4 0 -4565057.043699441
Cbr4 netL4 0 7.014999617587113e-21

* Branch 5
Rabr5 node_2 netRa5 -2104.5282692831192
Lbr5 netRa5 netL5 -4.037946576819045e-11
Rbbr5 netL5 0 -1254057.7595582416
Cbr5 netL5 0 -1.886139900219508e-20

* Branch 6
Rabr6 node_2 netRa6 4776504803.339461
Lbr6 netRa6 netL6 4.658962071809921e-05
Rbbr6 netL6 0 -644554954529.4689
Cbr6 netL6 0 1.6157115152617092e-26

* Branch 7
Rabr7 node_2 netRa7 103.2355998865989
Lbr7 netRa7 netL7 9.159681571247835e-14
Rbbr7 netL7 0 -277.3429445587365
Cbr7 netL7 0 4.965626378463986e-18

* Branch 8
Rabr8 node_2 netRa8 33160.62781392425
Lbr8 netRa8 netL8 -7.18706234765153e-12
Rbbr8 netL8 0 -35300.65310033588
Cbr8 netL8 0 -5.9253041624781095e-21

* Branch 9
Rabr9 node_2 netRa9 -221724.29437387356
Lbr9 netRa9 netL9 4.3793447443159096e-11
Rbbr9 netL9 0 234582.57500899278
Cbr9 netL9 0 8.2760738043667225e-22

* Branch 10
Rabr10 node_2 netRa10 -1852601380.6280322
Lbr10 netRa10 netL10 0.00019229036799383909
Rbbr10 netL10 0 22991191939484.047
Cbr10 netL10 0 3.419863674086599e-27

* Branch 11
Rabr11 node_2 netRa11 -6802.001957867898
Lbr11 netRa11 netL11 2.5867616935548865e-12
Rbbr11 netL11 0 8273.391261385439
Cbr11 netL11 0 4.499683203345428e-20

* Branch 12
Rabr12 node_2 netRa12 -7340.11556267859
Lbr12 netRa12 netL12 -2.2873681099531273e-11
Rbbr12 netL12 0 136000.24935387785
Cbr12 netL12 0 -2.7031395274307078e-20

* Branch 13
Rabr13 node_2 netRa13 14.17319431346285
Lbr13 netRa13 netL13 1.0697617235479458e-13
Rbbr13 netL13 0 -2119.4179968613416
Cbr13 netL13 0 6.068031879611384e-18

* Branch 14
Rabr14 node_2 netRa14 806515.5113376738
Lbr14 netRa14 netL14 5.794794992569439e-11
Rbbr14 netL14 0 -812960.8573489776
Cbr14 netL14 0 8.906722922108838e-23

* Branch 15
Rabr15 node_2 netRa15 -621033816500.0723
Lbr15 netRa15 netL15 -0.0009952150480061065
Rbbr15 netL15 0 3120441084171.458
Cbr15 netL15 0 -5.139001395135239e-28

* Branch 16
Rabr16 node_2 netRa16 -1.149478160468813
Lbr16 netRa16 netL16 1.2392874655366067e-14
Rbbr16 netL16 0 49.46210845256001
Cbr16 netL16 0 4.9131550552683606e-17

* Branch 17
Rabr17 node_2 netRa17 -619301.8259594775
Lbr17 netRa17 netL17 -2.5983995279577763e-11
Rbbr17 netL17 0 621147.0981943515
Cbr17 netL17 0 -6.812641353381883e-23

* Branch 18
Rabr18 node_2 netRa18 170.82091460801874
Lbr18 netRa18 netL18 6.208213577937128e-13
Rbbr18 netL18 0 1567.626442863059
Cbr18 netL18 0 9.276800660131313e-19

* Branch 19
Rabr19 node_2 netRa19 -59660687556.48583
Lbr19 netRa19 netL19 -0.00024388830954794632
Rbbr19 netL19 0 1808408354263.9326
Cbr19 netL19 0 -2.3099327192313463e-27

* Branch 20
Rabr20 node_2 netRa20 0.7181994414489832
Lbr20 netRa20 netL20 1.1160903775932268e-13
Rbbr20 netL20 0 24780.826340395994
Cbr20 netL20 0 5.080936639192407e-18

* Branch 21
Rabr21 node_2 netRa21 -922689.6836096117
Lbr21 netRa21 netL21 2.1333795938542447e-09
Rbbr21 netL21 0 9218217.635377783
Cbr21 netL21 0 2.391830765106547e-22

* Branch 22
Rabr22 node_2 netRa22 913803.4130019225
Lbr22 netRa22 netL22 -2.24135626166889e-09
Rbbr22 netL22 0 -10120520.596333176
Cbr22 netL22 0 -2.3013853534339357e-22

* Branch 23
Rabr23 node_2 netRa23 -9409184.354054417
Lbr23 netRa23 netL23 1.5714221096297626e-08
Rbbr23 netL23 0 50843435.74668397
Cbr23 netL23 0 2.936745929425943e-23

* Branch 24
Rabr24 node_2 netRa24 -6367761.957930266
Lbr24 netRa24 netL24 -3.4385466901752334e-10
Rbbr24 netL24 0 6401581.686395151
Cbr24 netL24 0 -8.515826033768675e-24

* Branch 25
Rd node_2 0 10396.85643184949

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 -11154.090247487133
Lbr0 netRa0 netL0 -6.6170838670767985e-12
Rbbr0 netL0 node_3 17536.58404108119
Cbr0 netL0 node_3 -5.874682052516619e-20

* Branch 1
Rabr1 node_2 netRa1 79697706469081.73
Lbr1 netRa1 netL1 -0.014271657293607585
Rbbr1 netL1 node_3 -83030093158039.72
Cbr1 netL1 node_3 -2.1565485887412924e-30

* Branch 2
Rabr2 node_2 netRa2 12.392423846040678
Lbr2 netRa2 netL2 6.00964957795249e-13
Rbbr2 netL2 node_3 130301.71382004907
Cbr2 netL2 node_3 1.2692378135205107e-18

* Branch 3
Rabr3 node_2 netRa3 -45993404.53721265
Lbr3 netRa3 netL3 -3.790362554869288e-08
Rbbr3 netL3 node_3 88599514.79795651
Cbr3 netL3 node_3 -9.671023447004833e-24

* Branch 4
Rabr4 node_2 netRa4 1850095.018152275
Lbr4 netRa4 netL4 -1.886748236962749e-09
Rbbr4 netL4 node_3 -4190182.6796810185
Cbr4 netL4 node_3 -2.252855414294133e-22

* Branch 5
Rabr5 node_2 netRa5 -111126.50790713885
Lbr5 netRa5 netL5 4.998541823819364e-10
Rbbr5 netL5 node_3 2186851.1210505585
Cbr5 netL5 node_3 1.443821308762533e-21

* Branch 6
Rabr6 node_2 netRa6 -3688751174737.8174
Lbr6 netRa6 netL6 -0.00041345688051303296
Rbbr6 netL6 node_3 3749903680636.43
Cbr6 netL6 node_3 -2.9912124577758636e-29

* Branch 7
Rabr7 node_2 netRa7 -793.7399512004272
Lbr7 netRa7 netL7 -1.0654065259326579e-12
Rbbr7 netL7 node_3 5067.579979914191
Cbr7 netL7 node_3 -5.735307973225675e-19

* Branch 8
Rabr8 node_2 netRa8 145.36796903970182
Lbr8 netRa8 netL8 9.212620632815338e-13
Rbbr8 netL8 node_3 143329.8109089029
Cbr8 netL8 node_3 7.632783708066163e-19

* Branch 9
Rabr9 node_2 netRa9 19306.116986679783
Lbr9 netRa9 netL9 4.733632787392568e-11
Rbbr9 netL9 node_3 -243061.85170177225
Cbr9 netL9 node_3 1.28590577508109e-20

* Branch 10
Rabr10 node_2 netRa10 -51887982740952.66
Lbr10 netRa10 netL10 -0.01188691972967154
Rbbr10 netL10 node_3 56031579506568.77
Cbr10 netL10 node_3 -4.091443998775763e-30

* Branch 11
Rabr11 node_2 netRa11 -80179.57300048778
Lbr11 netRa11 netL11 4.1738950281580577e-10
Rbbr11 netL11 node_3 2644179.31192726
Cbr11 netL11 node_3 1.520477085765846e-21

* Branch 12
Rabr12 node_2 netRa12 -1885440.6781900185
Lbr12 netRa12 netL12 4.767492957309715e-09
Rbbr12 netL12 node_3 18300897.176019784
Cbr12 netL12 node_3 1.2296761633458543e-22

* Branch 13
Rabr13 node_2 netRa13 301854.1387859764
Lbr13 netRa13 netL13 -4.923456687081461e-10
Rbbr13 netL13 node_3 -1429979.3140262903
Cbr13 netL13 node_3 -1.0471438265759541e-21

* Branch 14
Rabr14 node_2 netRa14 -7.1415166742167004
Lbr14 netRa14 netL14 6.224093311946608e-13
Rbbr14 netL14 node_3 8054.459128998648
Cbr14 netL14 node_3 1.0450043114948852e-18

* Branch 15
Rabr15 node_2 netRa15 -2032787205529.2268
Lbr15 netRa15 netL15 -0.004514867978153152
Rbbr15 netL15 node_3 17751962453776.754
Cbr15 netL15 node_3 -1.2523132001841755e-28

* Branch 16
Rabr16 node_2 netRa16 -21.740468355617708
Lbr16 netRa16 netL16 2.0776934952530295e-13
Rbbr16 netL16 node_3 808.9766510121863
Cbr16 netL16 node_3 2.9196584539440145e-18

* Branch 17
Rabr17 node_2 netRa17 61904.2479287565
Lbr17 netRa17 netL17 -6.994808793155253e-12
Rbbr17 netL17 node_3 -63200.97487130536
Cbr17 netL17 node_3 -1.747850883698925e-21

* Branch 18
Rabr18 node_2 netRa18 55.75987035754181
Lbr18 netRa18 netL18 1.1554733277980816e-13
Rbbr18 netL18 node_3 407.55396463856493
Cbr18 netL18 node_3 5.109473274843689e-18

* Branch 19
Rabr19 node_2 netRa19 2017854724835.7644
Lbr19 netRa19 netL19 -0.0015281271725366397
Rbbr19 netL19 node_3 -3996424670395.692
Cbr19 netL19 node_3 -1.88746952823454e-28

* Branch 20
Rabr20 node_2 netRa20 -1778340057.65212
Lbr20 netRa20 netL20 3.6258374143794717e-06
Rbbr20 netL20 node_3 14443878389.976671
Cbr20 netL20 node_3 1.371393418218053e-25

* Branch 21
Rabr21 node_2 netRa21 3760627.8377702297
Lbr21 netRa21 netL21 -6.264243198073057e-08
Rbbr21 netL21 node_3 -1366328042.2805824
Cbr21 netL21 node_3 -9.026843590292712e-24

* Branch 22
Rabr22 node_2 netRa22 -1897827.4140499306
Lbr22 netRa22 netL22 5.972404970862633e-08
Rbbr22 netL22 node_3 1973556777.760089
Cbr22 netL22 node_3 9.484866209135246e-24

* Branch 23
Rabr23 node_2 netRa23 -10043579.481683327
Lbr23 netRa23 netL23 -1.026871385697742e-08
Rbbr23 netL23 node_3 30033846.352331564
Cbr23 netL23 node_3 -3.670508326030274e-23

* Branch 24
Rabr24 node_2 netRa24 642.2389850601187
Lbr24 netRa24 netL24 1.8507386165324577e-12
Rbbr24 netL24 node_3 -20065.029703324784
Cbr24 netL24 node_3 2.8989826668238836e-19

* Branch 25
Rd node_2 node_3 42800.94281295713

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 -8468.143568436552
Lbr0 netRa0 netL0 -5.538862320696702e-12
Rbbr0 netL0 node_4 14839.855330539074
Cbr0 netL0 node_4 -8.279640681569968e-20

* Branch 1
Rabr1 node_2 netRa1 11735175958686.732
Lbr1 netRa1 netL1 -0.003534695975615416
Rbbr1 netL1 node_4 -13123349822453.537
Cbr1 netL1 node_4 -2.2948847623254334e-29

* Branch 2
Rabr2 node_2 netRa2 10.621842152527817
Lbr2 netRa2 netL2 5.151150536835056e-13
Rbbr2 netL2 node_4 111677.5744563414
Cbr2 netL2 node_4 1.4807710398158708e-18

* Branch 3
Rabr3 node_2 netRa3 -131860916.1519252
Lbr3 netRa3 netL3 7.786703232182521e-08
Rbbr3 netL3 node_4 190575811.28157562
Cbr3 netL3 node_4 3.01605693074859e-24

* Branch 4
Rabr4 node_2 netRa4 188166.45641476594
Lbr4 netRa4 netL4 -9.00156497252029e-10
Rbbr4 netL4 node_4 -4297571.304918377
Cbr4 netL4 node_4 -8.085109773868145e-22

* Branch 5
Rabr5 node_2 netRa5 27943.211726854435
Lbr5 netRa5 netL5 3.235385091319109e-10
Rbbr5 netL5 node_4 52971863.20836574
Cbr5 netL5 node_4 2.3513068795385113e-21

* Branch 6
Rabr6 node_2 netRa6 -1004329918720.1863
Lbr6 netRa6 netL6 0.00033603086700960606
Rbbr6 netL6 node_4 1152259549803.4993
Cbr6 netL6 node_4 2.897403793880415e-28

* Branch 7
Rabr7 node_2 netRa7 -625.2020805508326
Lbr7 netRa7 netL7 -9.09613135223438e-13
Rbbr7 netL7 node_4 5009.048518704031
Cbr7 netL7 node_4 -6.971043886584865e-19

* Branch 8
Rabr8 node_2 netRa8 129.95758292932715
Lbr8 netRa8 netL8 7.91049972478329e-13
Rbbr8 netL8 node_4 425135.1372300574
Cbr8 netL8 node_4 8.882898792476969e-19

* Branch 9
Rabr9 node_2 netRa9 14504.09475339277
Lbr9 netRa9 netL9 3.772455239274821e-11
Rbbr9 netL9 node_4 -206881.3932509571
Cbr9 netL9 node_4 1.629876253816502e-20

* Branch 10
Rabr10 node_2 netRa10 638513636233.149
Lbr10 netRa10 netL10 0.004860731248356195
Rbbr10 netL10 node_4 -58255304382816.56
Cbr10 netL10 node_4 1.338176196039368e-28

* Branch 11
Rabr11 node_2 netRa11 131545.7427643005
Lbr11 netRa11 netL11 2.6150481968966974e-10
Rbbr11 netL11 node_4 -1026622.66815547
Cbr11 netL11 node_4 2.182047211188814e-21

* Branch 12
Rabr12 node_2 netRa12 5804195.91450747
Lbr12 netRa12 netL12 4.704567680841986e-09
Rbbr12 netL12 node_4 -11879319.190305268
Cbr12 netL12 node_4 7.104672341830388e-23

* Branch 13
Rabr13 node_2 netRa13 -77870.87775450741
Lbr13 netRa13 netL13 -2.9062793546907304e-10
Rbbr13 netL13 node_4 2163738.3960889704
Cbr13 netL13 node_4 -2.1676718358294097e-21

* Branch 14
Rabr14 node_2 netRa14 -5.6227074606186385
Lbr14 netRa14 netL14 5.343828995113755e-13
Rbbr14 netL14 node_4 6970.637128020473
Cbr14 netL14 node_4 1.2172405444559915e-18

* Branch 15
Rabr15 node_2 netRa15 -344850520288.85675
Lbr15 netRa15 netL15 -0.003492483992487768
Rbbr15 netL15 node_4 55976072605965.73
Cbr15 netL15 node_4 -1.81700608033482e-28

* Branch 16
Rabr16 node_2 netRa16 -21.45891415332748
Lbr16 netRa16 netL16 1.7926017541628075e-13
Rbbr16 netL16 node_4 677.3277841107939
Cbr16 netL16 node_4 3.367276509020653e-18

* Branch 17
Rabr17 node_2 netRa17 58089.939542264576
Lbr17 netRa17 netL17 -6.245633446884328e-12
Rbbr17 netL17 node_4 -59192.85096254367
Cbr17 netL17 node_4 -1.7776667626678824e-21

* Branch 18
Rabr18 node_2 netRa18 46.96266333084864
Lbr18 netRa18 netL18 9.877063970117867e-14
Rbbr18 netL18 node_4 343.3111304298015
Cbr18 netL18 node_4 5.9772242535679795e-18

* Branch 19
Rabr19 node_2 netRa19 485650485570.2905
Lbr19 netRa19 netL19 -0.0009417072525182457
Rbbr19 netL19 node_4 -3588515372325.9146
Cbr19 netL19 node_4 -5.349236623043398e-28

* Branch 20
Rabr20 node_2 netRa20 286208451.73444873
Lbr20 netRa20 netL20 4.0034360969716715e-06
Rbbr20 netL20 node_4 -123898935963.43802
Cbr20 netL20 node_4 1.413166287390174e-25

* Branch 21
Rabr21 node_2 netRa21 -18336440.044578977
Lbr21 netRa21 netL21 -7.188954840119923e-08
Rbbr21 netL21 node_4 560106104.2540636
Cbr21 netL21 node_4 -7.629219900749758e-24

* Branch 22
Rabr22 node_2 netRa22 18456598.882929757
Lbr22 netRa22 netL22 6.85643574204718e-08
Rbbr22 netL22 node_4 -506943140.2142833
Cbr22 netL22 node_4 7.968805555995658e-24

* Branch 23
Rabr23 node_2 netRa23 -9755748.840283042
Lbr23 netRa23 netL23 -9.76100863499373e-09
Rbbr23 netL23 node_4 28320001.94202698
Cbr23 netL23 node_4 -3.8029808061357517e-23

* Branch 24
Rabr24 node_2 netRa24 557.0226820662363
Lbr24 netRa24 netL24 1.5873513167266032e-12
Rbbr24 netL24 node_4 -16846.541166694627
Cbr24 netL24 node_4 3.376317847947056e-19

* Branch 25
Rd node_2 node_4 32154.546116119975

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 -869.022416970003
Lbr0 netRa0 netL0 -2.2011834138500776e-12
Rbbr0 netL0 0 -5567.479987528269
Cbr0 netL0 0 -5.609713030260166e-19

* Branch 1
Rabr1 node_3 netRa1 -7733101796746210.0
Lbr1 netRa1 netL1 -0.08586888799527581
Rbbr1 netL1 0 7734345183559135.0
Cbr1 netL1 0 -1.4356899413415009e-33

* Branch 2
Rabr2 node_3 netRa2 284600834.35665107
Lbr2 netRa2 netL2 4.5410479261362565e-07
Rbbr2 netL2 0 -1276823413.3674994
Cbr2 netL2 0 1.3051878785390611e-24

* Branch 3
Rabr3 node_3 netRa3 -10169685.573108891
Lbr3 netRa3 netL3 -1.4724747016982926e-08
Rbbr3 netL3 0 40151188.86791177
Cbr3 netL3 0 -3.865625696387294e-23

* Branch 4
Rabr4 node_3 netRa4 81613.99155026242
Lbr4 netRa4 netL4 1.1166523789386122e-10
Rbbr4 netL4 0 -306593.78764344426
Cbr4 netL4 0 5.001615200008138e-21

* Branch 5
Rabr5 node_3 netRa5 4.924828553950692
Lbr5 netRa5 netL5 1.2254133330437985e-13
Rbbr5 netL5 0 2968.2491424067707
Cbr5 netL5 0 6.215035729728377e-18

* Branch 6
Rabr6 node_3 netRa6 196303866604.36008
Lbr6 netRa6 netL6 -0.00010985782585172186
Rbbr6 netL6 0 -277078119116.9404
Cbr6 netL6 0 -2.0124405331824944e-27

* Branch 7
Rabr7 node_3 netRa7 625.6723560866168
Lbr7 netRa7 netL7 -5.114032623213337e-13
Rbbr7 netL7 0 -1060.202162843124
Cbr7 netL7 0 -5.80659904013874e-19

* Branch 8
Rabr8 node_3 netRa8 14240.699170346921
Lbr8 netRa8 netL8 9.15713355159246e-12
Rbbr8 netL8 0 -23630.942635276664
Cbr8 netL8 0 3.0483312272197785e-20

* Branch 9
Rabr9 node_3 netRa9 -6042.6301160432395
Lbr9 netRa9 netL9 -2.4449958519235648e-11
Rbbr9 netL9 0 238256.44646003356
Cbr9 netL9 0 -2.6357948660097818e-20

* Branch 10
Rabr10 node_3 netRa10 715709408920.3063
Lbr10 netRa10 netL10 -0.0005560714403749601
Rbbr10 netL10 0 -1371075221774.2986
Cbr10 netL10 0 -5.653185429630544e-28

* Branch 11
Rabr11 node_3 netRa11 -616.0142709793517
Lbr11 netRa11 netL11 -2.427972249572087e-12
Rbbr11 netL11 0 19439.540630260824
Cbr11 netL11 0 -2.610150794205552e-19

* Branch 12
Rabr12 node_3 netRa12 2353957.704292421
Lbr12 netRa12 netL12 2.873233224137792e-10
Rbbr12 netL12 0 -2407938.8306303467
Cbr12 netL12 0 5.0994794173101837e-23

* Branch 13
Rabr13 node_3 netRa13 2.8389726416916163
Lbr13 netRa13 netL13 1.1173666595589631e-13
Rbbr13 netL13 0 5827.648028540405
Cbr13 netL13 0 5.851466612458688e-18

* Branch 14
Rabr14 node_3 netRa14 654.1759018631572
Lbr14 netRa14 netL14 9.951765214932681e-12
Rbbr14 netL14 0 366826.54189450626
Cbr14 netL14 0 6.553195128982993e-20

* Branch 15
Rabr15 node_3 netRa15 -2531573941253.036
Lbr15 netRa15 netL15 -0.001766131410448303
Rbbr15 netL15 0 4461800696265.588
Cbr15 netL15 0 -1.5640469234505952e-28

* Branch 16
Rabr16 node_3 netRa16 0.46570550483583245
Lbr16 netRa16 netL16 1.6405640344648273e-14
Rbbr16 netL16 0 90.17351961274686
Cbr16 netL16 0 3.8193411040435643e-17

* Branch 17
Rabr17 node_3 netRa17 -3127.986233446666
Lbr17 netRa17 netL17 -1.8245174356515265e-12
Rbbr17 netL17 0 5153.22493396507
Cbr17 netL17 0 -1.2835257000315088e-19

* Branch 18
Rabr18 node_3 netRa18 151.61995666978927
Lbr18 netRa18 netL18 1.579688417803425e-13
Rbbr18 netL18 0 101894.7770315836
Cbr18 netL18 0 3.2924578851089378e-18

* Branch 19
Rabr19 node_3 netRa19 201584810123.1523
Lbr19 netRa19 netL19 0.0002420900746719508
Rbbr19 netL19 0 -703782779369.5698
Cbr19 netL19 0 1.717192576895445e-27

* Branch 20
Rabr20 node_3 netRa20 111211031.73560193
Lbr20 netRa20 netL20 -2.3103759678521023e-07
Rbbr20 netL20 0 -933085111.5541688
Cbr20 netL20 0 -2.1618816841464017e-24

* Branch 21
Rabr21 node_3 netRa21 2.234804261947914
Lbr21 netRa21 netL21 1.240349442565143e-13
Rbbr21 netL21 0 72230.63056830452
Cbr21 netL21 0 4.571628080768439e-18

* Branch 22
Rabr22 node_3 netRa22 -102928.72386251447
Lbr22 netRa22 netL22 2.0755933511464952e-10
Rbbr22 netL22 0 810215.3280252448
Cbr22 netL22 0 2.3847946840402532e-21

* Branch 23
Rabr23 node_3 netRa23 -246814.34625500656
Lbr23 netRa23 netL23 -1.836243278171447e-09
Rbbr23 netL23 0 51349487.76378943
Cbr23 netL23 0 -3.0691061849758366e-22

* Branch 24
Rabr24 node_3 netRa24 -87416.31844811312
Lbr24 netRa24 netL24 -2.6555247690659926e-11
Rbbr24 netL24 0 102788.22005533554
Cbr24 netL24 0 -3.1214240743248183e-21

* Branch 25
Rd node_3 0 3864.9770257720816

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 -14012.446739293115
Lbr0 netRa0 netL0 -9.986246008083463e-12
Rbbr0 netL0 node_4 27598.3037618555
Cbr0 netL0 node_4 -5.2651166119618906e-20

* Branch 1
Rabr1 node_3 netRa1 -160712084947663.5
Lbr1 netRa1 netL1 0.034239518815489284
Rbbr1 netL1 node_4 170223666868464.22
Cbr1 netL1 node_4 1.2514656929077265e-30

* Branch 2
Rabr2 node_3 netRa2 19.47318170218321
Lbr2 netRa2 netL2 9.443820693982653e-13
Rbbr2 netL2 node_4 204732.87177569797
Cbr2 netL2 node_4 8.076894733265907e-19

* Branch 3
Rabr3 node_3 netRa3 -7449706.4629991725
Lbr3 netRa3 netL3 3.19680192693419e-08
Rbbr3 netL3 node_4 157549243.85625398
Cbr3 netL3 node_4 2.271746920824238e-23

* Branch 4
Rabr4 node_3 netRa4 481.39299892555357
Lbr4 netRa4 netL4 -1.161950332008496e-09
Rbbr4 netL4 node_4 -19281979.036837984
Cbr4 netL4 node_4 -6.55012663628891e-22

* Branch 5
Rabr5 node_3 netRa5 100101.55657078506
Lbr5 netRa5 netL5 4.813175799232353e-10
Rbbr5 netL5 node_4 -5673651.646822453
Cbr5 netL5 node_4 1.5518286902368602e-21

* Branch 6
Rabr6 node_3 netRa6 566278175273.1096
Lbr6 netRa6 netL6 0.00027671418084916063
Rbbr6 netL6 node_4 -745145592130.1792
Cbr6 netL6 node_4 6.5787293708703605e-28

* Branch 7
Rabr7 node_3 netRa7 -1073.0639783751917
Lbr7 netRa7 netL7 -1.6692063755945595e-12
Rbbr7 netL7 node_4 10596.514726074714
Cbr7 netL7 node_4 -3.9009977946787877e-19

* Branch 8
Rabr8 node_3 netRa8 246.0669742215961
Lbr8 netRa8 netL8 1.4517142951192975e-12
Rbbr8 netL8 node_4 -804981.6857879492
Cbr8 netL8 node_4 4.837399637032149e-19

* Branch 9
Rabr9 node_3 netRa9 24926.119163141226
Lbr9 netRa9 netL9 6.592791233555367e-11
Rbbr9 netL9 node_4 -368533.21735480486
Cbr9 netL9 node_4 9.351095730789318e-21

* Branch 10
Rabr10 node_3 netRa10 12606632404330.527
Lbr10 netRa10 netL10 -0.004510047411984129
Rbbr10 netL10 node_4 -15057291602676.781
Cbr10 netL10 node_4 -2.3733198555212477e-29

* Branch 11
Rabr11 node_3 netRa11 415897.0213784191
Lbr11 netRa11 netL11 4.6146317894539495e-10
Rbbr11 netL11 node_4 -1250690.6612042708
Cbr11 netL11 node_4 9.466435920362142e-22

* Branch 12
Rabr12 node_3 netRa12 51482217.27971351
Lbr12 netRa12 netL12 1.4745022162329523e-08
Rbbr12 netL12 node_4 -58035468.09291971
Cbr12 netL12 node_4 5.005161552772594e-24

* Branch 13
Rabr13 node_3 netRa13 -351553.7903812062
Lbr13 netRa13 netL13 -5.079471051869302e-10
Rbbr13 netL13 node_4 1571035.0987420655
Cbr13 netL13 node_4 -9.98664686076068e-22

* Branch 14
Rabr14 node_3 netRa14 -9.744176774410658
Lbr14 netRa14 netL14 9.807976837811233e-13
Rbbr14 netL14 node_4 12857.19839578867
Cbr14 netL14 node_4 6.632400123505542e-19

* Branch 15
Rabr15 node_3 netRa15 -5804119758742.564
Lbr15 netRa15 netL15 -0.00927633866392683
Rbbr15 netL15 node_4 29038679767213.766
Cbr15 netL15 node_4 -5.507514106834677e-29

* Branch 16
Rabr16 node_3 netRa16 -43.30148838957103
Lbr16 netRa16 netL16 3.308211783820955e-13
Rbbr16 netL16 node_4 1223.5915081396547
Cbr16 netL16 node_4 1.8176214811783186e-18

* Branch 17
Rabr17 node_3 netRa17 116370.3180812909
Lbr17 netRa17 netL17 -1.1938026938665386e-11
Rbbr17 netL17 node_4 -118383.74601986766
Cbr17 netL17 node_4 -8.489203148516463e-22

* Branch 18
Rabr18 node_3 netRa18 84.73691033952494
Lbr18 netRa18 netL18 1.8072663311420623e-13
Rbbr18 netL18 node_4 619.8226896758126
Cbr18 netL18 node_4 3.2664349884428396e-18

* Branch 19
Rabr19 node_3 netRa19 5763619462564.384
Lbr19 netRa19 netL19 -0.0038348156556686597
Rbbr19 netL19 node_4 -10128016353395.596
Cbr19 netL19 node_4 -6.54658819035995e-29

* Branch 20
Rabr20 node_3 netRa20 2546239570.5561495
Lbr20 netRa20 netL20 7.000489084523928e-06
Rbbr20 netL20 node_4 -37884251915.258286
Cbr20 netL20 node_4 7.555889116460476e-26

* Branch 21
Rabr21 node_3 netRa21 -81841789.42932498
Lbr21 netRa21 netL21 -1.377692636371145e-07
Rbbr21 netL21 node_4 505868607.8059663
Cbr21 netL21 node_4 -3.4498861975118595e-24

* Branch 22
Rabr22 node_3 netRa22 80451736.08155847
Lbr22 netRa22 netL22 1.3228127654707586e-07
Rbbr22 netL22 node_4 -478193569.81396437
Cbr22 netL22 node_4 3.5653112582786944e-24

* Branch 23
Rabr23 node_3 netRa23 -21555850.12735926
Lbr23 netRa23 netL23 -1.9597527026593294e-08
Rbbr23 netL23 node_4 55188806.49513145
Cbr23 netL23 node_4 -1.7609515130518577e-23

* Branch 24
Rabr24 node_3 netRa24 1029.245461575668
Lbr24 netRa24 netL24 2.908977931697794e-12
Rbbr24 netL24 node_4 -30396.38809370876
Cbr24 netL24 node_4 1.840849004375475e-19

* Branch 25
Rd node_3 node_4 52605.093967580106

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 13138.835467508801
Lbr0 netRa0 netL0 -5.1071417176360886e-12
Rbbr0 netL0 0 -14593.257305911227
Cbr0 netL0 0 -2.0843269473730402e-20

* Branch 1
Rabr1 node_4 netRa1 8092374955850.347
Lbr1 netRa1 netL1 0.00488443775580368
Rbbr1 netL1 0 -11937879766193.309
Cbr1 netL1 0 5.057377464009484e-29

* Branch 2
Rabr2 node_4 netRa2 -232938280.01875106
Lbr2 netRa2 netL2 2.62586010644643e-07
Rbbr2 netL2 0 609718653.6066707
Cbr2 netL2 0 1.7948908958833307e-24

* Branch 3
Rabr3 node_4 netRa3 4775791.415677953
Lbr3 netRa3 netL3 -6.131725047595037e-09
Rbbr3 netL3 0 -14523355.636547836
Cbr3 netL3 0 -8.343708181747777e-23

* Branch 4
Rabr4 node_4 netRa4 4.0711739182797695
Lbr4 netRa4 netL4 1.198913418250038e-13
Rbbr4 netL4 0 3511.605644685727
Cbr4 netL4 0 6.355701464115726e-18

* Branch 5
Rabr5 node_4 netRa5 -5318.250944034199
Lbr5 netRa5 netL5 1.922198913604802e-11
Rbbr5 netL5 0 73447.62262272919
Cbr5 netL5 0 3.6691424517850693e-20

* Branch 6
Rabr6 node_4 netRa6 1340802469017.8376
Lbr6 netRa6 netL6 0.0002899820510064472
Rbbr6 netL6 0 -1423616709669.1372
Cbr6 netL6 0 1.5213325901781812e-28

* Branch 7
Rabr7 node_4 netRa7 3318.8846834090727
Lbr7 netRa7 netL7 -1.0397922586828402e-12
Rbbr7 netL7 0 -3718.3296720828007
Cbr7 netL7 0 -7.485433397077895e-20

* Branch 8
Rabr8 node_4 netRa8 3762.395835034609
Lbr8 netRa8 netL8 3.783351509185602e-12
Rbbr8 netL8 0 -10270.702620118615
Cbr8 netL8 0 1.1765680880374107e-19

* Branch 9
Rabr9 node_4 netRa9 -85006.53816780416
Lbr9 netRa9 netL9 -2.912333199432601e-11
Rbbr9 netL9 0 100564.90276312995
Cbr9 netL9 0 -3.51255217567515e-21

* Branch 10
Rabr10 node_4 netRa10 171311549886.61917
Lbr10 netRa10 netL10 -0.0001887794710291942
Rbbr10 netL10 0 -486556522523.7446
Cbr10 netL10 0 -2.2571552254856565e-27

* Branch 11
Rabr11 node_4 netRa11 -8348.748812307573
Lbr11 netRa11 netL11 5.6202149483281375e-12
Rbbr11 netL11 0 13917.282285318126
Cbr11 netL11 0 4.6593764589927367e-20

* Branch 12
Rabr12 node_4 netRa12 1.6629149622609998
Lbr12 netRa12 netL12 1.1234744469916549e-13
Rbbr12 netL12 0 5041.909323167262
Cbr12 netL12 0 5.819427296792271e-18

* Branch 13
Rabr13 node_4 netRa13 3817.8389991295376
Lbr13 netRa13 netL13 -3.7047295107392065e-12
Rbbr13 netL13 0 -9041.465945025677
Cbr13 netL13 0 -1.0191209282791825e-19

* Branch 14
Rabr14 node_4 netRa14 9628.041255212158
Lbr14 netRa14 netL14 8.26573607526318e-12
Rbbr14 netL14 0 -21634.92026602252
Cbr14 netL14 0 4.3709185954974845e-20

* Branch 15
Rabr15 node_4 netRa15 -171573198155.7032
Lbr15 netRa15 netL15 -0.0013120768210392255
Rbbr15 netL15 0 15936597169380.43
Cbr15 netL15 0 -4.814092221307197e-28

* Branch 16
Rabr16 node_4 netRa16 0.42486113353711974
Lbr16 netRa16 netL16 1.5590313850577744e-14
Rbbr16 netL16 0 85.37430402451949
Cbr16 netL16 0 4.018329059103816e-17

* Branch 17
Rabr17 node_4 netRa17 -7046.41468679011
Lbr17 netRa17 netL17 -2.567459217916769e-12
Rbbr17 netL17 0 8741.44771330863
Cbr17 netL17 0 -4.5003543953746575e-20

* Branch 18
Rabr18 node_4 netRa18 122.24710555378277
Lbr18 netRa18 netL18 1.8302230297664043e-13
Rbbr18 netL18 0 1072.9799324285214
Cbr18 netL18 0 3.160826836063901e-18

* Branch 19
Rabr19 node_4 netRa19 9947792867027.752
Lbr19 netRa19 netL19 0.001578049155643324
Rbbr19 netL19 0 -10377839338353.037
Cbr19 netL19 0 1.5298455547667924e-29

* Branch 20
Rabr20 node_4 netRa20 266011766.55713418
Lbr20 netRa20 netL20 -2.3566491035278986e-07
Rbbr20 netL20 0 -629559772.7811598
Cbr20 netL20 0 -1.3895060154123628e-24

* Branch 21
Rabr21 node_4 netRa21 -116217.07433632882
Lbr21 netRa21 netL21 2.6827046868713364e-10
Rbbr21 netL21 0 1157747.8793748429
Cbr21 netL21 0 1.9014581354571496e-21

* Branch 22
Rabr22 node_4 netRa22 2.1960004939173032
Lbr22 netRa22 netL22 1.205704636476202e-13
Rbbr22 netL22 0 61958.09989023261
Cbr22 netL22 0 4.702975861980888e-18

* Branch 23
Rabr23 node_4 netRa23 -1364077.5496375398
Lbr23 netRa23 netL23 -2.6470440840597693e-09
Rbbr23 netL23 0 11883460.196328267
Cbr23 netL23 0 -1.8937419138684197e-22

* Branch 24
Rabr24 node_4 netRa24 -329894.9114405251
Lbr24 netRa24 netL24 -5.355191254883824e-11
Rbbr24 netL24 0 346037.71173940966
Cbr24 netL24 0 -4.828356612960029e-22

* Branch 25
Rd node_4 0 2904.278539880657

.ends


.end
