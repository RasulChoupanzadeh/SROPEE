* netlist generated with reverse MNA (number of voltage nodes: n = 200 )

.subckt equivalent_circuit

.param Ip1=1.0
.param Ip2=0.0
.param Ip3=0.0
.param Ip4=0.0

R1_1 V1 0 -433.2008655111855
L1_1 V1 0 5.192760486397402e-13
C1_1 V1 0 -4.2514895596191865e-19

R1_2 V1 V2 21033.24474522573
L1_2 V1 V2 9.755870299560235e-12
C1_2 V1 V2 5.088173281894094e-20

R1_3 V1 V3 28414.558416370888
L1_3 V1 V3 1.2505366049950288e-11
C1_3 V1 V3 3.85152740971625e-20

R1_4 V1 V4 36131.64131865122
L1_4 V1 V4 1.6117950861426902e-11
C1_4 V1 V4 2.9905758498660504e-20

R1_5 V1 V5 8085.758942654931
L1_5 V1 V5 -8.584243037792361e-13
C1_5 V1 V5 4.905037257567655e-19

R1_6 V1 V6 15992.253839732959
L1_6 V1 V6 -3.0730151675051324e-12
C1_6 V1 V6 2.0459804072040274e-19

R1_7 V1 V7 20523.898615858845
L1_7 V1 V7 -3.5344175977096557e-12
C1_7 V1 V7 1.7959017655872924e-19

R1_8 V1 V8 27653.790321111224
L1_8 V1 V8 -3.2980966074664847e-12
C1_8 V1 V8 1.69727373413704e-19

R1_9 V1 V9 1282.6459472259633
L1_9 V1 V9 -6.198510501403288e-12
C1_9 V1 V9 -1.220265855809291e-19

R1_10 V1 V10 8293.330800499849
L1_10 V1 V10 -6.9210566071211014e-12
C1_10 V1 V10 -4.771840724853211e-20

R1_11 V1 V11 11588.080292702645
L1_11 V1 V11 -9.22925518155158e-12
C1_11 V1 V11 -5.370652639805492e-20

R1_12 V1 V12 8164.221301970933
L1_12 V1 V12 -7.533384831339332e-12
C1_12 V1 V12 -4.911128785246633e-20

R1_13 V1 V13 -4084.8057713060803
L1_13 V1 V13 -4.156886563497436e-11
C1_13 V1 V13 6.759030720072043e-20

R1_14 V1 V14 -153524.37665329513
L1_14 V1 V14 1.0969379200191717e-11
C1_14 V1 V14 -4.2833679853232345e-21

R1_15 V1 V15 -105693.99477070464
L1_15 V1 V15 7.88378589351734e-12
C1_15 V1 V15 -3.1561597856188096e-20

R1_16 V1 V16 -31831.28166855784
L1_16 V1 V16 5.574914468887453e-12
C1_16 V1 V16 -6.43939846712335e-20

R1_17 V1 V17 -8355.82787442807
L1_17 V1 V17 3.496827386977143e-12
C1_17 V1 V17 -6.965064421855997e-20

R1_18 V1 V18 -151499.28387887217
L1_18 V1 V18 9.364716365540634e-12
C1_18 V1 V18 -6.82879741013041e-20

R1_19 V1 V19 -48022.71162987769
L1_19 V1 V19 1.7769342860096163e-11
C1_19 V1 V19 -1.475131499645549e-20

R1_20 V1 V20 -30988.89172051378
L1_20 V1 V20 1.1499800395073695e-11
C1_20 V1 V20 -2.1868379075982457e-20

R1_21 V1 V21 -1391.8425258813645
L1_21 V1 V21 2.0695216029857136e-12
C1_21 V1 V21 -3.887065325532005e-20

R1_22 V1 V22 -7467.2859672934665
L1_22 V1 V22 6.6823902381456075e-12
C1_22 V1 V22 4.4665136936699105e-20

R1_23 V1 V23 -11503.949812125478
L1_23 V1 V23 6.190829655970595e-12
C1_23 V1 V23 -3.3693574922154907e-21

R1_24 V1 V24 -8120.889798737573
L1_24 V1 V24 4.756986302289507e-12
C1_24 V1 V24 -1.6240638235801425e-20

R1_25 V1 V25 1796.276193000769
L1_25 V1 V25 -2.2156095798783326e-12
C1_25 V1 V25 1.5126514693505715e-19

R1_26 V1 V26 13227.044850481216
L1_26 V1 V26 -6.186428123045896e-12
C1_26 V1 V26 8.16828385375328e-21

R1_27 V1 V27 19491.59066376986
L1_27 V1 V27 -4.332709407173538e-12
C1_27 V1 V27 7.16001432721823e-20

R1_28 V1 V28 10443.950135109537
L1_28 V1 V28 -2.810918820884939e-12
C1_28 V1 V28 1.3270526817771273e-19

R1_29 V1 V29 1958.2957637888626
L1_29 V1 V29 -3.17101610039916e-12
C1_29 V1 V29 3.159960401742501e-20

R1_30 V1 V30 23453.5293516914
L1_30 V1 V30 -7.941903559833125e-12
C1_30 V1 V30 1.7312838543258778e-20

R1_31 V1 V31 25593.040080010094
L1_31 V1 V31 -1.0480169067536881e-11
C1_31 V1 V31 -4.311986248092922e-21

R1_32 V1 V32 14516.810414010057
L1_32 V1 V32 -7.896951988761924e-12
C1_32 V1 V32 1.0086344981956899e-20

R1_33 V1 V33 3899.0619433135575
L1_33 V1 V33 1.0355393742449963e-11
C1_33 V1 V33 -6.242829392565242e-20

R1_34 V1 V34 -71475.62768575385
L1_34 V1 V34 5.1513334698561056e-11
C1_34 V1 V34 -4.391497954071495e-20

R1_35 V1 V35 -18314.578678488604
L1_35 V1 V35 1.1307483189641088e-11
C1_35 V1 V35 -5.647408188235168e-20

R1_36 V1 V36 -12660.741146200651
L1_36 V1 V36 6.290198913196221e-12
C1_36 V1 V36 -6.350181720177063e-20

R1_37 V1 V37 -3711.7799263326465
L1_37 V1 V37 2.7374114666594428e-12
C1_37 V1 V37 -1.5827400907897723e-19

R1_38 V1 V38 -20154.47719709472
L1_38 V1 V38 5.171594773675834e-12
C1_38 V1 V38 -8.729501457325276e-20

R1_39 V1 V39 -21324.408984700065
L1_39 V1 V39 9.812888387258562e-12
C1_39 V1 V39 -1.5304915138686902e-20

R1_40 V1 V40 -13645.382058446226
L1_40 V1 V40 6.393654587071256e-12
C1_40 V1 V40 -2.462412833928295e-20

R1_41 V1 V41 -82765.9474440154
L1_41 V1 V41 1.519546515813399e-11
C1_41 V1 V41 8.794088836806e-20

R1_42 V1 V42 -29106.003722578844
L1_42 V1 V42 -3.202099789811143e-11
C1_42 V1 V42 3.3920954336543675e-20

R1_43 V1 V43 -16775.806744408088
L1_43 V1 V43 2.6607872258259227e-11
C1_43 V1 V43 5.043000903196978e-21

R1_44 V1 V44 -14605.776456772017
L1_44 V1 V44 5.729500063529651e-11
C1_44 V1 V44 3.341392679590911e-20

R1_45 V1 V45 3968.2034941092134
L1_45 V1 V45 -4.296094197687357e-12
C1_45 V1 V45 6.300217297217242e-20

R1_46 V1 V46 377395.64819347207
L1_46 V1 V46 -8.403322194735864e-12
C1_46 V1 V46 6.948761335640716e-20

R1_47 V1 V47 168670.74349632123
L1_47 V1 V47 -9.019063007167118e-12
C1_47 V1 V47 4.701571523092279e-20

R1_48 V1 V48 23883.980310853694
L1_48 V1 V48 -4.71729272496756e-12
C1_48 V1 V48 9.010838548784392e-20

R1_49 V1 V49 3278.174780831463
L1_49 V1 V49 -1.7493099117998892e-11
C1_49 V1 V49 3.404535738560236e-20

R1_50 V1 V50 -46106.96547803912
L1_50 V1 V50 9.19846171010106e-11
C1_50 V1 V50 -3.118739241931117e-20

R1_51 V1 V51 -3546255.6222161516
L1_51 V1 V51 -1.2532599948488711e-11
C1_51 V1 V51 8.782968287223054e-21

R1_52 V1 V52 -44827.91493094889
L1_52 V1 V52 -3.2380544473021275e-11
C1_52 V1 V52 2.897566934918742e-21

R1_53 V1 V53 7966.599967224096
L1_53 V1 V53 -1.1389437432942609e-11
C1_53 V1 V53 -4.9138124651773734e-20

R1_54 V1 V54 38930.8783427592
L1_54 V1 V54 1.8932550746501918e-11
C1_54 V1 V54 -7.096425953641355e-20

R1_55 V1 V55 26014.273012537014
L1_55 V1 V55 1.0315643023746129e-10
C1_55 V1 V55 -4.189749856233985e-20

R1_56 V1 V56 64420.75287517149
L1_56 V1 V56 9.286848916979311e-12
C1_56 V1 V56 -7.913704417706799e-20

R1_57 V1 V57 -38421.31476838835
L1_57 V1 V57 2.3112164197867203e-12
C1_57 V1 V57 -1.6203473447240304e-19

R1_58 V1 V58 -18140.31356759425
L1_58 V1 V58 -2.957279574226211e-11
C1_58 V1 V58 1.8787189620901288e-20

R1_59 V1 V59 -10533.073912132208
L1_59 V1 V59 2.2939805449849055e-11
C1_59 V1 V59 1.3102791390137918e-20

R1_60 V1 V60 -7418.960223943149
L1_60 V1 V60 1.2119473641693757e-11
C1_60 V1 V60 2.0399598085547285e-20

R1_61 V1 V61 -125003.47391031745
L1_61 V1 V61 -3.6153887924305402e-12
C1_61 V1 V61 1.7085745787157726e-19

R1_62 V1 V62 -215955.96815793717
L1_62 V1 V62 -2.5480880278853105e-10
C1_62 V1 V62 2.0688897834999194e-20

R1_63 V1 V63 -51982.024418905814
L1_63 V1 V63 1.2025332264422603e-11
C1_63 V1 V63 -3.578393449192641e-20

R1_64 V1 V64 169369.95586412295
L1_64 V1 V64 8.371277280194475e-10
C1_64 V1 V64 4.6862851045099305e-21

R1_65 V1 V65 4471.494562048301
L1_65 V1 V65 9.22629551241542e-11
C1_65 V1 V65 1.9255761633527448e-20

R1_66 V1 V66 -31918.775359712647
L1_66 V1 V66 1.3837055251096973e-11
C1_66 V1 V66 -4.9032362885560736e-20

R1_67 V1 V67 -43097.602437969115
L1_67 V1 V67 1.7186418447443537e-11
C1_67 V1 V67 -3.8002305470125236e-20

R1_68 V1 V68 -1377344.4655242066
L1_68 V1 V68 -5.2911941776306857e-11
C1_68 V1 V68 1.928375090009751e-21

R1_69 V1 V69 7362.269185643566
L1_69 V1 V69 -5.037990108303596e-12
C1_69 V1 V69 5.588731127266167e-20

R1_70 V1 V70 -110915.33597718952
L1_70 V1 V70 -1.5616509360117013e-11
C1_70 V1 V70 2.7594248106741367e-20

R1_71 V1 V71 47745.70924678057
L1_71 V1 V71 -4.875890566717937e-12
C1_71 V1 V71 8.940423273661338e-20

R1_72 V1 V72 71878.4592488347
L1_72 V1 V72 -5.361558905443738e-12
C1_72 V1 V72 6.062641963055841e-20

R1_73 V1 V73 23247.319025389446
L1_73 V1 V73 2.4260840755122577e-09
C1_73 V1 V73 -5.60280833431586e-20

R1_74 V1 V74 43119.15562383872
L1_74 V1 V74 -1.2559070518295504e-11
C1_74 V1 V74 2.6919211985194597e-20

R1_75 V1 V75 77505.37521081782
L1_75 V1 V75 -3.738734405946413e-11
C1_75 V1 V75 1.6491059691493712e-20

R1_76 V1 V76 -36351.549876455894
L1_76 V1 V76 1.0435549018588013e-11
C1_76 V1 V76 -2.2622625668107144e-20

R1_77 V1 V77 -14442.397455128157
L1_77 V1 V77 2.511858844052836e-12
C1_77 V1 V77 -1.6614695798356376e-19

R1_78 V1 V78 44417.04876356756
L1_78 V1 V78 1.4187495072029169e-11
C1_78 V1 V78 -4.4369557942007405e-20

R1_79 V1 V79 -105618.93712133387
L1_79 V1 V79 8.558278775771186e-12
C1_79 V1 V79 -5.746629211142479e-20

R1_80 V1 V80 610581.5865618695
L1_80 V1 V80 1.3852731457854921e-11
C1_80 V1 V80 -3.256153951712918e-20

R1_81 V1 V81 2324.607035749718
L1_81 V1 V81 -3.740295391744823e-12
C1_81 V1 V81 1.661723817179564e-19

R1_82 V1 V82 -15406.551513433122
L1_82 V1 V82 2.8403389235652714e-11
C1_82 V1 V82 -2.34922004416896e-20

R1_83 V1 V83 -8309.031445825127
L1_83 V1 V83 1.1109540503820842e-11
C1_83 V1 V83 -6.173635700902296e-20

R1_84 V1 V84 -9173.500285722334
L1_84 V1 V84 1.6807733486279515e-11
C1_84 V1 V84 -1.9535450261860953e-20

R1_85 V1 V85 103508.62080426975
L1_85 V1 V85 -3.0836562687406237e-11
C1_85 V1 V85 5.46683303979816e-20

R1_86 V1 V86 -7332.207514163571
L1_86 V1 V86 -7.90720276500811e-12
C1_86 V1 V86 6.204504206677429e-20

R1_87 V1 V87 -24465.364362692646
L1_87 V1 V87 -2.3291505545928898e-11
C1_87 V1 V87 3.738566851538043e-20

R1_88 V1 V88 -23282.908779715537
L1_88 V1 V88 -1.2596515042855552e-11
C1_88 V1 V88 4.5617453413980286e-20

R1_89 V1 V89 13655.015301284393
L1_89 V1 V89 -8.876263471542013e-12
C1_89 V1 V89 3.1162399882156603e-20

R1_90 V1 V90 13775.8483249114
L1_90 V1 V90 1.0595999196088378e-11
C1_90 V1 V90 -3.8269779698248665e-20

R1_91 V1 V91 12286.735560826168
L1_91 V1 V91 -4.062473983376342e-12
C1_91 V1 V91 1.2117871277490771e-19

R1_92 V1 V92 28066.28626447992
L1_92 V1 V92 -5.956421159422824e-12
C1_92 V1 V92 7.491654801471555e-20

R1_93 V1 V93 5967.8124078819155
L1_93 V1 V93 7.36697505596122e-12
C1_93 V1 V93 -1.1939961710108959e-19

R1_94 V1 V94 12464.556077418169
L1_94 V1 V94 2.3978948121890405e-11
C1_94 V1 V94 -3.8858226575980517e-20

R1_95 V1 V95 77320.31389091205
L1_95 V1 V95 8.250267008236584e-12
C1_95 V1 V95 -6.831368847877752e-20

R1_96 V1 V96 37360.3506933012
L1_96 V1 V96 5.4913656456341005e-12
C1_96 V1 V96 -8.551338230623968e-20

R1_97 V1 V97 6482.4225927328725
L1_97 V1 V97 3.673685128928817e-12
C1_97 V1 V97 -1.23705204837056e-19

R1_98 V1 V98 -4736.608834056283
L1_98 V1 V98 -7.514382516802232e-12
C1_98 V1 V98 4.062554608115842e-20

R1_99 V1 V99 -4523.706911727045
L1_99 V1 V99 6.585146770679544e-12
C1_99 V1 V99 -1.0293656134437743e-19

R1_100 V1 V100 -4565.913439555478
L1_100 V1 V100 1.3878146357572479e-11
C1_100 V1 V100 -4.60503582620461e-20

R1_101 V1 V101 -33113.659091585214
L1_101 V1 V101 -4.479956698432206e-12
C1_101 V1 V101 1.760624684061793e-19

R1_102 V1 V102 -54621.86098905163
L1_102 V1 V102 2.6033435422838287e-11
C1_102 V1 V102 -1.6117924625779984e-20

R1_103 V1 V103 197716.76019590272
L1_103 V1 V103 -9.334871333162108e-12
C1_103 V1 V103 5.1794120235464494e-20

R1_104 V1 V104 -42382.12614170785
L1_104 V1 V104 -9.20809713732414e-12
C1_104 V1 V104 7.033521267275711e-20

R1_105 V1 V105 2055.794630137923
L1_105 V1 V105 -6.0716831001184965e-12
C1_105 V1 V105 3.6020027252486626e-20

R1_106 V1 V106 -25351.92445103614
L1_106 V1 V106 1.6028923155384796e-11
C1_106 V1 V106 -3.765481505006421e-20

R1_107 V1 V107 41971.58370961075
L1_107 V1 V107 -1.9752288614151722e-11
C1_107 V1 V107 5.354785587142785e-20

R1_108 V1 V108 19545.85992750546
L1_108 V1 V108 -2.2400834606736034e-11
C1_108 V1 V108 2.864403770633891e-20

R1_109 V1 V109 -9678.15621510849
L1_109 V1 V109 1.020939859251861e-11
C1_109 V1 V109 -5.217374456913256e-20

R1_110 V1 V110 83850.60443580207
L1_110 V1 V110 -4.039029413066973e-11
C1_110 V1 V110 3.636805774456264e-20

R1_111 V1 V111 -66757.5667948957
L1_111 V1 V111 -1.505409146426831e-11
C1_111 V1 V111 6.338840012041554e-21

R1_112 V1 V112 -22278.89591018269
L1_112 V1 V112 -5.546274924104065e-11
C1_112 V1 V112 -2.6153922970576754e-20

R1_113 V1 V113 15320.796776161078
L1_113 V1 V113 6.51709770608847e-12
C1_113 V1 V113 -7.846399797056603e-20

R1_114 V1 V114 -32623.05260434585
L1_114 V1 V114 1.3864356637278293e-10
C1_114 V1 V114 -3.4172315394734435e-21

R1_115 V1 V115 -15298.229018599779
L1_115 V1 V115 7.031105438698191e-12
C1_115 V1 V115 -8.437505338542505e-20

R1_116 V1 V116 -24992.94156865167
L1_116 V1 V116 9.216614431202457e-12
C1_116 V1 V116 -6.884911561785159e-20

R1_117 V1 V117 5667.0589618732265
L1_117 V1 V117 5.657868701910951e-12
C1_117 V1 V117 -7.639606405520157e-20

R1_118 V1 V118 -152282.469580746
L1_118 V1 V118 -2.219289212282915e-11
C1_118 V1 V118 -8.5440880083873e-21

R1_119 V1 V119 -35828.80019264507
L1_119 V1 V119 -3.1480548199417985e-11
C1_119 V1 V119 3.35048009449378e-20

R1_120 V1 V120 -14979.821061662537
L1_120 V1 V120 -9.676997301462743e-11
C1_120 V1 V120 2.0548484378334244e-20

R1_121 V1 V121 12356.410536902353
L1_121 V1 V121 -2.9849600970828364e-12
C1_121 V1 V121 2.231991417692359e-19

R1_122 V1 V122 -31795.708975748996
L1_122 V1 V122 -4.5280053717208775e-11
C1_122 V1 V122 1.6061407650692384e-20

R1_123 V1 V123 22789.784890549785
L1_123 V1 V123 -1.0399963929398953e-11
C1_123 V1 V123 1.57399680729213e-20

R1_124 V1 V124 14685.828473923964
L1_124 V1 V124 -7.680067509914238e-12
C1_124 V1 V124 6.206927889991052e-20

R1_125 V1 V125 3468.2477308507973
L1_125 V1 V125 -5.198573314962173e-12
C1_125 V1 V125 1.7140614858217986e-20

R1_126 V1 V126 -456946.2219567506
L1_126 V1 V126 -2.749384078907511e-11
C1_126 V1 V126 5.2862059689775855e-20

R1_127 V1 V127 -66056.232949783
L1_127 V1 V127 1.602717050067083e-11
C1_127 V1 V127 2.844731145657341e-21

R1_128 V1 V128 39105.144225367316
L1_128 V1 V128 2.4267010617401318e-11
C1_128 V1 V128 -1.0099461968202274e-20

R1_129 V1 V129 -20024.16579736368
L1_129 V1 V129 3.85567577045788e-12
C1_129 V1 V129 -1.1056908959365683e-19

R1_130 V1 V130 5930563.449434934
L1_130 V1 V130 9.836352720639507e-12
C1_130 V1 V130 -6.563662900439304e-20

R1_131 V1 V131 -64796.64800483162
L1_131 V1 V131 -2.8472107622572148e-11
C1_131 V1 V131 -2.4616145989115028e-20

R1_132 V1 V132 -9570.258345959568
L1_132 V1 V132 7.128441676687627e-11
C1_132 V1 V132 -5.722234059087768e-20

R1_133 V1 V133 -4913.297020952164
L1_133 V1 V133 1.1396948254152466e-11
C1_133 V1 V133 -1.1852087101304207e-20

R1_134 V1 V134 -8597.219226070167
L1_134 V1 V134 3.951550743344918e-11
C1_134 V1 V134 2.3108450609909577e-20

R1_135 V1 V135 67863.1546880637
L1_135 V1 V135 5.147777708211162e-11
C1_135 V1 V135 1.3062623970958225e-20

R1_136 V1 V136 17808.695075996235
L1_136 V1 V136 -7.771704198013538e-11
C1_136 V1 V136 1.8065788764292925e-20

R1_137 V1 V137 4459.748074715231
L1_137 V1 V137 4.853796392444144e-12
C1_137 V1 V137 -1.0880406064650644e-19

R1_138 V1 V138 5583.213508003735
L1_138 V1 V138 -9.908869059593787e-12
C1_138 V1 V138 3.9202845437661864e-20

R1_139 V1 V139 -22602.799535939706
L1_139 V1 V139 1.3530899611202185e-10
C1_139 V1 V139 6.1498005226172715e-21

R1_140 V1 V140 -24036.48030560717
L1_140 V1 V140 2.391624960138779e-11
C1_140 V1 V140 -2.8080481715169925e-20

R1_141 V1 V141 -13728.651953580178
L1_141 V1 V141 -2.776556351193857e-12
C1_141 V1 V141 1.8808155588203313e-19

R1_142 V1 V142 -7812.5838564327905
L1_142 V1 V142 1.3466182675468778e-10
C1_142 V1 V142 -1.4567605870069264e-20

R1_143 V1 V143 -17222.53704790176
L1_143 V1 V143 8.906638809904943e-11
C1_143 V1 V143 -2.69105102596482e-20

R1_144 V1 V144 -9989.497689866665
L1_144 V1 V144 -3.284776237468952e-11
C1_144 V1 V144 5.142148115628731e-20

R1_145 V1 V145 2713.52597642631
L1_145 V1 V145 -2.9335960201979028e-12
C1_145 V1 V145 1.5830244964786747e-19

R1_146 V1 V146 -11225.460070475563
L1_146 V1 V146 9.285741762218025e-11
C1_146 V1 V146 -3.3853967861125076e-20

R1_147 V1 V147 16563.489890684537
L1_147 V1 V147 -7.136736549394724e-12
C1_147 V1 V147 1.1447468580601515e-19

R1_148 V1 V148 6191.579326175332
L1_148 V1 V148 -6.100538254267854e-12
C1_148 V1 V148 4.81921243447446e-20

R1_149 V1 V149 -1877.0419248440087
L1_149 V1 V149 2.526334932863073e-12
C1_149 V1 V149 -2.0621029483518728e-19

R1_150 V1 V150 6531.452496200777
L1_150 V1 V150 -6.986267458476036e-12
C1_150 V1 V150 5.949827795462177e-20

R1_151 V1 V151 7852.77580814898
L1_151 V1 V151 -1.1470355835581438e-11
C1_151 V1 V151 -2.9284411103722757e-20

R1_152 V1 V152 -12453.474618285562
L1_152 V1 V152 2.2881643790184266e-11
C1_152 V1 V152 -2.6439235389247303e-20

R1_153 V1 V153 3409.3973847185352
L1_153 V1 V153 3.0386598688761846e-12
C1_153 V1 V153 -2.011413108633726e-19

R1_154 V1 V154 -20320.435270397596
L1_154 V1 V154 5.5846061175418485e-12
C1_154 V1 V154 -6.267253917587139e-20

R1_155 V1 V155 -4508.332511173043
L1_155 V1 V155 5.545638863652873e-12
C1_155 V1 V155 1.87105430764508e-20

R1_156 V1 V156 -175642.96413998908
L1_156 V1 V156 1.0563111451822095e-11
C1_156 V1 V156 -8.053220789885655e-20

R1_157 V1 V157 2984.2570533949056
L1_157 V1 V157 -2.555784478843366e-11
C1_157 V1 V157 4.922043846924117e-20

R1_158 V1 V158 -12940.108609893708
L1_158 V1 V158 9.9848064131543e-11
C1_158 V1 V158 -2.5134976269365084e-20

R1_159 V1 V159 -156728.16004517357
L1_159 V1 V159 1.0991797196818971e-11
C1_159 V1 V159 -9.734345923026326e-20

R1_160 V1 V160 -10689.619858401502
L1_160 V1 V160 1.0494105161151775e-11
C1_160 V1 V160 6.469435229305657e-21

R1_161 V1 V161 6244.063708361071
L1_161 V1 V161 -2.906907225087815e-12
C1_161 V1 V161 2.5603144167376583e-19

R1_162 V1 V162 -20838.545844041164
L1_162 V1 V162 -1.255917091612422e-09
C1_162 V1 V162 -7.314761354933933e-20

R1_163 V1 V163 -6811.545493569763
L1_163 V1 V163 -1.3083691173037734e-10
C1_163 V1 V163 -2.0359470998010938e-20

R1_164 V1 V164 -41715.45050423147
L1_164 V1 V164 -7.769907701632838e-12
C1_164 V1 V164 3.1293004988886142e-21

R1_165 V1 V165 3769.9244320733555
L1_165 V1 V165 -8.448624441386765e-12
C1_165 V1 V165 -4.3772585393171665e-20

R1_166 V1 V166 -10752.730951500404
L1_166 V1 V166 -3.8416078789827904e-12
C1_166 V1 V166 1.0914183472624206e-19

R1_167 V1 V167 23975.151377997205
L1_167 V1 V167 -4.830765883435893e-12
C1_167 V1 V167 7.190036901018617e-20

R1_168 V1 V168 -7289.76679520018
L1_168 V1 V168 -6.2840477268610235e-12
C1_168 V1 V168 1.3883487322336897e-19

R1_169 V1 V169 -167427.2543456973
L1_169 V1 V169 4.588403568040735e-12
C1_169 V1 V169 -1.5363217175752873e-19

R1_170 V1 V170 3639.7882944403223
L1_170 V1 V170 1.1599091548690213e-11
C1_170 V1 V170 -2.1748389327683454e-20

R1_171 V1 V171 4490.663879800782
L1_171 V1 V171 7.368709435407177e-11
C1_171 V1 V171 2.4338476666381833e-20

R1_172 V1 V172 5782.025417872222
L1_172 V1 V172 1.4467792399548949e-11
C1_172 V1 V172 -4.353330765747404e-20

R1_173 V1 V173 4816.43296867582
L1_173 V1 V173 9.850642128684524e-12
C1_173 V1 V173 -4.790730308968187e-20

R1_174 V1 V174 -4026.375182053689
L1_174 V1 V174 2.1607463045312885e-12
C1_174 V1 V174 -1.6430047187674553e-19

R1_175 V1 V175 -3669.818157487335
L1_175 V1 V175 2.9650566044376608e-12
C1_175 V1 V175 -1.4399721955291112e-19

R1_176 V1 V176 -4212.518407314408
L1_176 V1 V176 2.4743918726716855e-12
C1_176 V1 V176 -1.7116525775389533e-19

R1_177 V1 V177 -15411.933662629253
L1_177 V1 V177 -3.195059078914938e-11
C1_177 V1 V177 1.0030509732635147e-19

R1_178 V1 V178 34216.04274132612
L1_178 V1 V178 -4.605958081335834e-12
C1_178 V1 V178 6.032740978489563e-20

R1_179 V1 V179 -956823.8289146698
L1_179 V1 V179 -5.935229195673792e-12
C1_179 V1 V179 6.617936482964584e-20

R1_180 V1 V180 13242.13342583944
L1_180 V1 V180 -3.4602039692942435e-12
C1_180 V1 V180 1.0621644320612716e-19

R1_181 V1 V181 -5272.854533966659
L1_181 V1 V181 -1.3607936292255234e-11
C1_181 V1 V181 1.429126931332978e-19

R1_182 V1 V182 10143.320789522568
L1_182 V1 V182 -1.419625437207456e-11
C1_182 V1 V182 3.6898230128784884e-21

R1_183 V1 V183 9463.955186638907
L1_183 V1 V183 -2.6291584333404103e-11
C1_183 V1 V183 -1.8426664171018772e-22

R1_184 V1 V184 8114.691551930211
L1_184 V1 V184 -8.669873775660176e-12
C1_184 V1 V184 3.071818298893331e-20

R1_185 V1 V185 2041.3849135050223
L1_185 V1 V185 -4.171630350399828e-12
C1_185 V1 V185 -1.5785715814269495e-19

R1_186 V1 V186 -6930.099624435893
L1_186 V1 V186 -9.039867703019595e-12
C1_186 V1 V186 9.12755394145139e-20

R1_187 V1 V187 -58790.64543741401
L1_187 V1 V187 -1.8837077598547787e-11
C1_187 V1 V187 1.9925045952642708e-20

R1_188 V1 V188 -31790.797891329203
L1_188 V1 V188 -2.68761758255661e-10
C1_188 V1 V188 2.841496797841405e-20

R1_189 V1 V189 -1975.7399932474978
L1_189 V1 V189 4.474843679206596e-12
C1_189 V1 V189 3.500324419641485e-21

R1_190 V1 V190 99526.78063460374
L1_190 V1 V190 1.4594304733842032e-11
C1_190 V1 V190 -2.341319433771314e-20

R1_191 V1 V191 7777.188432070167
L1_191 V1 V191 -8.115932914663875e-11
C1_191 V1 V191 -6.041372343630178e-21

R1_192 V1 V192 17823.940689859992
L1_192 V1 V192 8.854140200176688e-12
C1_192 V1 V192 -7.2979622828716e-20

R1_193 V1 V193 -23562.290137010932
L1_193 V1 V193 5.527786823612293e-12
C1_193 V1 V193 -5.428750155437893e-20

R1_194 V1 V194 8542.87542082846
L1_194 V1 V194 3.874062244786085e-12
C1_194 V1 V194 -1.4142903123447241e-19

R1_195 V1 V195 -69942.88389647102
L1_195 V1 V195 3.322423247894866e-11
C1_195 V1 V195 -5.561472864763809e-21

R1_196 V1 V196 -43650.24173144481
L1_196 V1 V196 6.321720542457309e-12
C1_196 V1 V196 -5.603657680786646e-20

R1_197 V1 V197 3100.894144686381
L1_197 V1 V197 -6.27835755529152e-12
C1_197 V1 V197 1.2532290350119897e-19

R1_198 V1 V198 -8066.555508861803
L1_198 V1 V198 -2.1051605329974118e-11
C1_198 V1 V198 1.2932679962706811e-21

R1_199 V1 V199 -4409.237250214629
L1_199 V1 V199 1.5590115355222516e-11
C1_199 V1 V199 -7.837173608001203e-20

R1_200 V1 V200 -7074.886407635252
L1_200 V1 V200 -6.966818249024695e-12
C1_200 V1 V200 1.046221381553623e-19

R2_2 V2 0 -3947.2127938146505
L2_2 V2 0 1.282323907081617e-12
C2_2 V2 0 -1.1352961796563434e-18

R2_3 V2 V3 51151.09987768509
L2_3 V2 V3 8.084659153896639e-12
C2_3 V2 V3 5.996654735514636e-20

R2_4 V2 V4 51371.407842152315
L2_4 V2 V4 9.089595694648935e-12
C2_4 V2 V4 5.287397361997769e-20

R2_5 V2 V5 -21728.584144459757
L2_5 V2 V5 3.1262426878497493e-12
C2_5 V2 V5 -1.5365401833383227e-19

R2_6 V2 V6 5681.357879210301
L2_6 V2 V6 -6.235535157734272e-13
C2_6 V2 V6 7.996145137128471e-19

R2_7 V2 V7 25003.004920492236
L2_7 V2 V7 -2.9968601994551206e-12
C2_7 V2 V7 2.231898040230324e-19

R2_8 V2 V8 43189.36601194046
L2_8 V2 V8 -3.4522885336519804e-12
C2_8 V2 V8 1.7930582491718645e-19

R2_9 V2 V9 -3571.471456631513
L2_9 V2 V9 -2.2759935692414488e-11
C2_9 V2 V9 5.226977305645436e-20

R2_10 V2 V10 4683.934999485386
L2_10 V2 V10 2.7158059983748377e-12
C2_10 V2 V10 -4.6154312642058276e-20

R2_11 V2 V11 -34782.501403193884
L2_11 V2 V11 1.268233836679461e-11
C2_11 V2 V11 -8.661448787713107e-20

R2_12 V2 V12 -24768.292814777633
L2_12 V2 V12 1.614000462607672e-11
C2_12 V2 V12 -7.131951394230556e-20

R2_13 V2 V13 11954.508974600209
L2_13 V2 V13 2.4627955970457677e-11
C2_13 V2 V13 -5.365508111418027e-20

R2_14 V2 V14 -5709.837992559466
L2_14 V2 V14 1.6158337957451786e-12
C2_14 V2 V14 -4.127052794970795e-19

R2_15 V2 V15 -28309.528751114365
L2_15 V2 V15 4.171299128415499e-12
C2_15 V2 V15 -1.1615488109782054e-19

R2_16 V2 V16 -21859.391362847135
L2_16 V2 V16 3.079985670848394e-12
C2_16 V2 V16 -1.7380989607108066e-19

R2_17 V2 V17 15625.122231482628
L2_17 V2 V17 -8.475169783087644e-12
C2_17 V2 V17 3.671442424229877e-20

R2_18 V2 V18 -13359.930135985836
L2_18 V2 V18 -1.2402039232683565e-11
C2_18 V2 V18 1.119866537255545e-19

R2_19 V2 V19 242486.16263565654
L2_19 V2 V19 -1.0867483418997329e-11
C2_19 V2 V19 6.10146219668099e-20

R2_20 V2 V20 145845.33450865743
L2_20 V2 V20 -9.328698836043919e-12
C2_20 V2 V20 6.978141668714238e-20

R2_21 V2 V21 4090.3188325814203
L2_21 V2 V21 -2.166039059721541e-09
C2_21 V2 V21 -4.459443989485718e-20

R2_22 V2 V22 -6582.392546898529
L2_22 V2 V22 -4.755815877578012e-12
C2_22 V2 V22 4.6702142844388687e-20

R2_23 V2 V23 88915.30137205697
L2_23 V2 V23 6.485262088128274e-11
C2_23 V2 V23 7.655630656802584e-21

R2_24 V2 V24 46229.37514129151
L2_24 V2 V24 3.4807031694277315e-11
C2_24 V2 V24 -3.7759601800345425e-21

R2_25 V2 V25 -5120.2484153207915
L2_25 V2 V25 6.548685704842858e-12
C2_25 V2 V25 -4.7655330152529145e-20

R2_26 V2 V26 6364.678631463607
L2_26 V2 V26 -9.771079260898798e-11
C2_26 V2 V26 6.191596458666666e-20

R2_27 V2 V27 109696.76200317244
L2_27 V2 V27 -3.518685437161708e-11
C2_27 V2 V27 -6.5813682437385466e-21

R2_28 V2 V28 128105.1325668743
L2_28 V2 V28 -1.2315043739420697e-11
C2_28 V2 V28 2.725329766582499e-20

R2_29 V2 V29 -5638.439352168632
L2_29 V2 V29 -6.783966268467567e-12
C2_29 V2 V29 1.142653813253053e-19

R2_30 V2 V30 6185.298445666664
L2_30 V2 V30 4.579187840913254e-12
C2_30 V2 V30 -7.104146547408982e-20

R2_31 V2 V31 45194.443429088795
L2_31 V2 V31 -2.715164543883303e-11
C2_31 V2 V31 2.0482068744356456e-22

R2_32 V2 V32 46906.035285929596
L2_32 V2 V32 -1.7227008605069945e-11
C2_32 V2 V32 1.7248095878145407e-20

R2_33 V2 V33 -8074.041657281745
L2_33 V2 V33 3.644855026912059e-12
C2_33 V2 V33 -1.2329174953348927e-19

R2_34 V2 V34 -23757.99483999443
L2_34 V2 V34 8.883554626737506e-12
C2_34 V2 V34 6.343687756674954e-20

R2_35 V2 V35 -27074.957679845757
L2_35 V2 V35 6.608832672623858e-12
C2_35 V2 V35 -8.422947261144494e-20

R2_36 V2 V36 -19730.747495228672
L2_36 V2 V36 5.0176106628153804e-12
C2_36 V2 V36 -1.0091207874443989e-19

R2_37 V2 V37 10482.887874198348
L2_37 V2 V37 1.569253318753826e-11
C2_37 V2 V37 -2.4701110432371008e-20

R2_38 V2 V38 -12931.520626023206
L2_38 V2 V38 4.9855275781873264e-11
C2_38 V2 V38 -4.2497135390658025e-20

R2_39 V2 V39 -137561.34792963532
L2_39 V2 V39 1.9724959119256237e-10
C2_39 V2 V39 1.5866633942802927e-20

R2_40 V2 V40 -537144.4688733565
L2_40 V2 V40 -4.405678113564933e-11
C2_40 V2 V40 3.904950814792311e-20

R2_41 V2 V41 23860.664786258752
L2_41 V2 V41 -4.418812165128961e-12
C2_41 V2 V41 8.422594435025851e-20

R2_42 V2 V42 -17559.10462812444
L2_42 V2 V42 5.489347309705055e-12
C2_42 V2 V42 -6.801338214713285e-20

R2_43 V2 V43 70794.35416572039
L2_43 V2 V43 -2.611237135260247e-11
C2_43 V2 V43 -3.985347323106561e-21

R2_44 V2 V44 36621.55987463979
L2_44 V2 V44 -1.2602738777406532e-11
C2_44 V2 V44 1.1170143920411376e-20

R2_45 V2 V45 -15464.753351420066
L2_45 V2 V45 -7.972875880758374e-12
C2_45 V2 V45 7.990246894681325e-20

R2_46 V2 V46 5928.129186287715
L2_46 V2 V46 -2.022151444338123e-12
C2_46 V2 V46 2.22261451290948e-19

R2_47 V2 V47 24881.14929277724
L2_47 V2 V47 -5.151763179925213e-12
C2_47 V2 V47 8.147996837489534e-20

R2_48 V2 V48 18008.16191602096
L2_48 V2 V48 -3.6917553452141e-12
C2_48 V2 V48 1.1562799369641462e-19

R2_49 V2 V49 -7523.869102389553
L2_49 V2 V49 7.358974154337044e-12
C2_49 V2 V49 -6.813254736137028e-20

R2_50 V2 V50 15037.708231106302
L2_50 V2 V50 4.493731014417416e-12
C2_50 V2 V50 -7.82469033325654e-20

R2_51 V2 V51 -92898.85963380491
L2_51 V2 V51 5.47125661785553e-12
C2_51 V2 V51 -1.244549631924086e-19

R2_52 V2 V52 -48575.37147950239
L2_52 V2 V52 3.9821861605523736e-12
C2_52 V2 V52 -1.60341684244773e-19

R2_53 V2 V53 -17140.81181746265
L2_53 V2 V53 4.222373077505069e-12
C2_53 V2 V53 -8.184353822684229e-20

R2_54 V2 V54 -8261.325309244978
L2_54 V2 V54 3.926409791830662e-12
C2_54 V2 V54 -1.16279247865046e-19

R2_55 V2 V55 -17835.298733219803
L2_55 V2 V55 7.794654917709924e-12
C2_55 V2 V55 -5.301924690097811e-20

R2_56 V2 V56 -11209.87553590114
L2_56 V2 V56 4.3635227286888284e-12
C2_56 V2 V56 -9.168280952112607e-20

R2_57 V2 V57 37296.95905716223
L2_57 V2 V57 -4.1396349108330665e-12
C2_57 V2 V57 1.2384191538092212e-19

R2_58 V2 V58 15975.990085988658
L2_58 V2 V58 1.4284383087613206e-11
C2_58 V2 V58 3.089771982125447e-20

R2_59 V2 V59 17371.157132923785
L2_59 V2 V59 -3.4230163463279627e-12
C2_59 V2 V59 1.5029192722020616e-19

R2_60 V2 V60 12621.929538245991
L2_60 V2 V60 -2.508014702354499e-12
C2_60 V2 V60 2.0664866701726152e-19

R2_61 V2 V61 55596.10466998017
L2_61 V2 V61 -9.517881611698577e-11
C2_61 V2 V61 -1.7044428619654317e-20

R2_62 V2 V62 -81274.4271466117
L2_62 V2 V62 -7.810435034211128e-12
C2_62 V2 V62 4.904522102270313e-20

R2_63 V2 V63 138638.458315807
L2_63 V2 V63 1.565604426015442e-11
C2_63 V2 V63 -4.7558268098235094e-20

R2_64 V2 V64 37825.7582569555
L2_64 V2 V64 4.1005513221738595e-11
C2_64 V2 V64 -3.431595903891148e-20

R2_65 V2 V65 -15236.963339870965
L2_65 V2 V65 -1.130218790241622e-11
C2_65 V2 V65 4.183569216461101e-20

R2_66 V2 V66 10074.501750461643
L2_66 V2 V66 -5.377805333655636e-12
C2_66 V2 V66 1.4111702668914743e-19

R2_67 V2 V67 -53586.00115856938
L2_67 V2 V67 7.492589531279727e-12
C2_67 V2 V67 -8.234581094804698e-20

R2_68 V2 V68 -151386.78326839302
L2_68 V2 V68 1.0543666299762602e-11
C2_68 V2 V68 -6.853289473356732e-20

R2_69 V2 V69 -9216.36412993746
L2_69 V2 V69 2.9618457519893883e-12
C2_69 V2 V69 -1.5728889370126231e-19

R2_70 V2 V70 21712.735208965652
L2_70 V2 V70 6.373040633696887e-12
C2_70 V2 V70 -8.328908854473582e-20

R2_71 V2 V71 39806.926272696655
L2_71 V2 V71 -7.623421995046635e-12
C2_71 V2 V71 7.175657183800006e-20

R2_72 V2 V72 177566.4359942078
L2_72 V2 V72 -1.7086580534785474e-11
C2_72 V2 V72 3.8191335051140694e-20

R2_73 V2 V73 28531.2025162708
L2_73 V2 V73 -4.195598680159715e-09
C2_73 V2 V73 4.882539157191314e-20

R2_74 V2 V74 -7083.79900711623
L2_74 V2 V74 1.8351243934886754e-12
C2_74 V2 V74 -2.337459909153188e-19

R2_75 V2 V75 88577.10662793912
L2_75 V2 V75 -1.2675994177986254e-10
C2_75 V2 V75 1.906768447123168e-20

R2_76 V2 V76 -34818.07590354856
L2_76 V2 V76 6.7270020919197366e-12
C2_76 V2 V76 -4.7106384957130135e-20

R2_77 V2 V77 21475.923062935944
L2_77 V2 V77 -3.1374943685891074e-12
C2_77 V2 V77 1.6711592617459964e-19

R2_78 V2 V78 17499.113661916672
L2_78 V2 V78 -2.5218507427241046e-12
C2_78 V2 V78 2.338360022353069e-19

R2_79 V2 V79 -47379.82163181947
L2_79 V2 V79 -1.2369800839152949e-10
C2_79 V2 V79 7.102872895658574e-21

R2_80 V2 V80 49891.59624661138
L2_80 V2 V80 -5.771354536824464e-12
C2_80 V2 V80 8.036810019452763e-20

R2_81 V2 V81 -7344.0144825031775
L2_81 V2 V81 2.1382179251330088e-11
C2_81 V2 V81 -2.607726706142374e-20

R2_82 V2 V82 9396.276913975316
L2_82 V2 V82 -2.9596107378987206e-12
C2_82 V2 V82 2.066394752032837e-19

R2_83 V2 V83 31248.521333730096
L2_83 V2 V83 -7.645278834757126e-11
C2_83 V2 V83 -1.2733674378304806e-20

R2_84 V2 V84 14173.728422628501
L2_84 V2 V84 -4.390459108731985e-12
C2_84 V2 V84 9.229121157059965e-20

R2_85 V2 V85 -43659.168265899134
L2_85 V2 V85 -2.0116948375234678e-11
C2_85 V2 V85 -2.4394863348352744e-20

R2_86 V2 V86 9976.73156354526
L2_86 V2 V86 2.5493121622289006e-12
C2_86 V2 V86 -2.2761447861666565e-19

R2_87 V2 V87 81310.66683401178
L2_87 V2 V87 2.3090956527900305e-11
C2_87 V2 V87 -4.998177546887961e-20

R2_88 V2 V88 -78026.18284592715
L2_88 V2 V88 5.0583263612440945e-12
C2_88 V2 V88 -1.3064364044248059e-19

R2_89 V2 V89 -13889.887657164989
L2_89 V2 V89 3.0183247560489286e-12
C2_89 V2 V89 -1.487293446505124e-19

R2_90 V2 V90 -5640.2569422704655
L2_90 V2 V90 3.1335460588517452e-12
C2_90 V2 V90 -1.8012005761567267e-19

R2_91 V2 V91 -81672.93963102547
L2_91 V2 V91 -7.965941443915315e-12
C2_91 V2 V91 4.6909774416763635e-20

R2_92 V2 V92 -30365.702763654175
L2_92 V2 V92 3.742208925914864e-11
C2_92 V2 V92 -1.9653138079132476e-20

R2_93 V2 V93 -61283.5590453284
L2_93 V2 V93 -8.844809780997286e-12
C2_93 V2 V93 9.987660793490034e-20

R2_94 V2 V94 -17902.613459625318
L2_94 V2 V94 -2.295481192535619e-12
C2_94 V2 V94 2.185153092619327e-19

R2_95 V2 V95 238774.0773044742
L2_95 V2 V95 -9.063745520175376e-12
C2_95 V2 V95 9.059776184703881e-20

R2_96 V2 V96 2906853.5348356883
L2_96 V2 V96 -5.088287446797838e-12
C2_96 V2 V96 1.433598051383293e-19

R2_97 V2 V97 -18998.954035652503
L2_97 V2 V97 -2.247639371266265e-12
C2_97 V2 V97 2.4207467505880054e-19

R2_98 V2 V98 3931.799101409657
L2_98 V2 V98 1.4655169998669882e-11
C2_98 V2 V98 6.328676980142436e-20

R2_99 V2 V99 -49467.228726181056
L2_99 V2 V99 4.61462276238059e-12
C2_99 V2 V99 -1.6007576146559662e-19

R2_100 V2 V100 20129.04810414065
L2_100 V2 V100 -1.3111559931908727e-11
C2_100 V2 V100 -2.4736774195791205e-20

R2_101 V2 V101 74654.01196796348
L2_101 V2 V101 3.1614678303238566e-12
C2_101 V2 V101 -1.938697423729048e-19

R2_102 V2 V102 -7682.766106337674
L2_102 V2 V102 2.8331766280778396e-12
C2_102 V2 V102 -1.6790268600794074e-19

R2_103 V2 V103 42457.44439819088
L2_103 V2 V103 5.891548174668108e-12
C2_103 V2 V103 -1.0382678002090115e-19

R2_104 V2 V104 23488.71529955998
L2_104 V2 V104 5.824084689999807e-12
C2_104 V2 V104 -1.1199092631341547e-19

R2_105 V2 V105 -5016.375036264275
L2_105 V2 V105 3.086050927275787e-12
C2_105 V2 V105 -1.613446525936265e-19

R2_106 V2 V106 4762.185371350179
L2_106 V2 V106 -5.275373677442056e-12
C2_106 V2 V106 3.611161356047456e-20

R2_107 V2 V107 13948.583353616761
L2_107 V2 V107 -2.6346180717332978e-12
C2_107 V2 V107 2.031371163043152e-19

R2_108 V2 V108 -42434.58778276659
L2_108 V2 V108 3.4550161368057034e-11
C2_108 V2 V108 5.330977839064699e-21

R2_109 V2 V109 52473.92183094867
L2_109 V2 V109 -3.444837923100944e-12
C2_109 V2 V109 1.8620909517654889e-19

R2_110 V2 V110 -9850.834301696515
L2_110 V2 V110 -3.999167610072619e-11
C2_110 V2 V110 7.415090793871676e-20

R2_111 V2 V111 99480.72813517995
L2_111 V2 V111 -1.1602378481761928e-11
C2_111 V2 V111 2.3447629012077787e-20

R2_112 V2 V112 64184.899989216334
L2_112 V2 V112 -7.355901628769762e-12
C2_112 V2 V112 5.32849954655172e-20

R2_113 V2 V113 14972.52552468496
L2_113 V2 V113 -2.9238168907455273e-12
C2_113 V2 V113 1.9593618659110997e-19

R2_114 V2 V114 -8027.835304559882
L2_114 V2 V114 1.0218256968820369e-11
C2_114 V2 V114 2.7494982639536345e-20

R2_115 V2 V115 -10882.280801405515
L2_115 V2 V115 2.2847363373127415e-12
C2_115 V2 V115 -1.674699315465428e-19

R2_116 V2 V116 -43411.73255404721
L2_116 V2 V116 1.0412510408672985e-11
C2_116 V2 V116 -1.1803178932543595e-21

R2_117 V2 V117 -7815.602896909019
L2_117 V2 V117 4.084560295607952e-12
C2_117 V2 V117 -1.2965577430422313e-19

R2_118 V2 V118 4635.514458429497
L2_118 V2 V118 1.3201235797648853e-11
C2_118 V2 V118 -1.2334214634974352e-19

R2_119 V2 V119 13723.537914459539
L2_119 V2 V119 -1.0467841466809727e-11
C2_119 V2 V119 7.93732845063361e-21

R2_120 V2 V120 19050.171887943132
L2_120 V2 V120 2.192192826918392e-11
C2_120 V2 V120 -6.929955724661506e-20

R2_121 V2 V121 -21789.23764532159
L2_121 V2 V121 2.7084192635631523e-12
C2_121 V2 V121 -1.9882335888032425e-19

R2_122 V2 V122 16968.614462500176
L2_122 V2 V122 -5.138927000896704e-12
C2_122 V2 V122 1.5059577665764203e-19

R2_123 V2 V123 17033.560168055577
L2_123 V2 V123 -6.9206475602060365e-12
C2_123 V2 V123 6.028102016042891e-20

R2_124 V2 V124 22388.46464963976
L2_124 V2 V124 -1.1669651588682776e-11
C2_124 V2 V124 3.2988364754075085e-20

R2_125 V2 V125 -41554.40344448865
L2_125 V2 V125 -4.859120683555464e-12
C2_125 V2 V125 9.114456418526473e-20

R2_126 V2 V126 -11749.016869216604
L2_126 V2 V126 -1.9584777618950512e-10
C2_126 V2 V126 -7.637808294020208e-21

R2_127 V2 V127 -12655.517901577627
L2_127 V2 V127 7.435371080910416e-11
C2_127 V2 V127 6.328682317131058e-20

R2_128 V2 V128 -10994.140868265215
L2_128 V2 V128 -3.5030094598867004e-10
C2_128 V2 V128 7.315944915224488e-20

R2_129 V2 V129 58922.85920967405
L2_129 V2 V129 -1.917358630487276e-12
C2_129 V2 V129 3.2310559418992005e-19

R2_130 V2 V130 -10740.441429894528
L2_130 V2 V130 2.444686980872914e-12
C2_130 V2 V130 -1.4744958480584885e-19

R2_131 V2 V131 15036.125097238177
L2_131 V2 V131 8.942460051286614e-11
C2_131 V2 V131 -6.078972428401008e-20

R2_132 V2 V132 10295.121233849964
L2_132 V2 V132 9.19112654132971e-12
C2_132 V2 V132 -1.2249112680246717e-19

R2_133 V2 V133 -27515.34518293011
L2_133 V2 V133 1.5526912446427553e-12
C2_133 V2 V133 -3.099143652897946e-19

R2_134 V2 V134 3125.0805629130177
L2_134 V2 V134 -1.4636334725793986e-12
C2_134 V2 V134 3.5129080072007234e-19

R2_135 V2 V135 39930.025016130334
L2_135 V2 V135 6.239907733417776e-12
C2_135 V2 V135 -7.5244785180186e-20

R2_136 V2 V136 15844.836363175253
L2_136 V2 V136 6.068639774288264e-11
C2_136 V2 V136 -2.8691271243003038e-21

R2_137 V2 V137 96108.70453701158
L2_137 V2 V137 4.9330380357344175e-12
C2_137 V2 V137 -1.5420785333315475e-19

R2_138 V2 V138 -5236.7920779339
L2_138 V2 V138 2.8295444295051465e-12
C2_138 V2 V138 -2.173587018491714e-19

R2_139 V2 V139 -11284.59567269157
L2_139 V2 V139 1.3450098658671354e-11
C2_139 V2 V139 1.2310139920219288e-20

R2_140 V2 V140 -14454.069194242367
L2_140 V2 V140 -1.8675159076907355e-10
C2_140 V2 V140 5.2412794061448324e-20

R2_141 V2 V141 6325.955995791438
L2_141 V2 V141 -1.3183046603982534e-12
C2_141 V2 V141 4.2298034909879702e-19

R2_142 V2 V142 -3848.4891557163405
L2_142 V2 V142 1.3979311131246911e-12
C2_142 V2 V142 -1.0167167044095471e-19

R2_143 V2 V143 7597.987694064969
L2_143 V2 V143 -2.88888513572017e-12
C2_143 V2 V143 1.532164737588975e-19

R2_144 V2 V144 262368.63231350295
L2_144 V2 V144 -1.8956174190222757e-11
C2_144 V2 V144 4.111543368346178e-20

R2_145 V2 V145 -4260.136635383206
L2_145 V2 V145 -2.0577357410967666e-11
C2_145 V2 V145 1.0168605290804951e-19

R2_146 V2 V146 2267.6739608730513
L2_146 V2 V146 -1.2165261098312498e-12
C2_146 V2 V146 8.456991973077867e-20

R2_147 V2 V147 -11128.494661222914
L2_147 V2 V147 1.814876350915134e-11
C2_147 V2 V147 -3.328756780669465e-20

R2_148 V2 V148 7173.8591703744705
L2_148 V2 V148 -9.636740435306434e-12
C2_148 V2 V148 -2.3067527243286822e-20

R2_149 V2 V149 21403.27599979112
L2_149 V2 V149 7.886034096384682e-13
C2_149 V2 V149 -6.513496439745446e-19

R2_150 V2 V150 6969.633427061802
L2_150 V2 V150 -5.8206527652910575e-12
C2_150 V2 V150 3.9083861397390575e-19

R2_151 V2 V151 -15478.082570438346
L2_151 V2 V151 4.265997047377252e-12
C2_151 V2 V151 -1.3735818236940122e-19

R2_152 V2 V152 -3872.9798547880073
L2_152 V2 V152 9.692022968231367e-12
C2_152 V2 V152 1.4080058656329147e-20

R2_153 V2 V153 -444713.21159377164
L2_153 V2 V153 -1.2063594843724811e-11
C2_153 V2 V153 1.5082932234957455e-22

R2_154 V2 V154 -4499.73029888938
L2_154 V2 V154 3.4714278226522205e-12
C2_154 V2 V154 -3.4700298233731356e-19

R2_155 V2 V155 -7853.147263622015
L2_155 V2 V155 4.875350044591296e-12
C2_155 V2 V155 -5.377156909481969e-20

R2_156 V2 V156 2986.6144918476007
L2_156 V2 V156 8.871059834027693e-11
C2_156 V2 V156 -4.698957118230753e-20

R2_157 V2 V157 87305.63596575781
L2_157 V2 V157 -8.543361160748192e-13
C2_157 V2 V157 6.383573179619277e-19

R2_158 V2 V158 -351329.4768474444
L2_158 V2 V158 2.947946119308453e-12
C2_158 V2 V158 4.0386245485034434e-20

R2_159 V2 V159 3356.4885448754426
L2_159 V2 V159 -5.478159660433594e-12
C2_159 V2 V159 -2.808315536803274e-20

R2_160 V2 V160 18848.95789101654
L2_160 V2 V160 -2.7872858151392075e-10
C2_160 V2 V160 -5.965230998896724e-20

R2_161 V2 V161 -6037.10118056952
L2_161 V2 V161 1.9211638208642173e-11
C2_161 V2 V161 -2.4413496441983558e-20

R2_162 V2 V162 11027.37442402536
L2_162 V2 V162 1.2132794097582327e-11
C2_162 V2 V162 -3.125997540390474e-20

R2_163 V2 V163 -59331.43262398777
L2_163 V2 V163 -3.909036769690637e-12
C2_163 V2 V163 1.68035064614189e-19

R2_164 V2 V164 -24599.65551169494
L2_164 V2 V164 -1.8427826882870925e-11
C2_164 V2 V164 2.295920281283784e-20

R2_165 V2 V165 -18098.498012458047
L2_165 V2 V165 1.3564199373729397e-12
C2_165 V2 V165 -3.714567810830508e-19

R2_166 V2 V166 3783.8818283221926
L2_166 V2 V166 -1.0262971184723187e-11
C2_166 V2 V166 7.347055328984737e-21

R2_167 V2 V167 75619.82974118984
L2_167 V2 V167 3.302200366236546e-11
C2_167 V2 V167 -1.0083226310378368e-20

R2_168 V2 V168 -13989.739393953132
L2_168 V2 V168 -1.523368955781692e-11
C2_168 V2 V168 1.0212821487070293e-19

R2_169 V2 V169 9720.6140510794
L2_169 V2 V169 -1.7149597530541897e-11
C2_169 V2 V169 5.145465941442965e-20

R2_170 V2 V170 -2801.812485344662
L2_170 V2 V170 8.61401635397508e-12
C2_170 V2 V170 -1.5624232399754173e-19

R2_171 V2 V171 -6291.730484127394
L2_171 V2 V171 1.6669995632870973e-12
C2_171 V2 V171 -2.8624474062319684e-19

R2_172 V2 V172 150736.49447579787
L2_172 V2 V172 2.9819131589857163e-12
C2_172 V2 V172 -1.6628142198140664e-19

R2_173 V2 V173 -7437.286570854511
L2_173 V2 V173 -2.727063243049491e-12
C2_173 V2 V173 1.4975429028027436e-19

R2_174 V2 V174 -17172.40672294747
L2_174 V2 V174 1.814381376363447e-11
C2_174 V2 V174 2.1151761863404725e-19

R2_175 V2 V175 9432.194411577531
L2_175 V2 V175 7.283136790176314e-11
C2_175 V2 V175 -9.56517672588634e-21

R2_176 V2 V176 9565.695090426012
L2_176 V2 V176 -5.6141010079320024e-11
C2_176 V2 V176 -6.2581415455776624e-21

R2_177 V2 V177 9239.95210154769
L2_177 V2 V177 1.4992072463873177e-10
C2_177 V2 V177 -9.689055058691324e-20

R2_178 V2 V178 3500.1438851363164
L2_178 V2 V178 -2.7483798615766653e-12
C2_178 V2 V178 1.1502787870062004e-19

R2_179 V2 V179 27356.062532351825
L2_179 V2 V179 -1.7353525723586376e-12
C2_179 V2 V179 3.180175044959001e-19

R2_180 V2 V180 32259.845166076542
L2_180 V2 V180 -1.8521688593349294e-12
C2_180 V2 V180 2.1208097593517162e-19

R2_181 V2 V181 16402.853031456267
L2_181 V2 V181 1.863947190240543e-11
C2_181 V2 V181 3.4107941590152386e-20

R2_182 V2 V182 -7465.658519867417
L2_182 V2 V182 1.3397070686319475e-12
C2_182 V2 V182 -2.2697991227485714e-19

R2_183 V2 V183 10911.501412018872
L2_183 V2 V183 -4.0821340846069964e-12
C2_183 V2 V183 4.4975901629698244e-20

R2_184 V2 V184 71135.67035543828
L2_184 V2 V184 -1.6726945523115066e-11
C2_184 V2 V184 2.403117355618153e-22

R2_185 V2 V185 -4163.083311440859
L2_185 V2 V185 2.0052086403859095e-11
C2_185 V2 V185 4.10419367534386e-20

R2_186 V2 V186 -15731.709020896751
L2_186 V2 V186 4.057485459273943e-12
C2_186 V2 V186 -5.6046428566785564e-21

R2_187 V2 V187 -8962.071230772295
L2_187 V2 V187 1.76999530552079e-12
C2_187 V2 V187 -2.1895808885928873e-19

R2_188 V2 V188 -4459.578115189731
L2_188 V2 V188 1.6185349289975547e-12
C2_188 V2 V188 -1.90345545628531e-19

R2_189 V2 V189 4053.918683598157
L2_189 V2 V189 6.056601213972302e-12
C2_189 V2 V189 -2.145389354732236e-19

R2_190 V2 V190 5202.73273113374
L2_190 V2 V190 -2.4680697927892706e-12
C2_190 V2 V190 2.286222902363003e-19

R2_191 V2 V191 -5617.126891323262
L2_191 V2 V191 2.209543683629804e-12
C2_191 V2 V191 -2.0684864749899037e-19

R2_192 V2 V192 -32793.90417322505
L2_192 V2 V192 5.928100134320559e-12
C2_192 V2 V192 -1.3532004122079967e-19

R2_193 V2 V193 -75249.3622096184
L2_193 V2 V193 -4.351948294227661e-12
C2_193 V2 V193 1.389040293022488e-19

R2_194 V2 V194 -7737.2188050649
L2_194 V2 V194 8.536697163978945e-12
C2_194 V2 V194 1.8123014255677116e-20

R2_195 V2 V195 4950.692813748112
L2_195 V2 V195 -1.2658575597245892e-12
C2_195 V2 V195 3.631091936273778e-19

R2_196 V2 V196 4465.491186801925
L2_196 V2 V196 -1.114256818841078e-12
C2_196 V2 V196 3.45330452848742e-19

R2_197 V2 V197 -7423.553416508771
L2_197 V2 V197 -2.9809110830643335e-12
C2_197 V2 V197 1.395184219879356e-19

R2_198 V2 V198 -38762.89268056515
L2_198 V2 V198 5.8679099120951086e-12
C2_198 V2 V198 -4.4304722629049654e-20

R2_199 V2 V199 5623.710366045787
L2_199 V2 V199 -3.0502637066837277e-12
C2_199 V2 V199 1.6700151880325228e-19

R2_200 V2 V200 228095.5972051205
L2_200 V2 V200 -1.648505466853579e-11
C2_200 V2 V200 5.966577893355301e-20

R3_3 V3 0 2032.4413328891703
L3_3 V3 0 3.59471922475185e-12
C3_3 V3 0 7.524735765642459e-23

R3_4 V3 V4 201966.90739936352
L3_4 V3 V4 3.0992048699780595e-11
C3_4 V3 V4 1.8149349130428704e-20

R3_5 V3 V5 -27455.585552053348
L3_5 V3 V5 3.9191271473696735e-12
C3_5 V3 V5 -1.1250757388307525e-19

R3_6 V3 V6 -11223.157506870426
L3_6 V3 V6 2.4456978446843338e-12
C3_6 V3 V6 -2.8470546825135107e-19

R3_7 V3 V7 6384.468450470114
L3_7 V3 V7 -8.299311986236509e-13
C3_7 V3 V7 7.289119961669115e-19

R3_8 V3 V8 58787.259552178475
L3_8 V3 V8 -5.471528509412761e-12
C3_8 V3 V8 1.2069719435921783e-19

R3_9 V3 V9 -5005.483038989448
L3_9 V3 V9 -6.55072034426785e-11
C3_9 V3 V9 2.7980419439800075e-20

R3_10 V3 V10 -8702.126293811869
L3_10 V3 V10 -9.510759246889336e-12
C3_10 V3 V10 4.99072689952136e-20

R3_11 V3 V11 3042.9180451006746
L3_11 V3 V11 9.103436109991112e-12
C3_11 V3 V11 -5.596929079792798e-20

R3_12 V3 V12 83598.16421178271
L3_12 V3 V12 1.31165074540225e-11
C3_12 V3 V12 -8.035165274688772e-20

R3_13 V3 V13 16929.77815191842
L3_13 V3 V13 1.5272704361108016e-11
C3_13 V3 V13 -5.629911751446155e-20

R3_14 V3 V14 38004.79259285817
L3_14 V3 V14 -8.918707846085226e-12
C3_14 V3 V14 2.734761245159738e-20

R3_15 V3 V15 -5537.152495025052
L3_15 V3 V15 1.586706123025886e-12
C3_15 V3 V15 -3.1606366157521697e-19

R3_16 V3 V16 -28692.412451202097
L3_16 V3 V16 5.546295429562626e-12
C3_16 V3 V16 -9.217932669644556e-20

R3_17 V3 V17 22894.660805841264
L3_17 V3 V17 -9.715441888458007e-12
C3_17 V3 V17 4.1214876485684355e-20

R3_18 V3 V18 17535.703389724804
L3_18 V3 V18 2.5041967029004403e-11
C3_18 V3 V18 -1.2925971481825746e-20

R3_19 V3 V19 -7715.661863904799
L3_19 V3 V19 -7.932790662434664e-12
C3_19 V3 V19 2.056425404740497e-19

R3_20 V3 V20 -49363.30874200402
L3_20 V3 V20 -1.5196483326326285e-11
C3_20 V3 V20 8.377978957542967e-20

R3_21 V3 V21 5366.431281544783
L3_21 V3 V21 -2.992503843535926e-11
C3_21 V3 V21 -1.7345066869949998e-20

R3_22 V3 V22 11823.123526538806
L3_22 V3 V22 -2.8736045308366645e-11
C3_22 V3 V22 -5.2786098550311674e-21

R3_23 V3 V23 -5416.89076815947
L3_23 V3 V23 1.0710316696790393e-11
C3_23 V3 V23 -8.910187855265504e-20

R3_24 V3 V24 -133910.31931503286
L3_24 V3 V24 5.906680721030715e-11
C3_24 V3 V24 -8.800530198628105e-21

R3_25 V3 V25 -6955.085861870589
L3_25 V3 V25 1.1662583489798564e-11
C3_25 V3 V25 -3.3825907487393685e-20

R3_26 V3 V26 -21633.464907888363
L3_26 V3 V26 7.17745423775627e-12
C3_26 V3 V26 -3.0942231497591995e-20

R3_27 V3 V27 6017.0955364905
L3_27 V3 V27 -4.565103788667134e-12
C3_27 V3 V27 1.4461168388838366e-19

R3_28 V3 V28 36910.80389375844
L3_28 V3 V28 -3.207684155777911e-11
C3_28 V3 V28 8.836677332268699e-21

R3_29 V3 V29 -7271.793403116701
L3_29 V3 V29 -2.329614515056025e-11
C3_29 V3 V29 4.917086525693746e-20

R3_30 V3 V30 -14480.131471228275
L3_30 V3 V30 -7.834773309367615e-12
C3_30 V3 V30 6.905291452865234e-20

R3_31 V3 V31 4832.49158865956
L3_31 V3 V31 2.6235314946063906e-11
C3_31 V3 V31 -1.3619749227570738e-19

R3_32 V3 V32 29868.42626235365
L3_32 V3 V32 -2.079906966328041e-11
C3_32 V3 V32 -1.8055905921049333e-20

R3_33 V3 V33 -10754.390681235285
L3_33 V3 V33 8.915540982689948e-12
C3_33 V3 V33 -4.2248536899996835e-20

R3_34 V3 V34 448615.2375748865
L3_34 V3 V34 9.503913283052134e-12
C3_34 V3 V34 -2.0580169918407078e-20

R3_35 V3 V35 -15834.906754560317
L3_35 V3 V35 7.758510369033197e-12
C3_35 V3 V35 -5.8663215877987275e-21

R3_36 V3 V36 -35366.585808107804
L3_36 V3 V36 7.984378424054902e-12
C3_36 V3 V36 -5.926316147351952e-20

R3_37 V3 V37 14779.02190577215
L3_37 V3 V37 -3.537058446554427e-11
C3_37 V3 V37 1.9106980455464978e-20

R3_38 V3 V38 27821.119064137634
L3_38 V3 V38 8.713000210154781e-12
C3_38 V3 V38 -4.671717074354079e-20

R3_39 V3 V39 -5883.815910913484
L3_39 V3 V39 -4.602601906845165e-12
C3_39 V3 V39 1.7713789456804195e-19

R3_40 V3 V40 -18054.522951125047
L3_40 V3 V40 -1.644136222099588e-11
C3_40 V3 V40 8.844835875318687e-20

R3_41 V3 V41 43131.47008147383
L3_41 V3 V41 -8.165548148012566e-12
C3_41 V3 V41 2.6101457337882622e-20

R3_42 V3 V42 13772.049668752443
L3_42 V3 V42 -8.697323126330384e-12
C3_42 V3 V42 7.017622734593339e-20

R3_43 V3 V43 -18261.605810118195
L3_43 V3 V43 2.8580957663766713e-12
C3_43 V3 V43 -1.9019156118491594e-19

R3_44 V3 V44 38101.48154210958
L3_44 V3 V44 2.3371084556540847e-11
C3_44 V3 V44 -6.08991915044835e-20

R3_45 V3 V45 -17221.343897491486
L3_45 V3 V45 -2.3698948983492865e-11
C3_45 V3 V45 3.1046811892560756e-20

R3_46 V3 V46 -80315.15862520161
L3_46 V3 V46 -9.963136931602125e-12
C3_46 V3 V46 5.932392338148914e-20

R3_47 V3 V47 5458.42435194655
L3_47 V3 V47 -8.261787617872323e-12
C3_47 V3 V47 -2.0598962499369658e-20

R3_48 V3 V48 21568.084704918907
L3_48 V3 V48 -9.324060927168317e-12
C3_48 V3 V48 2.691064848915442e-20

R3_49 V3 V49 -10854.643192294861
L3_49 V3 V49 3.425539723682164e-11
C3_49 V3 V49 -1.2150579517261805e-21

R3_50 V3 V50 -55358.327308820444
L3_50 V3 V50 8.065866633182305e-12
C3_50 V3 V50 -3.5692046793643604e-20

R3_51 V3 V51 9566.7910874311
L3_51 V3 V51 -3.3305630356257287e-12
C3_51 V3 V51 1.7293233743933996e-19

R3_52 V3 V52 85104.05680702823
L3_52 V3 V52 -3.074020165975257e-10
C3_52 V3 V52 7.25500885493643e-21

R3_53 V3 V53 -40828.299486919874
L3_53 V3 V53 7.016504441497956e-12
C3_53 V3 V53 -4.975478242631569e-20

R3_54 V3 V54 52919.71960255766
L3_54 V3 V54 6.66613944876591e-12
C3_54 V3 V54 -4.7189638138247926e-20

R3_55 V3 V55 -16265.967714922417
L3_55 V3 V55 6.730189273858541e-12
C3_55 V3 V55 -6.963586747089595e-20

R3_56 V3 V56 -30915.65249914666
L3_56 V3 V56 6.1527689973572315e-12
C3_56 V3 V56 -6.177649741004513e-20

R3_57 V3 V57 566687.9532919312
L3_57 V3 V57 -6.596154618524757e-12
C3_57 V3 V57 8.776481707797408e-20

R3_58 V3 V58 17112.24565076454
L3_58 V3 V58 -5.461549364427663e-12
C3_58 V3 V58 7.406267509137047e-20

R3_59 V3 V59 -10679.866393399661
L3_59 V3 V59 3.0063092431134677e-12
C3_59 V3 V59 -8.493702950138699e-20

R3_60 V3 V60 894223.3084091007
L3_60 V3 V60 -2.1875004092179257e-11
C3_60 V3 V60 4.772003681539569e-20

R3_61 V3 V61 142305.49032411765
L3_61 V3 V61 -9.252648116532041e-11
C3_61 V3 V61 -5.9146421809800774e-21

R3_62 V3 V62 -70944.04758549956
L3_62 V3 V62 -1.9832473434519136e-11
C3_62 V3 V62 5.94567675986921e-20

R3_63 V3 V63 90470.84072229992
L3_63 V3 V63 -9.925400544276236e-12
C3_63 V3 V63 1.5812382843719834e-20

R3_64 V3 V64 74953.24569138573
L3_64 V3 V64 -1.1739389433595215e-11
C3_64 V3 V64 2.5294142263964296e-20

R3_65 V3 V65 -16635.570329211867
L3_65 V3 V65 -4.4075763503462434e-11
C3_65 V3 V65 1.0558122744729548e-20

R3_66 V3 V66 -91909.11859662014
L3_66 V3 V66 6.751023564886832e-12
C3_66 V3 V66 -5.684100620002619e-20

R3_67 V3 V67 10020.718687177296
L3_67 V3 V67 -3.758613174978529e-12
C3_67 V3 V67 1.4629047273701677e-19

R3_68 V3 V68 27059.58924696328
L3_68 V3 V68 -3.2711474731345343e-10
C3_68 V3 V68 -8.98361741874395e-21

R3_69 V3 V69 -33958.83484368487
L3_69 V3 V69 5.830490991858711e-12
C3_69 V3 V69 -7.837127347523559e-20

R3_70 V3 V70 -40802.16391920998
L3_70 V3 V70 1.7802511289241076e-11
C3_70 V3 V70 -5.622191438257881e-20

R3_71 V3 V71 8690.29842724036
L3_71 V3 V71 2.1547285016516334e-11
C3_71 V3 V71 -2.5941319748755564e-20

R3_72 V3 V72 29154.226725676017
L3_72 V3 V72 1.0691588206546484e-10
C3_72 V3 V72 -6.907999016013318e-21

R3_73 V3 V73 67488.83974677422
L3_73 V3 V73 -1.2181277979844755e-11
C3_73 V3 V73 7.750714653696257e-20

R3_74 V3 V74 25709.187519804957
L3_74 V3 V74 -4.333985433640615e-12
C3_74 V3 V74 1.356316303812862e-19

R3_75 V3 V75 -6122.401309986687
L3_75 V3 V75 2.455610128337995e-12
C3_75 V3 V75 -2.2070121975843655e-19

R3_76 V3 V76 -16875.228409941075
L3_76 V3 V76 1.2485768376193747e-11
C3_76 V3 V76 -3.0669455135333097e-20

R3_77 V3 V77 -70098.2493606329
L3_77 V3 V77 -8.263813434784851e-12
C3_77 V3 V77 4.4842284864934313e-20

R3_78 V3 V78 -47063.611015287584
L3_78 V3 V78 5.569942302050701e-12
C3_78 V3 V78 -1.6905801253992162e-19

R3_79 V3 V79 -16413.762512103385
L3_79 V3 V79 -3.126553221890031e-12
C3_79 V3 V79 1.7796593205047561e-19

R3_80 V3 V80 -26964.01080730482
L3_80 V3 V80 -2.6012821834970605e-11
C3_80 V3 V80 -1.0223325047793273e-20

R3_81 V3 V81 -7181.275994238132
L3_81 V3 V81 1.0005147432565012e-11
C3_81 V3 V81 -8.838072939729823e-20

R3_82 V3 V82 -118490.79781521947
L3_82 V3 V82 -8.498214362472114e-11
C3_82 V3 V82 3.776844462244833e-20

R3_83 V3 V83 9839.223889061259
L3_83 V3 V83 -7.859392468479715e-12
C3_83 V3 V83 2.765163718783385e-20

R3_84 V3 V84 15875.145415866913
L3_84 V3 V84 -8.074597916372566e-12
C3_84 V3 V84 3.960332425243503e-20

R3_85 V3 V85 44639.497513149014
L3_85 V3 V85 -6.974603176255823e-12
C3_85 V3 V85 6.108142876601744e-20

R3_86 V3 V86 10375.70002860382
L3_86 V3 V86 -3.516524888026007e-12
C3_86 V3 V86 1.6617502664906243e-19

R3_87 V3 V87 16170.382110674609
L3_87 V3 V87 2.077884864391117e-12
C3_87 V3 V87 -2.8054354234114494e-19

R3_88 V3 V88 42140.594268989546
L3_88 V3 V88 1.0274211120444877e-11
C3_88 V3 V88 -7.105795426765541e-20

R3_89 V3 V89 -89296.17792830674
L3_89 V3 V89 6.4465276568841095e-12
C3_89 V3 V89 -6.426185245074015e-20

R3_90 V3 V90 -24740.43699478191
L3_90 V3 V90 2.213867253354833e-12
C3_90 V3 V90 -2.2394630350539456e-19

R3_91 V3 V91 11274.21702191645
L3_91 V3 V91 -1.283914121897564e-12
C3_91 V3 V91 4.333691787192729e-19

R3_92 V3 V92 68572.1279874129
L3_92 V3 V92 -1.5702982332645414e-11
C3_92 V3 V92 3.223900756382418e-20

R3_93 V3 V93 -16796.174483158495
L3_93 V3 V93 1.1594477599291982e-11
C3_93 V3 V93 -4.464198608022597e-20

R3_94 V3 V94 -38018.28064830274
L3_94 V3 V94 1.5245595403856836e-11
C3_94 V3 V94 3.389178497263714e-21

R3_95 V3 V95 -4101.630222241863
L3_95 V3 V95 6.088966843068531e-12
C3_95 V3 V95 2.0163229715062624e-20

R3_96 V3 V96 -11243.2335115702
L3_96 V3 V96 1.0341396099862507e-10
C3_96 V3 V96 4.2874294022535285e-20

R3_97 V3 V97 -14865.986678371817
L3_97 V3 V97 -3.059934181641365e-12
C3_97 V3 V97 2.3331490144762747e-19

R3_98 V3 V98 13329.070337588284
L3_98 V3 V98 -2.6559218670886852e-12
C3_98 V3 V98 1.8358538023316103e-19

R3_99 V3 V99 4943.066926494684
L3_99 V3 V99 1.359107117831408e-12
C3_99 V3 V99 -4.758510752486043e-19

R3_100 V3 V100 12161.123811579959
L3_100 V3 V100 1.1675230473615806e-11
C3_100 V3 V100 -8.924925973526128e-20

R3_101 V3 V101 40278.470003087175
L3_101 V3 V101 6.342990585257383e-12
C3_101 V3 V101 -1.0642878211465977e-19

R3_102 V3 V102 33201.57459581763
L3_102 V3 V102 1.9713202759230258e-11
C3_102 V3 V102 -4.0325042068391034e-20

R3_103 V3 V103 36675.78474934378
L3_103 V3 V103 -1.6643085578369569e-12
C3_103 V3 V103 3.276074257435251e-19

R3_104 V3 V104 19708.705825656518
L3_104 V3 V104 -6.533592554097929e-12
C3_104 V3 V104 7.223812876688118e-20

R3_105 V3 V105 -10714.151452294285
L3_105 V3 V105 8.990717925651445e-12
C3_105 V3 V105 -8.012866023045518e-20

R3_106 V3 V106 -28945.76416980092
L3_106 V3 V106 2.5858727356702734e-12
C3_106 V3 V106 -2.3482087414659253e-19

R3_107 V3 V107 -29822.450877066753
L3_107 V3 V107 -1.8031472955804087e-11
C3_107 V3 V107 8.005974134374205e-20

R3_108 V3 V108 -63319.20918753655
L3_108 V3 V108 1.1543023132241856e-11
C3_108 V3 V108 -2.1764641327441446e-20

R3_109 V3 V109 27145.319545169532
L3_109 V3 V109 -7.308268812538169e-12
C3_109 V3 V109 1.325388411042907e-19

R3_110 V3 V110 -126054.07343423217
L3_110 V3 V110 -5.051731961986477e-12
C3_110 V3 V110 1.0987438690169035e-19

R3_111 V3 V111 4082.786316086001
L3_111 V3 V111 1.4639571338673184e-11
C3_111 V3 V111 -4.156650053130947e-20

R3_112 V3 V112 15730.922102570821
L3_112 V3 V112 1.3955392386815569e-11
C3_112 V3 V112 -5.175130767893702e-20

R3_113 V3 V113 -15355.647980582607
L3_113 V3 V113 -1.6990660348689383e-10
C3_113 V3 V113 -3.9062920666307794e-21

R3_114 V3 V114 39487.298752752155
L3_114 V3 V114 -2.806126565078695e-12
C3_114 V3 V114 2.1292609593159371e-19

R3_115 V3 V115 -4445.029080674132
L3_115 V3 V115 2.5322205366752244e-12
C3_115 V3 V115 -5.568554552013587e-20

R3_116 V3 V116 -13341.209172353203
L3_116 V3 V116 -1.6334622893035734e-11
C3_116 V3 V116 8.267809741229502e-20

R3_117 V3 V117 -9475.7702880711
L3_117 V3 V117 1.2206505202213772e-11
C3_117 V3 V117 -1.1173099664022596e-20

R3_118 V3 V118 -113338.11326791723
L3_118 V3 V118 2.853388821745045e-12
C3_118 V3 V118 -2.2455521954815563e-19

R3_119 V3 V119 6985.765412599712
L3_119 V3 V119 5.0461011723905344e-11
C3_119 V3 V119 -6.628109991176753e-20

R3_120 V3 V120 14624.21362307079
L3_120 V3 V120 8.604067169564878e-12
C3_120 V3 V120 -9.600743978302591e-20

R3_121 V3 V121 25129.348845856675
L3_121 V3 V121 -1.853170464242619e-11
C3_121 V3 V121 3.2705136476824645e-20

R3_122 V3 V122 208191.75600522198
L3_122 V3 V122 2.0317121714946055e-11
C3_122 V3 V122 -3.99683204067271e-20

R3_123 V3 V123 6885.240894116322
L3_123 V3 V123 -1.4304889668812981e-12
C3_123 V3 V123 3.593045820905113e-19

R3_124 V3 V124 20393.55063033307
L3_124 V3 V124 -7.931323107837271e-12
C3_124 V3 V124 4.5023192140224105e-20

R3_125 V3 V125 48293.49228076062
L3_125 V3 V125 3.477396326502524e-11
C3_125 V3 V125 -6.281926166158035e-20

R3_126 V3 V126 29547.20412038366
L3_126 V3 V126 -2.5096124739497242e-12
C3_126 V3 V126 1.7930271640076943e-19

R3_127 V3 V127 -4725.417723732314
L3_127 V3 V127 1.752537443432126e-12
C3_127 V3 V127 -2.6622063932386916e-19

R3_128 V3 V128 -12047.043392214504
L3_128 V3 V128 -1.7040046660237704e-11
C3_128 V3 V128 8.148393362783e-20

R3_129 V3 V129 -7669.137281762642
L3_129 V3 V129 3.3763725433302557e-11
C3_129 V3 V129 4.0708811790991675e-20

R3_130 V3 V130 -14690.124847991661
L3_130 V3 V130 1.478779323734588e-11
C3_130 V3 V130 -5.1335844300858404e-20

R3_131 V3 V131 16031.664602998002
L3_131 V3 V131 -4.1187250627190614e-11
C3_131 V3 V131 8.255391934119031e-24

R3_132 V3 V132 18909.329396195342
L3_132 V3 V132 3.916587991701988e-12
C3_132 V3 V132 -1.8593718578448778e-19

R3_133 V3 V133 -1885438.2629821193
L3_133 V3 V133 -3.083076644698874e-11
C3_133 V3 V133 2.569475206227079e-20

R3_134 V3 V134 -18394.74936806133
L3_134 V3 V134 4.285214903851032e-12
C3_134 V3 V134 -1.6388122983972042e-19

R3_135 V3 V135 7090.868665269951
L3_135 V3 V135 -1.1429094647145284e-12
C3_135 V3 V135 5.143837656105429e-19

R3_136 V3 V136 68240.68094466394
L3_136 V3 V136 -1.765900273957191e-11
C3_136 V3 V136 2.0085366045518018e-20

R3_137 V3 V137 24322.319338626912
L3_137 V3 V137 -5.042616577146429e-12
C3_137 V3 V137 5.930479674559495e-20

R3_138 V3 V138 -93248.29761775372
L3_138 V3 V138 -2.8134955487808e-12
C3_138 V3 V138 1.8572303629759771e-19

R3_139 V3 V139 -6693.620600011584
L3_139 V3 V139 8.109411021218035e-13
C3_139 V3 V139 -6.9713482191096e-19

R3_140 V3 V140 -12857.347767623367
L3_140 V3 V140 -7.604389343715608e-11
C3_140 V3 V140 1.479568366239625e-20

R3_141 V3 V141 7247.787961118629
L3_141 V3 V141 4.474943825075772e-11
C3_141 V3 V141 -3.791376520761248e-20

R3_142 V3 V142 7373.141600845276
L3_142 V3 V142 -7.605385083217483e-12
C3_142 V3 V142 5.196682774709222e-20

R3_143 V3 V143 6246.5829053005855
L3_143 V3 V143 -7.305751954334546e-12
C3_143 V3 V143 1.4947847791531253e-19

R3_144 V3 V144 7136.915797787365
L3_144 V3 V144 6.536608971549389e-11
C3_144 V3 V144 -2.3710386325738568e-20

R3_145 V3 V145 -3742.3103127738846
L3_145 V3 V145 5.6695866835658256e-12
C3_145 V3 V145 -4.445480557337201e-20

R3_146 V3 V146 -9366.266635170043
L3_146 V3 V146 2.9226467120885984e-12
C3_146 V3 V146 -1.1053445920520067e-19

R3_147 V3 V147 -2325.1483576447986
L3_147 V3 V147 -1.4943378268311024e-12
C3_147 V3 V147 2.9382644517332015e-19

R3_148 V3 V148 -4184.258555238209
L3_148 V3 V148 1.2723602507206486e-11
C3_148 V3 V148 -1.3417799815747383e-20

R3_149 V3 V149 6099.275241557233
L3_149 V3 V149 1.3859546193608257e-11
C3_149 V3 V149 1.255404866060082e-20

R3_150 V3 V150 17469.09094806154
L3_150 V3 V150 -3.1535284990734395e-11
C3_150 V3 V150 -6.05074674667316e-20

R3_151 V3 V151 1265.6225846406544
L3_151 V3 V151 -2.1398559742005448e-10
C3_151 V3 V151 -3.555950917686572e-20

R3_152 V3 V152 4022.5076036959454
L3_152 V3 V152 -1.1517518974431692e-11
C3_152 V3 V152 4.702752187562737e-20

R3_153 V3 V153 -11504.60488057064
L3_153 V3 V153 -4.9003337944830205e-12
C3_153 V3 V153 1.2262572522808173e-19

R3_154 V3 V154 7766.152140351076
L3_154 V3 V154 -7.42542336111247e-12
C3_154 V3 V154 1.457269665183285e-19

R3_155 V3 V155 -714.3825633073365
L3_155 V3 V155 1.2047249659854378e-12
C3_155 V3 V155 -4.4840596953591075e-19

R3_156 V3 V156 -11394.796611604292
L3_156 V3 V156 -6.842334564596547e-11
C3_156 V3 V156 3.1672531894099687e-20

R3_157 V3 V157 -20369.39923745928
L3_157 V3 V157 -9.457355501074633e-12
C3_157 V3 V157 -3.860693487903924e-20

R3_158 V3 V158 35452.5539603699
L3_158 V3 V158 -2.217676259607902e-11
C3_158 V3 V158 -6.222893472453607e-20

R3_159 V3 V159 2617.770925928865
L3_159 V3 V159 -2.9258389052137575e-12
C3_159 V3 V159 3.732278526487069e-19

R3_160 V3 V160 -25364.105885688663
L3_160 V3 V160 8.183348749182695e-09
C3_160 V3 V160 -2.1029134995370652e-20

R3_161 V3 V161 -17351.826914876747
L3_161 V3 V161 3.7246889989973095e-12
C3_161 V3 V161 -1.6303014931815922e-19

R3_162 V3 V162 -34912.716336104095
L3_162 V3 V162 5.203966278647574e-12
C3_162 V3 V162 -3.3728992374089264e-20

R3_163 V3 V163 3180.3074198008458
L3_163 V3 V163 -3.874732540840109e-12
C3_163 V3 V163 -2.0323427908137801e-19

R3_164 V3 V164 5423.017679866768
L3_164 V3 V164 -2.845722994112742e-11
C3_164 V3 V164 -3.9533793730051514e-20

R3_165 V3 V165 -12695.98025478759
L3_165 V3 V165 -5.4387961597583175e-12
C3_165 V3 V165 1.3141042194564253e-19

R3_166 V3 V166 -67793.8997239325
L3_166 V3 V166 -4.4908758670226933e-11
C3_166 V3 V166 2.4714501549258005e-20

R3_167 V3 V167 6697.059635647822
L3_167 V3 V167 3.178025839461455e-12
C3_167 V3 V167 -6.415123781556072e-21

R3_168 V3 V168 -9210.462917137986
L3_168 V3 V168 5.666342686056688e-12
C3_168 V3 V168 -1.165955384583233e-19

R3_169 V3 V169 12970.93792958208
L3_169 V3 V169 -4.268812380641486e-12
C3_169 V3 V169 1.673129360640384e-19

R3_170 V3 V170 12630.915311846418
L3_170 V3 V170 -2.1762183672145638e-11
C3_170 V3 V170 -2.058787829262793e-22

R3_171 V3 V171 -1629.7272743059611
L3_171 V3 V171 -6.587725731836034e-12
C3_171 V3 V171 1.043011031017809e-19

R3_172 V3 V172 -8352.945060594857
L3_172 V3 V172 -6.876202347866054e-12
C3_172 V3 V172 1.1568829291165852e-19

R3_173 V3 V173 -7430.955825498074
L3_173 V3 V173 3.1479577627996056e-12
C3_173 V3 V173 -1.255161740647934e-19

R3_174 V3 V174 -60840.2135104605
L3_174 V3 V174 -1.1524235525311946e-11
C3_174 V3 V174 6.367154745910394e-20

R3_175 V3 V175 2839.5197412241223
L3_175 V3 V175 1.0892686544933333e-11
C3_175 V3 V175 -1.4316042734672714e-19

R3_176 V3 V176 19516.168154903873
L3_176 V3 V176 -7.581028301276645e-12
C3_176 V3 V176 4.917645762649168e-20

R3_177 V3 V177 8107.189670317562
L3_177 V3 V177 -5.8628090714896765e-12
C3_177 V3 V177 2.174279471983013e-20

R3_178 V3 V178 -51386.62689750189
L3_178 V3 V178 5.441882690684214e-11
C3_178 V3 V178 -4.2072796189178843e-20

R3_179 V3 V179 -3424.4057238789946
L3_179 V3 V179 7.319759268817964e-11
C3_179 V3 V179 1.5790404214589493e-20

R3_180 V3 V180 15540.393978564665
L3_180 V3 V180 8.010627719721828e-12
C3_180 V3 V180 -5.657980278998892e-20

R3_181 V3 V181 -143320.90872846733
L3_181 V3 V181 1.0237859270944234e-11
C3_181 V3 V181 -4.4183848032149383e-20

R3_182 V3 V182 -7243.641986583248
L3_182 V3 V182 -2.659214527028543e-10
C3_182 V3 V182 1.0968000300166554e-20

R3_183 V3 V183 3995.7442147648335
L3_183 V3 V183 -7.187043097698895e-12
C3_183 V3 V183 -5.067248331161318e-21

R3_184 V3 V184 -70744.03142129577
L3_184 V3 V184 -1.0611401235590062e-11
C3_184 V3 V184 1.6503385626561047e-20

R3_185 V3 V185 -5702.527818389049
L3_185 V3 V185 5.3028009520160404e-12
C3_185 V3 V185 8.737104962709772e-21

R3_186 V3 V186 10239.672914233985
L3_186 V3 V186 -8.473948022064392e-12
C3_186 V3 V186 5.017756437930511e-20

R3_187 V3 V187 -26730.537974974417
L3_187 V3 V187 2.390540377287253e-12
C3_187 V3 V187 -1.302475553334801e-19

R3_188 V3 V188 -5685.97614739234
L3_188 V3 V188 5.1149860901926526e-12
C3_188 V3 V188 -7.156896207800987e-20

R3_189 V3 V189 4039.9715196490743
L3_189 V3 V189 -3.5022229122918203e-12
C3_189 V3 V189 1.0703612297514221e-19

R3_190 V3 V190 201032.45462875077
L3_190 V3 V190 1.1624040554602845e-11
C3_190 V3 V190 -4.9949336859810766e-20

R3_191 V3 V191 -9440.209427209167
L3_191 V3 V191 -4.66114653160272e-12
C3_191 V3 V191 2.772679885156815e-19

R3_192 V3 V192 52535.58480243262
L3_192 V3 V192 -3.897751267998178e-11
C3_192 V3 V192 1.3543480444627122e-19

R3_193 V3 V193 266046.8270283492
L3_193 V3 V193 9.397234406576433e-11
C3_193 V3 V193 -1.0626855005912874e-20

R3_194 V3 V194 -18988.49452949953
L3_194 V3 V194 -3.3365303290864147e-12
C3_194 V3 V194 1.5084111107587885e-19

R3_195 V3 V195 35135.64492269495
L3_195 V3 V195 3.962460187843205e-12
C3_195 V3 V195 -3.8414090349486203e-19

R3_196 V3 V196 3540.568703492625
L3_196 V3 V196 -4.069793959800872e-12
C3_196 V3 V196 4.903415710339761e-20

R3_197 V3 V197 -16430.272771344513
L3_197 V3 V197 5.4377145452389456e-12
C3_197 V3 V197 -8.461875542105807e-20

R3_198 V3 V198 6485.657416941937
L3_198 V3 V198 2.164921957479479e-11
C3_198 V3 V198 -8.134231436058414e-21

R3_199 V3 V199 40953.85653649069
L3_199 V3 V199 7.767594125484675e-12
C3_199 V3 V199 -7.246659570888423e-20

R3_200 V3 V200 -29081.152112774736
L3_200 V3 V200 3.981493335177442e-12
C3_200 V3 V200 -1.5542878464752022e-19

R4_4 V4 0 -1887.8044692365597
L4_4 V4 0 5.966161407657952e-13
C4_4 V4 0 -1.1951049811262118e-18

R4_5 V4 V5 -31365.113714200652
L4_5 V4 V5 5.55159497856526e-12
C4_5 V4 V5 -9.66728224265108e-20

R4_6 V4 V6 -12424.661985831903
L4_6 V4 V6 3.0235289325670397e-12
C4_6 V4 V6 -2.5137293684289465e-19

R4_7 V4 V7 -10327.316998841572
L4_7 V4 V7 9.137638747495214e-12
C4_7 V4 V7 -2.9426182686258877e-19

R4_8 V4 V8 4088.28952531268
L4_8 V4 V8 -7.731300867648592e-13
C4_8 V4 V8 1.0219480778553813e-18

R4_9 V4 V9 -6169.739964106783
L4_9 V4 V9 2.351475338727511e-10
C4_9 V4 V9 6.017574186418295e-21

R4_10 V4 V10 -9661.552034448507
L4_10 V4 V10 -1.065656474618262e-11
C4_10 V4 V10 4.617643841813832e-20

R4_11 V4 V11 -13931.09674837413
L4_11 V4 V11 2.700818781252762e-11
C4_11 V4 V11 7.224895138034585e-20

R4_12 V4 V12 3011.816620734595
L4_12 V4 V12 1.4266320003770596e-11
C4_12 V4 V12 -8.029533821923959e-20

R4_13 V4 V13 24242.660574012792
L4_13 V4 V13 1.341782512278175e-11
C4_13 V4 V13 -7.186402702163051e-20

R4_14 V4 V14 66549.20280939255
L4_14 V4 V14 -2.557731739470828e-11
C4_14 V4 V14 -3.0579821531905395e-20

R4_15 V4 V15 -111048.0861316932
L4_15 V4 V15 -8.977182287692465e-12
C4_15 V4 V15 -5.932559526766695e-20

R4_16 V4 V16 -5491.479542523907
L4_16 V4 V16 1.2342549155399818e-12
C4_16 V4 V16 -3.1703750460880237e-19

R4_17 V4 V17 26189.24294113037
L4_17 V4 V17 -1.0605426889093647e-11
C4_17 V4 V17 5.757393603449417e-20

R4_18 V4 V18 18201.265442084597
L4_18 V4 V18 7.545143292829244e-11
C4_18 V4 V18 3.5366092523650937e-20

R4_19 V4 V19 18454.314326400592
L4_19 V4 V19 -4.7813549743767514e-11
C4_19 V4 V19 2.785134665842884e-20

R4_20 V4 V20 -7365.224563370271
L4_20 V4 V20 -6.842379640387545e-12
C4_20 V4 V20 2.758744669995666e-19

R4_21 V4 V21 6942.139283135855
L4_21 V4 V21 -6.276228685424044e-11
C4_21 V4 V21 -4.019167272662809e-21

R4_22 V4 V22 12797.970134519122
L4_22 V4 V22 -5.378107802082811e-11
C4_22 V4 V22 -1.274668204311781e-20

R4_23 V4 V23 19834.578420165843
L4_23 V4 V23 -7.844696330038708e-11
C4_23 V4 V23 -3.541928219558613e-20

R4_24 V4 V24 -5592.619429460605
L4_24 V4 V24 6.2628894562878945e-12
C4_24 V4 V24 -1.0054822613601056e-19

R4_25 V4 V25 -9361.172945437185
L4_25 V4 V25 1.8300129918787073e-11
C4_25 V4 V25 -4.681077632777435e-21

R4_26 V4 V26 -27510.20974602085
L4_26 V4 V26 1.2850639184113827e-11
C4_26 V4 V26 3.7992764356305087e-20

R4_27 V4 V27 -130891.22004357292
L4_27 V4 V27 9.866328419255717e-12
C4_27 V4 V27 5.2441228060097377e-20

R4_28 V4 V28 5092.623069542736
L4_28 V4 V28 -2.510815415825953e-12
C4_28 V4 V28 2.2292065461280886e-19

R4_29 V4 V29 -9804.068709478554
L4_29 V4 V29 -1.6195916412542867e-11
C4_29 V4 V29 4.8204208457995644e-20

R4_30 V4 V30 -16421.167996748045
L4_30 V4 V30 -8.130738649594376e-12
C4_30 V4 V30 5.396615502756135e-20

R4_31 V4 V31 -34435.7568616604
L4_31 V4 V31 -2.0479636580535038e-11
C4_31 V4 V31 9.54795209765125e-20

R4_32 V4 V32 5529.164858972244
L4_32 V4 V32 7.014867990412687e-11
C4_32 V4 V32 -2.701845341434141e-19

R4_33 V4 V33 -11872.741024330995
L4_33 V4 V33 9.451189971136262e-12
C4_33 V4 V33 -1.9528261781955362e-20

R4_34 V4 V34 -63554.87259795894
L4_34 V4 V34 1.1973171431493259e-11
C4_34 V4 V34 1.7357847773459362e-20

R4_35 V4 V35 30337.27915799301
L4_35 V4 V35 7.483132411264749e-12
C4_35 V4 V35 2.3072067238590346e-20

R4_36 V4 V36 -6226.740450839613
L4_36 V4 V36 5.372766170720251e-12
C4_36 V4 V36 -1.6777711929357332e-19

R4_37 V4 V37 23488.369097362738
L4_37 V4 V37 2.4644529414244494e-10
C4_37 V4 V37 5.2459343390648095e-21

R4_38 V4 V38 56682.43586907825
L4_38 V4 V38 8.444747704764767e-12
C4_38 V4 V38 -5.3912819192779915e-20

R4_39 V4 V39 34087.78326613935
L4_39 V4 V39 1.1456372375393667e-11
C4_39 V4 V39 -2.454316325349427e-20

R4_40 V4 V40 -5025.229563999355
L4_40 V4 V40 -4.4059488040223975e-12
C4_40 V4 V40 1.345139450220529e-19

R4_41 V4 V41 38065.42367893461
L4_41 V4 V41 -7.212320599198741e-12
C4_41 V4 V41 5.240578582053717e-20

R4_42 V4 V42 14684.52157664822
L4_42 V4 V42 -7.371929645516434e-12
C4_42 V4 V42 1.1262277060283378e-19

R4_43 V4 V43 12167.805082233634
L4_43 V4 V43 -9.82979803268963e-12
C4_43 V4 V43 8.926426264748659e-20

R4_44 V4 V44 -15763.829611252186
L4_44 V4 V44 2.8952369602623597e-12
C4_44 V4 V44 -2.244704079509546e-19

R4_45 V4 V45 -31372.99761930796
L4_45 V4 V45 -1.3958617446853009e-11
C4_45 V4 V45 4.355591051860409e-20

R4_46 V4 V46 106882.29605181106
L4_46 V4 V46 -7.608216394013747e-12
C4_46 V4 V46 7.400294262758766e-20

R4_47 V4 V47 634224.0705768742
L4_47 V4 V47 -1.1473307669199206e-11
C4_47 V4 V47 6.776462417862029e-20

R4_48 V4 V48 3734.073165315951
L4_48 V4 V48 -3.524060245367602e-12
C4_48 V4 V48 5.164761552495277e-20

R4_49 V4 V49 -12978.840262931357
L4_49 V4 V49 3.5449149861775274e-11
C4_49 V4 V49 2.440202225987854e-20

R4_50 V4 V50 -38962.18479381551
L4_50 V4 V50 9.624402251209882e-12
C4_50 V4 V50 5.430633450848656e-22

R4_51 V4 V51 172603.0663316854
L4_51 V4 V51 4.476298373787032e-12
C4_51 V4 V51 -1.2789761747751316e-20

R4_52 V4 V52 65268.34448453494
L4_52 V4 V52 -4.620485069298119e-12
C4_52 V4 V52 3.8471974172946655e-20

R4_53 V4 V53 -36667.296115027326
L4_53 V4 V53 8.281855441604594e-12
C4_53 V4 V53 -3.570742749391102e-20

R4_54 V4 V54 -109647.82074443215
L4_54 V4 V54 6.958515368640613e-12
C4_54 V4 V54 -4.4283510332539924e-20

R4_55 V4 V55 55536.28961741691
L4_55 V4 V55 1.0584483508919326e-11
C4_55 V4 V55 -1.084483279718076e-20

R4_56 V4 V56 -6408.992722815009
L4_56 V4 V56 5.281089000070453e-12
C4_56 V4 V56 -1.9214687321256763e-19

R4_57 V4 V57 326005.9628179364
L4_57 V4 V57 -7.197968558940617e-12
C4_57 V4 V57 1.0429860036613817e-19

R4_58 V4 V58 16178.010384187719
L4_58 V4 V58 -5.196021672111841e-12
C4_58 V4 V58 1.0020805283117524e-19

R4_59 V4 V59 14140.774225592806
L4_59 V4 V59 -4.3518182363853456e-12
C4_59 V4 V59 1.694562225658168e-19

R4_60 V4 V60 -8030.07231709817
L4_60 V4 V60 2.7566958426449146e-12
C4_60 V4 V60 -1.2701365163936592e-19

R4_61 V4 V61 90661.21955484766
L4_61 V4 V61 -3.681948364787145e-11
C4_61 V4 V61 -1.4110911344520668e-20

R4_62 V4 V62 -319924.4030045426
L4_62 V4 V62 -1.4932316603718435e-11
C4_62 V4 V62 6.329330855933506e-20

R4_63 V4 V63 153901.19056380625
L4_63 V4 V63 2.6066823148154066e-11
C4_63 V4 V63 -1.7253183668828885e-20

R4_64 V4 V64 26068.557361367228
L4_64 V4 V64 -3.968804622194063e-12
C4_64 V4 V64 1.827544258009015e-20

R4_65 V4 V65 -26918.02952978507
L4_65 V4 V65 -2.3649138300970006e-11
C4_65 V4 V65 4.0826430886928004e-20

R4_66 V4 V66 -66936.02044092858
L4_66 V4 V66 8.522599665020986e-12
C4_66 V4 V66 -1.657387765147654e-20

R4_67 V4 V67 -39712.05960289135
L4_67 V4 V67 4.416439477809547e-12
C4_67 V4 V67 -7.556118444373287e-20

R4_68 V4 V68 8306.697590429721
L4_68 V4 V68 -2.6188945066923727e-12
C4_68 V4 V68 1.5168093838513494e-19

R4_69 V4 V69 -19727.772991869533
L4_69 V4 V69 5.805365165971182e-12
C4_69 V4 V69 -9.785794313696872e-20

R4_70 V4 V70 -26494.10232972323
L4_70 V4 V70 1.3991477379430142e-11
C4_70 V4 V70 -9.001868316118268e-20

R4_71 V4 V71 -29254.65018520357
L4_71 V4 V71 -7.928358991841513e-12
C4_71 V4 V71 1.2555392182870642e-20

R4_72 V4 V72 10534.638886620329
L4_72 V4 V72 4.590091283060791e-12
C4_72 V4 V72 -9.76698919147341e-20

R4_73 V4 V73 320789.1419926896
L4_73 V4 V73 -1.771018788589498e-11
C4_73 V4 V73 8.567754591901119e-20

R4_74 V4 V74 37217.45482424195
L4_74 V4 V74 -5.379380614964624e-12
C4_74 V4 V74 1.2199530400278922e-19

R4_75 V4 V75 11791.882108306865
L4_75 V4 V75 -7.781173026983396e-12
C4_75 V4 V75 1.3677291577848797e-19

R4_76 V4 V76 -3944.640489866132
L4_76 V4 V76 1.8831389287837097e-12
C4_76 V4 V76 -2.9564110223946574e-19

R4_77 V4 V77 294386.70554528804
L4_77 V4 V77 -9.231613282733901e-12
C4_77 V4 V77 5.710303694884775e-20

R4_78 V4 V78 83399.11399012526
L4_78 V4 V78 8.132833616308815e-12
C4_78 V4 V78 -1.2996533783765697e-19

R4_79 V4 V79 -43582.280110022686
L4_79 V4 V79 4.269753086308812e-12
C4_79 V4 V79 -1.1735999640794816e-19

R4_80 V4 V80 254479.04162155784
L4_80 V4 V80 -2.108898938206755e-12
C4_80 V4 V80 2.3334761001894583e-19

R4_81 V4 V81 -15697.26331018714
L4_81 V4 V81 7.906945914008173e-11
C4_81 V4 V81 5.8671822271693605e-21

R4_82 V4 V82 -307256.93602201645
L4_82 V4 V82 -1.0416356149944156e-10
C4_82 V4 V82 5.512411845002549e-20

R4_83 V4 V83 15753.113995254465
L4_83 V4 V83 2.2032213354979615e-11
C4_83 V4 V83 8.954576736237794e-20

R4_84 V4 V84 8068.64853853335
L4_84 V4 V84 -3.5232413243942003e-12
C4_84 V4 V84 3.445262065090418e-20

R4_85 V4 V85 87924.38460865316
L4_85 V4 V85 -1.0102027459773908e-11
C4_85 V4 V85 2.7021553199994276e-20

R4_86 V4 V86 16356.022288388569
L4_86 V4 V86 -4.992889358676747e-12
C4_86 V4 V86 1.3843314160487107e-19

R4_87 V4 V87 -468562.5119857526
L4_87 V4 V87 -9.095595917556054e-12
C4_87 V4 V87 3.35530160512515e-20

R4_88 V4 V88 18319.19525706112
L4_88 V4 V88 1.5209385085987425e-12
C4_88 V4 V88 -3.1484896734324735e-19

R4_89 V4 V89 -30897.94520980814
L4_89 V4 V89 4.6712641767241275e-12
C4_89 V4 V89 -7.353167943331327e-20

R4_90 V4 V90 -38078.13556264281
L4_90 V4 V90 2.612099589722106e-12
C4_90 V4 V90 -1.3833029594108925e-19

R4_91 V4 V91 31204.925061445676
L4_91 V4 V91 5.067650889680147e-12
C4_91 V4 V91 -7.00768954671276e-20

R4_92 V4 V92 48146.76122774174
L4_92 V4 V92 -1.0965528638895886e-12
C4_92 V4 V92 3.578826684100865e-19

R4_93 V4 V93 -43191.42365918012
L4_93 V4 V93 1.7021137835034748e-11
C4_93 V4 V93 8.13034111973232e-21

R4_94 V4 V94 206332.26438673626
L4_94 V4 V94 2.992984629368574e-11
C4_94 V4 V94 4.290698437270913e-20

R4_95 V4 V95 59307.45594649868
L4_95 V4 V95 -1.3228915632187683e-11
C4_95 V4 V95 2.937474751724129e-20

R4_96 V4 V96 -3596.560544127848
L4_96 V4 V96 3.193716689235738e-12
C4_96 V4 V96 2.9661178800537837e-20

R4_97 V4 V97 -23275.424217386837
L4_97 V4 V97 -3.0930073121089956e-12
C4_97 V4 V97 2.5638749714799105e-19

R4_98 V4 V98 18792.23227997094
L4_98 V4 V98 -2.9336299490392776e-12
C4_98 V4 V98 1.5023705364268758e-19

R4_99 V4 V99 41505.41161711382
L4_99 V4 V99 1.3327763280077089e-11
C4_99 V4 V99 1.357479819769886e-19

R4_100 V4 V100 3675.7203347857053
L4_100 V4 V100 1.7904491101445525e-12
C4_100 V4 V100 -5.246750873118825e-19

R4_101 V4 V101 30031.819984205435
L4_101 V4 V101 6.267297857919195e-12
C4_101 V4 V101 -5.893288825138969e-20

R4_102 V4 V102 53215.354417153714
L4_102 V4 V102 1.185611674885671e-11
C4_102 V4 V102 -4.841910403832014e-20

R4_103 V4 V103 17251.430538166165
L4_103 V4 V103 1.1226229316870844e-11
C4_103 V4 V103 -3.686399845685568e-20

R4_104 V4 V104 43885.356316006946
L4_104 V4 V104 -1.4892458824556186e-12
C4_104 V4 V104 3.557694476270908e-19

R4_105 V4 V105 -11541.76276684621
L4_105 V4 V105 8.059186277179075e-12
C4_105 V4 V105 -6.658398461004117e-20

R4_106 V4 V106 -50875.156252138055
L4_106 V4 V106 4.5413554248924586e-12
C4_106 V4 V106 -1.4253343096427797e-19

R4_107 V4 V107 59323.72139550354
L4_107 V4 V107 -1.6471841168188368e-11
C4_107 V4 V107 -1.0072855519952082e-20

R4_108 V4 V108 -7333.059139777564
L4_108 V4 V108 2.889910857999611e-12
C4_108 V4 V108 -2.151322930328539e-21

R4_109 V4 V109 -776681.4508836707
L4_109 V4 V109 -7.458396498659548e-12
C4_109 V4 V109 1.5007115519638844e-19

R4_110 V4 V110 -22260.913554493134
L4_110 V4 V110 -2.1935844166366865e-11
C4_110 V4 V110 -3.325321346763533e-21

R4_111 V4 V111 -19121.381431911937
L4_111 V4 V111 2.2667399697520823e-11
C4_111 V4 V111 -7.672331959968702e-20

R4_112 V4 V112 3489.775465946198
L4_112 V4 V112 -2.534866166465864e-12
C4_112 V4 V112 1.9004747320819106e-19

R4_113 V4 V113 -41376.68240075761
L4_113 V4 V113 -1.689766321756252e-11
C4_113 V4 V113 -1.30603895766178e-20

R4_114 V4 V114 31167.440929928543
L4_114 V4 V114 -3.0591944717157094e-12
C4_114 V4 V114 1.465784189764803e-19

R4_115 V4 V115 -19175.6626502227
L4_115 V4 V115 -5.351708648499825e-12
C4_115 V4 V115 7.042532938739017e-20

R4_116 V4 V116 -5427.349361354814
L4_116 V4 V116 2.6827855190737578e-12
C4_116 V4 V116 -1.0798863458071765e-19

R4_117 V4 V117 -11509.14407179359
L4_117 V4 V117 1.2927763386165439e-11
C4_117 V4 V117 -3.140725670368566e-20

R4_118 V4 V118 107016.02429414626
L4_118 V4 V118 6.029501663581339e-12
C4_118 V4 V118 -1.2979565645490963e-19

R4_119 V4 V119 -77485.41818991219
L4_119 V4 V119 6.276620388087772e-12
C4_119 V4 V119 -1.4707735396298348e-19

R4_120 V4 V120 5829.345629259022
L4_120 V4 V120 3.2407448466933303e-12
C4_120 V4 V120 -3.233652084129345e-19

R4_121 V4 V121 -538603.8895600174
L4_121 V4 V121 -7.994591369250216e-11
C4_121 V4 V121 4.807881449318786e-20

R4_122 V4 V122 -28546.68493536298
L4_122 V4 V122 8.92063142286116e-12
C4_122 V4 V122 -1.0106553950415608e-19

R4_123 V4 V123 41105.3444613023
L4_123 V4 V123 9.417277867156208e-12
C4_123 V4 V123 -5.916737287122297e-20

R4_124 V4 V124 31204.324499651917
L4_124 V4 V124 -8.748406450041321e-13
C4_124 V4 V124 6.680104164593006e-19

R4_125 V4 V125 49400.054514200914
L4_125 V4 V125 -2.5713373530925863e-11
C4_125 V4 V125 -2.958097420523729e-20

R4_126 V4 V126 42733.08428095257
L4_126 V4 V126 -2.9865897019334655e-12
C4_126 V4 V126 7.854156151790715e-20

R4_127 V4 V127 -97057.1075104154
L4_127 V4 V127 -1.829483349043994e-12
C4_127 V4 V127 2.442146844877186e-19

R4_128 V4 V128 -4690.967146271931
L4_128 V4 V128 1.5563977304475088e-12
C4_128 V4 V128 -1.861163374809037e-19

R4_129 V4 V129 -9239.73395272697
L4_129 V4 V129 3.1970675476822974e-11
C4_129 V4 V129 3.970716714889849e-20

R4_130 V4 V130 -23941.074128425313
L4_130 V4 V130 1.655755379970198e-11
C4_130 V4 V130 -5.069043904379952e-20

R4_131 V4 V131 13535.65788359992
L4_131 V4 V131 2.6245562664308186e-12
C4_131 V4 V131 -1.9367608842476114e-19

R4_132 V4 V132 5684.183856347363
L4_132 V4 V132 7.415495447505452e-12
C4_132 V4 V132 -1.7219251298300803e-19

R4_133 V4 V133 49936.556691489954
L4_133 V4 V133 2.5481233989627227e-11
C4_133 V4 V133 -8.541799484944781e-20

R4_134 V4 V134 -35394.00140316522
L4_134 V4 V134 3.907328837777472e-12
C4_134 V4 V134 -2.6250562693045077e-19

R4_135 V4 V135 -7825.069333268542
L4_135 V4 V135 3.099215468635144e-12
C4_135 V4 V135 -2.717792921352088e-19

R4_136 V4 V136 9518.126339225879
L4_136 V4 V136 -9.999663139880413e-13
C4_136 V4 V136 5.832907509622428e-19

R4_137 V4 V137 -93765.16163683949
L4_137 V4 V137 -3.5640074998411543e-12
C4_137 V4 V137 1.101232015741371e-19

R4_138 V4 V138 -21930.33172720326
L4_138 V4 V138 -2.8473817885589598e-12
C4_138 V4 V138 1.9402416602886208e-19

R4_139 V4 V139 -22629.453616530704
L4_139 V4 V139 -1.5361820058536744e-12
C4_139 V4 V139 3.551053574217392e-19

R4_140 V4 V140 -35373.63513833331
L4_140 V4 V140 9.446063787885951e-13
C4_140 V4 V140 -7.004457458173851e-19

R4_141 V4 V141 14718.8886650583
L4_141 V4 V141 -9.030928277656028e-11
C4_141 V4 V141 -1.7953458552501448e-20

R4_142 V4 V142 14281.772815236007
L4_142 V4 V142 -7.0695124070806555e-12
C4_142 V4 V142 5.607259898327614e-20

R4_143 V4 V143 11293.261497666177
L4_143 V4 V143 1.7314723257799573e-10
C4_143 V4 V143 -6.496964959611202e-20

R4_144 V4 V144 -2786.948870166464
L4_144 V4 V144 -2.240274828725673e-11
C4_144 V4 V144 5.597346667331419e-20

R4_145 V4 V145 -5609.9542049269985
L4_145 V4 V145 4.100403040263072e-12
C4_145 V4 V145 -9.62069121238521e-20

R4_146 V4 V146 -9383.054868230185
L4_146 V4 V146 2.6001496801021904e-12
C4_146 V4 V146 -8.820944530283762e-20

R4_147 V4 V147 43054.86978840063
L4_147 V4 V147 6.550750041620619e-12
C4_147 V4 V147 -8.5948180011497e-20

R4_148 V4 V148 1437.027627498576
L4_148 V4 V148 -9.555580738867095e-13
C4_148 V4 V148 4.333377427924774e-19

R4_149 V4 V149 6503.603260243094
L4_149 V4 V149 -1.470090682516895e-11
C4_149 V4 V149 1.5504123145817213e-19

R4_150 V4 V150 10830.07591598154
L4_150 V4 V150 -6.394255621303757e-12
C4_150 V4 V150 4.806021343234097e-20

R4_151 V4 V151 -4122.74842680901
L4_151 V4 V151 6.1519129743908084e-12
C4_151 V4 V151 8.539568433457522e-20

R4_152 V4 V152 -6398.273648769772
L4_152 V4 V152 2.5653554016056788e-12
C4_152 V4 V152 -1.4396440039089164e-19

R4_153 V4 V153 -5839.4595225284265
L4_153 V4 V153 1.698042421156309e-11
C4_153 V4 V153 1.42315887272203e-21

R4_154 V4 V154 -9387.316012548108
L4_154 V4 V154 8.740821110415077e-12
C4_154 V4 V154 7.583000265624586e-20

R4_155 V4 V155 2651.334043698254
L4_155 V4 V155 -5.7757997824315275e-12
C4_155 V4 V155 8.75570457051205e-20

R4_156 V4 V156 11305.457969378323
L4_156 V4 V156 2.8391558825985448e-12
C4_156 V4 V156 -2.5338230061541035e-19

R4_157 V4 V157 8106.685382589347
L4_157 V4 V157 -3.6048388966761985e-12
C4_157 V4 V157 1.0201120462188881e-19

R4_158 V4 V158 5029.598435272095
L4_158 V4 V158 -7.092406356330426e-12
C4_158 V4 V158 -4.969224997487093e-21

R4_159 V4 V159 12318.127192706392
L4_159 V4 V159 9.052544467839435e-12
C4_159 V4 V159 -4.898090342209266e-20

R4_160 V4 V160 -2147.375453839565
L4_160 V4 V160 -3.953925339208264e-11
C4_160 V4 V160 1.575272004754911e-19

R4_161 V4 V161 -9016.721924336049
L4_161 V4 V161 2.5582796833585334e-12
C4_161 V4 V161 -1.248868116343172e-19

R4_162 V4 V162 -47229.76429258996
L4_162 V4 V162 5.809420367623205e-12
C4_162 V4 V162 3.035774413651764e-20

R4_163 V4 V163 24865.339015296682
L4_163 V4 V163 8.1392731331356e-12
C4_163 V4 V163 7.704493105913682e-20

R4_164 V4 V164 1389.7207434377126
L4_164 V4 V164 -2.7676192114934135e-12
C4_164 V4 V164 -8.726478298682935e-20

R4_165 V4 V165 12574.787282065767
L4_165 V4 V165 -4.670878144944852e-12
C4_165 V4 V165 1.2292871243252353e-19

R4_166 V4 V166 18316.112561340156
L4_166 V4 V166 -1.9557497424936572e-11
C4_166 V4 V166 9.565975231769887e-20

R4_167 V4 V167 10108.49719310173
L4_167 V4 V167 4.82100865636682e-11
C4_167 V4 V167 -3.3598542607536726e-20

R4_168 V4 V168 -2446.061024627677
L4_168 V4 V168 2.0017877099447486e-12
C4_168 V4 V168 -7.611932084307567e-20

R4_169 V4 V169 88443.91487183499
L4_169 V4 V169 -6.788743962360802e-12
C4_169 V4 V169 1.8405061358322565e-19

R4_170 V4 V170 178840.98593223045
L4_170 V4 V170 1.1441976043980351e-11
C4_170 V4 V170 9.709061133381462e-21

R4_171 V4 V171 -28175.275790157313
L4_171 V4 V171 8.453002792489225e-12
C4_171 V4 V171 5.2745913057396935e-20

R4_172 V4 V172 -4775.70704968532
L4_172 V4 V172 -2.6885553896950685e-12
C4_172 V4 V172 2.79443117629439e-20

R4_173 V4 V173 -8941.292024915436
L4_173 V4 V173 3.765420526634094e-12
C4_173 V4 V173 -1.1022389875391457e-19

R4_174 V4 V174 -48567.67610320253
L4_174 V4 V174 -7.9262165967924e-12
C4_174 V4 V174 2.1505640969323798e-20

R4_175 V4 V175 -47031.22652553266
L4_175 V4 V175 -3.813443406967756e-12
C4_175 V4 V175 8.081082031991334e-20

R4_176 V4 V176 2932.9453053832453
L4_176 V4 V176 2.876918018007594e-11
C4_176 V4 V176 -2.0369518006542045e-19

R4_177 V4 V177 8043.367959569785
L4_177 V4 V177 -8.000809450528863e-12
C4_177 V4 V177 3.8965966423983325e-20

R4_178 V4 V178 -117331.69687928855
L4_178 V4 V178 -2.6102589469531533e-11
C4_178 V4 V178 -4.9532669626598117e-20

R4_179 V4 V179 6829.2995701376585
L4_179 V4 V179 -2.939021865014184e-11
C4_179 V4 V179 -7.088594329177985e-20

R4_180 V4 V180 -8935.175511073103
L4_180 V4 V180 3.4175592877998014e-11
C4_180 V4 V180 1.4671353133397885e-19

R4_181 V4 V181 -107490.97956869549
L4_181 V4 V181 8.437500548058359e-11
C4_181 V4 V181 -3.3730291323559503e-20

R4_182 V4 V182 -8284.234118247137
L4_182 V4 V182 -1.975990231914534e-11
C4_182 V4 V182 5.478550231868964e-20

R4_183 V4 V183 -10183.860016070885
L4_183 V4 V183 -1.7485901380714816e-11
C4_183 V4 V183 4.540483983728885e-20

R4_184 V4 V184 24840.680729687138
L4_184 V4 V184 -5.29035539772933e-12
C4_184 V4 V184 -1.0289847332061786e-19

R4_185 V4 V185 -7280.389729885391
L4_185 V4 V185 6.571384178560795e-12
C4_185 V4 V185 5.108260860081832e-21

R4_186 V4 V186 7448.825158087586
L4_186 V4 V186 -5.403209330866092e-12
C4_186 V4 V186 -4.751484252669067e-20

R4_187 V4 V187 -32024.292081685864
L4_187 V4 V187 -6.032606903074988e-12
C4_187 V4 V187 -3.482872439118775e-20

R4_188 V4 V188 -4061.684667406049
L4_188 V4 V188 1.2709268631338689e-12
C4_188 V4 V188 -4.28151261072589e-20

R4_189 V4 V189 6473.65014278565
L4_189 V4 V189 -4.388990036759557e-12
C4_189 V4 V189 6.572611383226894e-20

R4_190 V4 V190 25453.906092246893
L4_190 V4 V190 1.1839322369457788e-11
C4_190 V4 V190 2.4899097753127894e-20

R4_191 V4 V191 -14279.547767935432
L4_191 V4 V191 2.2286712841712895e-12
C4_191 V4 V191 -2.6718449396659354e-20

R4_192 V4 V192 218873.9553314773
L4_192 V4 V192 -1.3576577665279005e-12
C4_192 V4 V192 2.553755377715929e-19

R4_193 V4 V193 -13488.759450198848
L4_193 V4 V193 -8.303908823017525e-11
C4_193 V4 V193 3.859907687054859e-21

R4_194 V4 V194 60527.47567538961
L4_194 V4 V194 -3.001162521414512e-12
C4_194 V4 V194 2.1220728792177096e-19

R4_195 V4 V195 7561.917684069331
L4_195 V4 V195 -1.7758449267693458e-12
C4_195 V4 V195 2.6175177666640077e-19

R4_196 V4 V196 9020.176771549974
L4_196 V4 V196 1.2864599009158815e-12
C4_196 V4 V196 -4.928148271068136e-19

R4_197 V4 V197 -7711.787691945903
L4_197 V4 V197 7.108246930581791e-12
C4_197 V4 V197 -1.2351439570460646e-19

R4_198 V4 V198 4974.022898921483
L4_198 V4 V198 -2.6304701234037867e-11
C4_198 V4 V198 1.0804728535445037e-19

R4_199 V4 V199 2087.474410058194
L4_199 V4 V199 1.5932712881480162e-11
C4_199 V4 V199 7.719852240588003e-20

R4_200 V4 V200 -3146.8057196197556
L4_200 V4 V200 1.9167502390538255e-11
C4_200 V4 V200 -6.623867618391642e-20

R5_5 V5 0 3216.9986563936914
L5_5 V5 0 1.5195466121928093e-13
C5_5 V5 0 1.0433353601265214e-18

R5_6 V5 V6 -8302.10410078876
L5_6 V5 V6 -8.25406796019906e-13
C5_6 V5 V6 -5.43129420747831e-19

R5_7 V5 V7 -10557.810498567263
L5_7 V5 V7 -9.42948372948979e-13
C5_7 V5 V7 -4.764202349189536e-19

R5_8 V5 V8 -13728.022139750617
L5_8 V5 V8 -8.671802933634776e-13
C5_8 V5 V8 -4.1495865895013974e-19

R5_9 V5 V9 12372.20367876603
L5_9 V5 V9 -1.7125706268223881e-12
C5_9 V5 V9 3.6825836392622074e-19

R5_10 V5 V10 18402.76230024495
L5_10 V5 V10 -1.9946958568344247e-12
C5_10 V5 V10 1.3870703233262682e-19

R5_11 V5 V11 17923.15414334357
L5_11 V5 V11 -2.6721679881913137e-12
C5_11 V5 V11 1.4938020875510162e-19

R5_12 V5 V12 17086.010280822615
L5_12 V5 V12 -2.1625938485468413e-12
C5_12 V5 V12 1.315280053094515e-19

R5_13 V5 V13 -4779.409239526077
L5_13 V5 V13 1.5938237328531193e-11
C5_13 V5 V13 -1.5908431936806933e-19

R5_14 V5 V14 -22923.581382696393
L5_14 V5 V14 2.6640400353522292e-12
C5_14 V5 V14 -4.802451899956043e-21

R5_15 V5 V15 -50405.003263582716
L5_15 V5 V15 2.014374881923399e-12
C5_15 V5 V15 7.399470132569645e-20

R5_16 V5 V16 -165635.76201955645
L5_16 V5 V16 1.3950319851933773e-12
C5_16 V5 V16 1.58650761346657e-19

R5_17 V5 V17 8030.749213215909
L5_17 V5 V17 1.018479194709751e-12
C5_17 V5 V17 1.3218868881102057e-19

R5_18 V5 V18 18878.902968490267
L5_18 V5 V18 2.5826916182670793e-12
C5_18 V5 V18 1.7997117646474665e-19

R5_19 V5 V19 83007.59328968804
L5_19 V5 V19 4.8735289555083645e-12
C5_19 V5 V19 3.54156912636525e-20

R5_20 V5 V20 79641.75049528664
L5_20 V5 V20 3.172403779555669e-12
C5_20 V5 V20 5.65116088045881e-20

R5_21 V5 V21 18143.320101297893
L5_21 V5 V21 6.283133894653123e-13
C5_21 V5 V21 1.2543985331186914e-19

R5_22 V5 V22 -25354.2503086276
L5_22 V5 V22 2.028766766322284e-12
C5_22 V5 V22 -1.190237606038037e-19

R5_23 V5 V23 -133281.87635743816
L5_23 V5 V23 1.8217936448429026e-12
C5_23 V5 V23 1.2952701615418227e-20

R5_24 V5 V24 -966266.8685370814
L5_24 V5 V24 1.391645326354847e-12
C5_24 V5 V24 4.9585845932787055e-20

R5_25 V5 V25 -8414.114927978635
L5_25 V5 V25 -6.521462581626008e-13
C5_25 V5 V25 -4.1402993240198187e-19

R5_26 V5 V26 65857.70840350748
L5_26 V5 V26 -1.7664819180419092e-12
C5_26 V5 V26 -1.3022972482700563e-20

R5_27 V5 V27 -34482.671999999395
L5_27 V5 V27 -1.225991384834244e-12
C5_27 V5 V27 -1.8977270997372784e-19

R5_28 V5 V28 -14748.258548962624
L5_28 V5 V28 -7.867382764124576e-13
C5_28 V5 V28 -3.5048931729683807e-19

R5_29 V5 V29 -35836.49842096409
L5_29 V5 V29 -9.135290358381286e-13
C5_29 V5 V29 -7.311973968773658e-20

R5_30 V5 V30 -391973.97280028847
L5_30 V5 V30 -2.3004175403234706e-12
C5_30 V5 V30 -4.655922398037961e-20

R5_31 V5 V31 81538.75421061584
L5_31 V5 V31 -3.0106334723214006e-12
C5_31 V5 V31 1.2144100246750791e-20

R5_32 V5 V32 251232.22796400404
L5_32 V5 V32 -2.254429345413972e-12
C5_32 V5 V32 -3.7559783741997424e-20

R5_33 V5 V33 -29727.43915666429
L5_33 V5 V33 2.3520455720729383e-12
C5_33 V5 V33 1.8181700966355557e-19

R5_34 V5 V34 46412.3950897997
L5_34 V5 V34 1.0350564133275899e-11
C5_34 V5 V34 1.221942003404425e-19

R5_35 V5 V35 38966.246910811926
L5_35 V5 V35 3.0101519544662486e-12
C5_35 V5 V35 1.552720134325055e-19

R5_36 V5 V36 124870.06701445024
L5_36 V5 V36 1.7008471824772506e-12
C5_36 V5 V36 1.6589075308982532e-19

R5_37 V5 V37 6059.356075343986
L5_37 V5 V37 8.066421923265687e-13
C5_37 V5 V37 4.0820522923226486e-19

R5_38 V5 V38 21995.53164397492
L5_38 V5 V38 1.450503876871588e-12
C5_38 V5 V38 2.3624489292151773e-19

R5_39 V5 V39 160500.1679364953
L5_39 V5 V39 2.7816924943787522e-12
C5_39 V5 V39 3.786678988182486e-20

R5_40 V5 V40 172267.65968549188
L5_40 V5 V40 1.8455834011290937e-12
C5_40 V5 V40 6.522059728637078e-20

R5_41 V5 V41 -17603.68228353306
L5_41 V5 V41 5.1497408887093445e-12
C5_41 V5 V41 -2.3029008363501695e-19

R5_42 V5 V42 -96696.55338766442
L5_42 V5 V42 -8.275145030852157e-12
C5_42 V5 V42 -9.046326514644345e-20

R5_43 V5 V43 -754690.0397096968
L5_43 V5 V43 8.04562601997402e-12
C5_43 V5 V43 -1.1382400637530699e-20

R5_44 V5 V44 -41646.52983997752
L5_44 V5 V44 1.8595909344922104e-11
C5_44 V5 V44 -9.52888765957016e-20

R5_45 V5 V45 -36730.369563874236
L5_45 V5 V45 -1.1661352524867232e-12
C5_45 V5 V45 -1.4848440909486077e-19

R5_46 V5 V46 -59038.78012876387
L5_46 V5 V46 -2.168546775605107e-12
C5_46 V5 V46 -1.8396519927182548e-19

R5_47 V5 V47 -59952.813514877394
L5_47 V5 V47 -2.4342343546962225e-12
C5_47 V5 V47 -1.2302302469913388e-19

R5_48 V5 V48 -31371.44918175364
L5_48 V5 V48 -1.2773944935182055e-12
C5_48 V5 V48 -2.3700423788496466e-19

R5_49 V5 V49 -26431.388120396572
L5_49 V5 V49 -7.445608248822446e-12
C5_49 V5 V49 -1.201277910757792e-19

R5_50 V5 V50 199610.2505127275
L5_50 V5 V50 1.3185276326569022e-11
C5_50 V5 V50 8.70167982980207e-20

R5_51 V5 V51 -62419.22350629028
L5_51 V5 V51 -4.036505973975228e-12
C5_51 V5 V51 -2.5499497806978963e-20

R5_52 V5 V52 -32055.943749273025
L5_52 V5 V52 -1.3836788399802236e-11
C5_52 V5 V52 -1.363588305078106e-20

R5_53 V5 V53 24462.05212239674
L5_53 V5 V53 -3.3038128959285337e-12
C5_53 V5 V53 1.4082301792345637e-19

R5_54 V5 V54 23100.951021933688
L5_54 V5 V54 4.776265305911684e-12
C5_54 V5 V54 1.8736285258713258e-19

R5_55 V5 V55 29054.441363252892
L5_55 V5 V55 2.6201106008702346e-11
C5_55 V5 V55 1.12207222305224e-19

R5_56 V5 V56 24460.568757700687
L5_56 V5 V56 2.5233192239170446e-12
C5_56 V5 V56 2.051672279571837e-19

R5_57 V5 V57 8866.64486158813
L5_57 V5 V57 6.768585953152905e-13
C5_57 V5 V57 4.595184639401364e-19

R5_58 V5 V58 525569.5344894503
L5_58 V5 V58 -7.454054678391476e-12
C5_58 V5 V58 -4.470031679876213e-20

R5_59 V5 V59 492472.752520131
L5_59 V5 V59 7.57101502680202e-12
C5_59 V5 V59 -3.0417373546139086e-20

R5_60 V5 V60 -225891.23695892558
L5_60 V5 V60 3.740806165692643e-12
C5_60 V5 V60 -5.705228970348944e-20

R5_61 V5 V61 -6932.871778198138
L5_61 V5 V61 -1.0772619391206919e-12
C5_61 V5 V61 -4.743329433443211e-19

R5_62 V5 V62 -379797.76634623273
L5_62 V5 V62 -2.6991721079183638e-11
C5_62 V5 V62 -5.333649469044164e-20

R5_63 V5 V63 32336.227533183093
L5_63 V5 V63 3.5492990082581064e-12
C5_63 V5 V63 9.592642755943176e-20

R5_64 V5 V64 141533.4069357807
L5_64 V5 V64 -5.1373986949449294e-11
C5_64 V5 V64 -1.26028501079264e-20

R5_65 V5 V65 -61843.332904770745
L5_65 V5 V65 3.539601254545557e-11
C5_65 V5 V65 -4.2357369963348246e-20

R5_66 V5 V66 55950.04005336857
L5_66 V5 V66 3.5773438151613457e-12
C5_66 V5 V66 1.394142107113474e-19

R5_67 V5 V67 327800.9825455072
L5_67 V5 V67 4.235156133480074e-12
C5_67 V5 V67 1.0472722713451592e-19

R5_68 V5 V68 -39591.21043263394
L5_68 V5 V68 -2.012833928815405e-11
C5_68 V5 V68 3.4834383319014974e-21

R5_69 V5 V69 -57941.83837710084
L5_69 V5 V69 -1.5023800627845428e-12
C5_69 V5 V69 -1.8199050817930713e-19

R5_70 V5 V70 -86938.47967157324
L5_70 V5 V70 -4.484200217400345e-12
C5_70 V5 V70 -8.361636505283057e-20

R5_71 V5 V71 -17711.01014816503
L5_71 V5 V71 -1.3802630264546308e-12
C5_71 V5 V71 -2.414725015482332e-19

R5_72 V5 V72 -27841.76622337468
L5_72 V5 V72 -1.5701191560954359e-12
C5_72 V5 V72 -1.6947554493562775e-19

R5_73 V5 V73 14908.936186452627
L5_73 V5 V73 -1.801901549493804e-11
C5_73 V5 V73 1.8278291486032837e-19

R5_74 V5 V74 91892.41896284964
L5_74 V5 V74 -3.3170302470597447e-12
C5_74 V5 V74 -7.724912732390395e-20

R5_75 V5 V75 43082.97551738537
L5_75 V5 V75 -7.666186017031571e-12
C5_75 V5 V75 -4.362566620308327e-20

R5_76 V5 V76 30112.627570437427
L5_76 V5 V76 3.1195120503898936e-12
C5_76 V5 V76 4.7287927306602593e-20

R5_77 V5 V77 14042.691934082739
L5_77 V5 V77 7.015633966657163e-13
C5_77 V5 V77 4.569636585628018e-19

R5_78 V5 V78 201531.67688010097
L5_78 V5 V78 3.846686648931325e-12
C5_78 V5 V78 1.3014100490307872e-19

R5_79 V5 V79 151278.97467006047
L5_79 V5 V79 2.248403957144625e-12
C5_79 V5 V79 1.5443617844457161e-19

R5_80 V5 V80 -70573.77672666812
L5_80 V5 V80 3.745229604103038e-12
C5_80 V5 V80 9.952048525748062e-20

R5_81 V5 V81 -9200.604878078166
L5_81 V5 V81 -1.0834902863531363e-12
C5_81 V5 V81 -4.6192703694413405e-19

R5_82 V5 V82 139799.55897706913
L5_82 V5 V82 7.446745117175598e-12
C5_82 V5 V82 6.954763903093158e-20

R5_83 V5 V83 27654.783327475412
L5_83 V5 V83 3.0312849230716025e-12
C5_83 V5 V83 1.6897335189890153e-19

R5_84 V5 V84 134873.64530774867
L5_84 V5 V84 5.030306021324081e-12
C5_84 V5 V84 5.548878145708987e-20

R5_85 V5 V85 -30141.631027311272
L5_85 V5 V85 -6.3129322210060795e-12
C5_85 V5 V85 -1.319685496431769e-19

R5_86 V5 V86 -55656.35601297887
L5_86 V5 V86 -2.207886896500973e-12
C5_86 V5 V86 -1.7456160371912801e-19

R5_87 V5 V87 -174427.6621345765
L5_87 V5 V87 -5.992173359058551e-12
C5_87 V5 V87 -1.0832182461973093e-19

R5_88 V5 V88 -106253.97841259904
L5_88 V5 V88 -3.721560508686854e-12
C5_88 V5 V88 -1.4127959260229289e-19

R5_89 V5 V89 -77879.35064599985
L5_89 V5 V89 -2.7641449019319086e-12
C5_89 V5 V89 -1.0361319203740019e-19

R5_90 V5 V90 19417.60400319063
L5_90 V5 V90 3.11952014954937e-12
C5_90 V5 V90 9.268896278552785e-20

R5_91 V5 V91 -18593.07437550412
L5_91 V5 V91 -1.1067728946755167e-12
C5_91 V5 V91 -3.2114420161622753e-19

R5_92 V5 V92 -27278.731039035134
L5_92 V5 V92 -1.5581615195151087e-12
C5_92 V5 V92 -1.9258800593094245e-19

R5_93 V5 V93 12479.017831299781
L5_93 V5 V93 1.9799822901396597e-12
C5_93 V5 V93 3.1827310841936154e-19

R5_94 V5 V94 -823953.8985930328
L5_94 V5 V94 6.080555392406897e-12
C5_94 V5 V94 1.1727902538724534e-19

R5_95 V5 V95 89184.28557264892
L5_95 V5 V95 2.204584177081752e-12
C5_95 V5 V95 1.9419240489081374e-19

R5_96 V5 V96 70616.51055404468
L5_96 V5 V96 1.4736694682839195e-12
C5_96 V5 V96 2.43098393373371e-19

R5_97 V5 V97 13568.743108581364
L5_97 V5 V97 1.124483967372757e-12
C5_97 V5 V97 3.8653471703336777e-19

R5_98 V5 V98 -59050.77934744165
L5_98 V5 V98 -2.1005651827185752e-12
C5_98 V5 V98 -1.0055800443119513e-19

R5_99 V5 V99 15481.649132516242
L5_99 V5 V99 1.7442810772861656e-12
C5_99 V5 V99 2.653864901250801e-19

R5_100 V5 V100 32377.83008690723
L5_100 V5 V100 3.5799524915538285e-12
C5_100 V5 V100 1.0019734134460579e-19

R5_101 V5 V101 -8323.9631798944
L5_101 V5 V101 -1.332466353827104e-12
C5_101 V5 V101 -4.9810312351368705e-19

R5_102 V5 V102 67130.90857773378
L5_102 V5 V102 7.044950979769652e-12
C5_102 V5 V102 3.402150558579681e-20

R5_103 V5 V103 -103533.87901457484
L5_103 V5 V103 -2.4997087979573948e-12
C5_103 V5 V103 -1.416041197327193e-19

R5_104 V5 V104 -44139.83219330009
L5_104 V5 V104 -2.342747352711525e-12
C5_104 V5 V104 -1.8391640301235328e-19

R5_105 V5 V105 -36786.16708549413
L5_105 V5 V105 -1.8655161844452823e-12
C5_105 V5 V105 -1.1103792924831318e-19

R5_106 V5 V106 27400.5670291134
L5_106 V5 V106 4.519779421579793e-12
C5_106 V5 V106 9.553477691241635e-20

R5_107 V5 V107 -35240.66847119225
L5_107 V5 V107 -4.8637248210603e-12
C5_107 V5 V107 -1.3456798800635865e-19

R5_108 V5 V108 -55094.225258172024
L5_108 V5 V108 -6.808145892442932e-12
C5_108 V5 V108 -7.510448870166022e-20

R5_109 V5 V109 14307.239340113621
L5_109 V5 V109 3.540133680437638e-12
C5_109 V5 V109 1.5681801570661889e-19

R5_110 V5 V110 -28926.940764753967
L5_110 V5 V110 -1.0983010579068477e-11
C5_110 V5 V110 -9.614333572206093e-20

R5_111 V5 V111 -1859905.044721373
L5_111 V5 V111 -4.383004884886514e-12
C5_111 V5 V111 -1.9419384568543043e-20

R5_112 V5 V112 34010.95224026063
L5_112 V5 V112 -1.3248497662083184e-11
C5_112 V5 V112 7.891754260090436e-20

R5_113 V5 V113 35295.072264634415
L5_113 V5 V113 1.7722528084297854e-12
C5_113 V5 V113 2.1422296820735714e-19

R5_114 V5 V114 -348190.5124284503
L5_114 V5 V114 1.316765679086984e-10
C5_114 V5 V114 2.031714496173521e-20

R5_115 V5 V115 23431.17558880391
L5_115 V5 V115 1.9268485630617303e-12
C5_115 V5 V115 2.250843616013164e-19

R5_116 V5 V116 35791.37164122621
L5_116 V5 V116 2.4588833458272604e-12
C5_116 V5 V116 1.8579177290663363e-19

R5_117 V5 V117 24907.57383810532
L5_117 V5 V117 1.6258477663946633e-12
C5_117 V5 V117 2.1875741562574926e-19

R5_118 V5 V118 45460.96814190774
L5_118 V5 V118 -6.846429704050068e-12
C5_118 V5 V118 1.0964479934964522e-20

R5_119 V5 V119 -51078.85670044473
L5_119 V5 V119 -8.962257264463922e-12
C5_119 V5 V119 -9.540342625784627e-20

R5_120 V5 V120 834314.600376898
L5_120 V5 V120 -3.0840362091563675e-11
C5_120 V5 V120 -7.16142376150806e-20

R5_121 V5 V121 -5858.230291940998
L5_121 V5 V121 -8.834754831569236e-13
C5_121 V5 V121 -6.149932777052607e-19

R5_122 V5 V122 -40365.40199833709
L5_122 V5 V122 -1.554295300539907e-11
C5_122 V5 V122 -4.104697323792599e-20

R5_123 V5 V123 -109226.42383390744
L5_123 V5 V123 -2.939559900427758e-12
C5_123 V5 V123 -3.4840158636161676e-20

R5_124 V5 V124 -22486.476175176605
L5_124 V5 V124 -2.0384338574919974e-12
C5_124 V5 V124 -1.4357839910667696e-19

R5_125 V5 V125 41553.647620532145
L5_125 V5 V125 -1.4333362908125553e-12
C5_125 V5 V125 -4.934795031122369e-20

R5_126 V5 V126 -23799.08502070251
L5_126 V5 V126 -6.39989203900429e-12
C5_126 V5 V126 -1.3780228859367728e-19

R5_127 V5 V127 -130981.90236352742
L5_127 V5 V127 4.953623898954552e-12
C5_127 V5 V127 -3.964230197082788e-21

R5_128 V5 V128 158686.9098300988
L5_128 V5 V128 6.458384861086151e-12
C5_128 V5 V128 2.4028511649848013e-20

R5_129 V5 V129 20224.210542279157
L5_129 V5 V129 1.124790573802453e-12
C5_129 V5 V129 3.269123581873825e-19

R5_130 V5 V130 20720.409578632494
L5_130 V5 V130 2.6937386777917417e-12
C5_130 V5 V130 1.6486420093541117e-19

R5_131 V5 V131 29573.22610860463
L5_131 V5 V131 -8.976875468841213e-12
C5_131 V5 V131 5.536352000579488e-20

R5_132 V5 V132 21556.382413318777
L5_132 V5 V132 1.4154905125808719e-11
C5_132 V5 V132 1.3988327090136216e-19

R5_133 V5 V133 20369.392789234098
L5_133 V5 V133 3.1119987258581475e-12
C5_133 V5 V133 -1.8083764526139826e-20

R5_134 V5 V134 -833140.6793356135
L5_134 V5 V134 1.558538863786034e-11
C5_134 V5 V134 -6.34863625475681e-20

R5_135 V5 V135 1180169.299643721
L5_135 V5 V135 1.774113905665461e-11
C5_135 V5 V135 -3.890312853922429e-20

R5_136 V5 V136 119336.41588029753
L5_136 V5 V136 -1.0981504626477736e-11
C5_136 V5 V136 -2.8935055960721116e-20

R5_137 V5 V137 15281.279063002474
L5_137 V5 V137 1.3896664250444697e-12
C5_137 V5 V137 3.091375174143537e-19

R5_138 V5 V138 -18883.408460598195
L5_138 V5 V138 -2.9001394055461037e-12
C5_138 V5 V138 -9.903927400823125e-20

R5_139 V5 V139 -24090.074799774073
L5_139 V5 V139 1.956639215650451e-11
C5_139 V5 V139 -1.2746858610989038e-20

R5_140 V5 V140 -38173.67864835858
L5_140 V5 V140 4.657239409181435e-12
C5_140 V5 V140 6.188070422343655e-20

R5_141 V5 V141 -6936.034312678704
L5_141 V5 V141 -7.694043715575938e-13
C5_141 V5 V141 -4.68215086062004e-19

R5_142 V5 V142 664039.1271121202
L5_142 V5 V142 1.908033471258191e-11
C5_142 V5 V142 4.014721843218819e-20

R5_143 V5 V143 26260.72719315522
L5_143 V5 V143 3.9378115653516927e-11
C5_143 V5 V143 7.68121810962916e-20

R5_144 V5 V144 -24116.9189531723
L5_144 V5 V144 -8.461024469556667e-12
C5_144 V5 V144 -1.4315727571074294e-19

R5_145 V5 V145 -10122.80489735046
L5_145 V5 V145 -8.484802344252122e-13
C5_145 V5 V145 -4.502238985915117e-19

R5_146 V5 V146 25616.75989971379
L5_146 V5 V146 4.4474841963153045e-11
C5_146 V5 V146 8.443521834281671e-20

R5_147 V5 V147 -11511.759455907948
L5_147 V5 V147 -1.9384613934168865e-12
C5_147 V5 V147 -3.156120116104057e-19

R5_148 V5 V148 36670.538279434055
L5_148 V5 V148 -1.5636154116839206e-12
C5_148 V5 V148 -1.1610132654004575e-19

R5_149 V5 V149 11147.745105297385
L5_149 V5 V149 6.694151679855344e-13
C5_149 V5 V149 5.449613874541102e-19

R5_150 V5 V150 53339.021848113705
L5_150 V5 V150 -1.8542201115860626e-12
C5_150 V5 V150 -1.4766205564607478e-19

R5_151 V5 V151 15494.926183128411
L5_151 V5 V151 -3.2534286152666132e-12
C5_151 V5 V151 8.269729447784726e-20

R5_152 V5 V152 321745.0871802677
L5_152 V5 V152 5.820333303450241e-12
C5_152 V5 V152 6.711101294120655e-20

R5_153 V5 V153 6133.98715101818
L5_153 V5 V153 8.975319170838375e-13
C5_153 V5 V153 5.553901676264132e-19

R5_154 V5 V154 85161.71937360619
L5_154 V5 V154 1.5482342342806968e-12
C5_154 V5 V154 1.6577832769045602e-19

R5_155 V5 V155 -11310.645028093617
L5_155 V5 V155 1.5086733992066662e-12
C5_155 V5 V155 -6.502083289248337e-20

R5_156 V5 V156 15064.76449234699
L5_156 V5 V156 2.83940232492247e-12
C5_156 V5 V156 2.159115359087451e-19

R5_157 V5 V157 18277.422591710685
L5_157 V5 V157 -3.8287452782891075e-12
C5_157 V5 V157 -1.2445501515961022e-19

R5_158 V5 V158 83729.88281230617
L5_158 V5 V158 1.7462596815676217e-11
C5_158 V5 V158 7.504382353171344e-20

R5_159 V5 V159 11300.605884790244
L5_159 V5 V159 3.050208061539073e-12
C5_159 V5 V159 2.781031911655e-19

R5_160 V5 V160 -20335.559533502346
L5_160 V5 V160 2.8964992460693028e-12
C5_160 V5 V160 -1.3706291083284245e-20

R5_161 V5 V161 -3927.3716915397686
L5_161 V5 V161 -8.997098790177625e-13
C5_161 V5 V161 -6.991349252955732e-19

R5_162 V5 V162 15493.723770909037
L5_162 V5 V162 6.586895554084585e-11
C5_162 V5 V162 1.9473081488418154e-19

R5_163 V5 V163 65123.496637350545
L5_163 V5 V163 -3.353866608321166e-11
C5_163 V5 V163 5.3380569080737033e-20

R5_164 V5 V164 29545.743802971243
L5_164 V5 V164 -2.1759536752971197e-12
C5_164 V5 V164 -1.4891505098772643e-20

R5_165 V5 V165 17368.28761542112
L5_165 V5 V165 -2.2971228754356445e-12
C5_165 V5 V165 1.352265960073235e-19

R5_166 V5 V166 -27649.31714527394
L5_166 V5 V166 -1.0631069710346522e-12
C5_166 V5 V166 -2.950912703666319e-19

R5_167 V5 V167 -43553.694362994
L5_167 V5 V167 -1.3820443376322214e-12
C5_167 V5 V167 -1.9301727702989674e-19

R5_168 V5 V168 -8308.540753051442
L5_168 V5 V168 -1.8252467192591067e-12
C5_168 V5 V168 -3.821825225874874e-19

R5_169 V5 V169 11688.46603374355
L5_169 V5 V169 1.2625576288917928e-12
C5_169 V5 V169 4.330444506282747e-19

R5_170 V5 V170 -58828.76681739193
L5_170 V5 V170 3.020407204375775e-12
C5_170 V5 V170 5.637867082671964e-20

R5_171 V5 V171 -22385.513125112084
L5_171 V5 V171 1.3079358635070185e-11
C5_171 V5 V171 -7.322609857142196e-20

R5_172 V5 V172 102271.49525064045
L5_172 V5 V172 4.002837352608887e-12
C5_172 V5 V172 1.1826208090691753e-19

R5_173 V5 V173 23180.18615679294
L5_173 V5 V173 2.7830793654833435e-12
C5_173 V5 V173 1.118117282726015e-19

R5_174 V5 V174 11673.654550954912
L5_174 V5 V174 6.158107145924305e-13
C5_174 V5 V174 4.610606557547809e-19

R5_175 V5 V175 8543.868113735358
L5_175 V5 V175 8.653430487714334e-13
C5_175 V5 V175 3.892677764496071e-19

R5_176 V5 V176 6793.584460521012
L5_176 V5 V176 7.198488730457402e-13
C5_176 V5 V176 4.556579377694262e-19

R5_177 V5 V177 -19129.806625908688
L5_177 V5 V177 -7.471593668954225e-12
C5_177 V5 V177 -2.747550441886196e-19

R5_178 V5 V178 171755.9539890119
L5_178 V5 V178 -1.2455816958565354e-12
C5_178 V5 V178 -1.6905613995831433e-19

R5_179 V5 V179 -20903.92903706137
L5_179 V5 V179 -1.6320310731858058e-12
C5_179 V5 V179 -1.7409927878680177e-19

R5_180 V5 V180 -16003.311393661941
L5_180 V5 V180 -9.662486487214468e-13
C5_180 V5 V180 -2.775817512179984e-19

R5_181 V5 V181 -6763.199047161738
L5_181 V5 V181 -4.643181295756802e-12
C5_181 V5 V181 -3.835843882011904e-19

R5_182 V5 V182 -100833.6232019743
L5_182 V5 V182 -4.573060331185495e-12
C5_182 V5 V182 -1.310542279421847e-20

R5_183 V5 V183 -75521.50546487761
L5_183 V5 V183 -8.106843619047574e-12
C5_183 V5 V183 9.177284407186976e-21

R5_184 V5 V184 -23503.333336681113
L5_184 V5 V184 -2.5761444817286136e-12
C5_184 V5 V184 -8.468596316143734e-20

R5_185 V5 V185 5527.906003869692
L5_185 V5 V185 -1.1306243477527043e-12
C5_185 V5 V185 4.302753537659758e-19

R5_186 V5 V186 -9480.855451891499
L5_186 V5 V186 -2.855386625134295e-12
C5_186 V5 V186 -2.4022780277388414e-19

R5_187 V5 V187 -48310.690645080314
L5_187 V5 V187 -6.264340111410075e-12
C5_187 V5 V187 -6.483039510869389e-20

R5_188 V5 V188 -25747.86765275675
L5_188 V5 V188 2.3500179400866497e-11
C5_188 V5 V188 -8.727968800115688e-20

R5_189 V5 V189 -32507.98956573852
L5_189 V5 V189 1.254745600648887e-12
C5_189 V5 V189 -1.260331209831625e-20

R5_190 V5 V190 18863.20419661502
L5_190 V5 V190 4.72646648289204e-12
C5_190 V5 V190 6.786825189119469e-20

R5_191 V5 V191 19159.671682644606
L5_191 V5 V191 -1.6899908620411874e-11
C5_191 V5 V191 5.6798983499696135e-21

R5_192 V5 V192 9976.325750284543
L5_192 V5 V192 3.0199947471959957e-12
C5_192 V5 V192 1.9460350416389635e-19

R5_193 V5 V193 -90645.32143822244
L5_193 V5 V193 1.460161395129552e-12
C5_193 V5 V193 1.430203867668206e-19

R5_194 V5 V194 9722.176440909412
L5_194 V5 V194 1.1422107666107456e-12
C5_194 V5 V194 4.0052403791799753e-19

R5_195 V5 V195 -103200.93068205199
L5_195 V5 V195 1.3541179194579867e-11
C5_195 V5 V195 3.599943948927101e-20

R5_196 V5 V196 23119.691056163767
L5_196 V5 V196 1.825975707546441e-12
C5_196 V5 V196 1.5709292949193743e-19

R5_197 V5 V197 -12162.149426945653
L5_197 V5 V197 -1.716453709329489e-12
C5_197 V5 V197 -3.3605727985453076e-19

R5_198 V5 V198 384564.8217410545
L5_198 V5 V198 -6.974314401156496e-12
C5_198 V5 V198 -2.232269695741676e-21

R5_199 V5 V199 20781.130223532688
L5_199 V5 V199 3.8476719278404334e-12
C5_199 V5 V199 2.2180254684910956e-19

R5_200 V5 V200 -6941.114387555944
L5_200 V5 V200 -2.2400881737195633e-12
C5_200 V5 V200 -2.8728639194378475e-19

R6_6 V6 0 658.0924929254437
L6_6 V6 0 1.7254751608244288e-13
C6_6 V6 0 3.821343131101104e-18

R6_7 V6 V7 -5806.5409138617415
L6_7 V6 V7 -5.905337497317518e-13
C6_7 V6 V7 -9.003270731086524e-19

R6_8 V6 V8 -9612.118691517579
L6_8 V6 V8 -6.138233153937757e-13
C6_8 V6 V8 -6.866046797316464e-19

R6_9 V6 V9 -8225.58486802893
L6_9 V6 V9 -2.2299083785555805e-12
C6_9 V6 V9 1.0230077087655195e-19

R6_10 V6 V10 -22599.212855421636
L6_10 V6 V10 1.3798790189370462e-12
C6_10 V6 V10 2.649113433200902e-19

R6_11 V6 V11 9428.370150892652
L6_11 V6 V11 3.1710020553590875e-11
C6_11 V6 V11 3.519134284280869e-19

R6_12 V6 V12 10643.370040646221
L6_12 V6 V12 -1.4590493516581122e-11
C6_12 V6 V12 2.7976352580496915e-19

R6_13 V6 V13 94988.3562163509
L6_13 V6 V13 8.054487986524847e-12
C6_13 V6 V13 9.638440146999206e-21

R6_14 V6 V14 9673.22853518177
L6_14 V6 V14 4.67983098791763e-13
C6_14 V6 V14 1.1633605606676552e-18

R6_15 V6 V15 47502.3778568536
L6_15 V6 V15 9.46202551912739e-13
C6_15 V6 V15 3.2850369466125865e-19

R6_16 V6 V16 13489.840506432081
L6_16 V6 V16 6.861089881196928e-13
C6_16 V6 V16 5.497158037463475e-19

R6_17 V6 V17 26239.926677160543
L6_17 V6 V17 5.5118153396142086e-12
C6_17 V6 V17 2.8507267718024793e-20

R6_18 V6 V18 12035.28800498913
L6_18 V6 V18 -4.95455208582332e-11
C6_18 V6 V18 -2.537705944122359e-19

R6_19 V6 V19 -32340.089001030898
L6_19 V6 V19 -6.2775138546525405e-12
C6_19 V6 V19 -1.2782813603049704e-19

R6_20 V6 V20 -22844.62156884328
L6_20 V6 V20 -7.172562403409768e-12
C6_20 V6 V20 -1.3017990543869679e-19

R6_21 V6 V21 5583.1869966742515
L6_21 V6 V21 1.1274663427348078e-12
C6_21 V6 V21 1.9949119592243114e-19

R6_22 V6 V22 8625.70716807077
L6_22 V6 V22 -2.0092142227201453e-12
C6_22 V6 V22 -1.8218610374208447e-19

R6_23 V6 V23 -564629.3533151416
L6_23 V6 V23 3.0512871838886603e-12
C6_23 V6 V23 -1.9344190103157313e-20

R6_24 V6 V24 59218.3710112509
L6_24 V6 V24 2.169719409874818e-12
C6_24 V6 V24 4.239052810312314e-20

R6_25 V6 V25 -7947.211228959236
L6_25 V6 V25 -2.4519732434786974e-12
C6_25 V6 V25 -1.529860715558964e-19

R6_26 V6 V26 -4239.065021554192
L6_26 V6 V26 -5.65731659712202e-12
C6_26 V6 V26 -1.4997907141612726e-19

R6_27 V6 V27 -34214.48799579537
L6_27 V6 V27 -1.9150525728403666e-12
C6_27 V6 V27 -8.283165115507649e-20

R6_28 V6 V28 -12451.269422564988
L6_28 V6 V28 -1.0542372493089588e-12
C6_28 V6 V28 -2.876660861050115e-19

R6_29 V6 V29 -6178.1560782642455
L6_29 V6 V29 -9.55484916831665e-13
C6_29 V6 V29 -3.6495536495852165e-19

R6_30 V6 V30 -32832.018044372184
L6_30 V6 V30 2.3911205019609475e-12
C6_30 V6 V30 1.5275835493779658e-19

R6_31 V6 V31 50980.89842422525
L6_31 V6 V31 -3.6273700724979125e-12
C6_31 V6 V31 -8.595295404912437e-21

R6_32 V6 V32 -592763.2248379855
L6_32 V6 V32 -2.479419360375045e-12
C6_32 V6 V32 -1.1197623606254292e-19

R6_33 V6 V33 57992.67122669
L6_33 V6 V33 9.536567370401794e-13
C6_33 V6 V33 4.506175274417337e-19

R6_34 V6 V34 25583.212418620908
L6_34 V6 V34 2.971339108148359e-12
C6_34 V6 V34 -9.612708048199498e-20

R6_35 V6 V35 10490.589294363283
L6_35 V6 V35 1.5760275223698586e-12
C6_35 V6 V35 3.3830384297436172e-19

R6_36 V6 V36 10654.481381308353
L6_36 V6 V36 1.1011136084142835e-12
C6_36 V6 V36 3.6590318474178145e-19

R6_37 V6 V37 7876.194547639044
L6_37 V6 V37 1.148138602258429e-12
C6_37 V6 V37 3.708289212109266e-19

R6_38 V6 V38 8685.79435614922
L6_38 V6 V38 2.5128210627035882e-12
C6_38 V6 V38 2.869911723791251e-19

R6_39 V6 V39 -46615.89612252752
L6_39 V6 V39 5.457395364275121e-12
C6_39 V6 V39 1.4500084880865445e-20

R6_40 V6 V40 -22628.498642317518
L6_40 V6 V40 5.256129213031679e-12
C6_40 V6 V40 -2.3114367113147753e-20

R6_41 V6 V41 -16773.346447839223
L6_41 V6 V41 -1.688867527279171e-12
C6_41 V6 V41 -3.927793172491628e-19

R6_42 V6 V42 18574.260416698882
L6_42 V6 V42 2.2032574955510355e-12
C6_42 V6 V42 1.4355010229464897e-19

R6_43 V6 V43 38734.540875620485
L6_43 V6 V43 -6.678960609761471e-11
C6_43 V6 V43 -1.8148604910144915e-20

R6_44 V6 V44 446186.5784398354
L6_44 V6 V44 -5.907021289882135e-12
C6_44 V6 V44 -1.3381459648268973e-19

R6_45 V6 V45 -8268.389073110482
L6_45 V6 V45 -1.203947952864315e-12
C6_45 V6 V45 -3.198790604391296e-19

R6_46 V6 V46 -4186.12485058194
L6_46 V6 V46 -6.283420366492775e-13
C6_46 V6 V46 -7.53453224491442e-19

R6_47 V6 V47 -18478.407168436694
L6_47 V6 V47 -1.2708291220519792e-12
C6_47 V6 V47 -3.12566988674302e-19

R6_48 V6 V48 -10982.508012016031
L6_48 V6 V48 -8.208402776102776e-13
C6_48 V6 V48 -4.837000605662495e-19

R6_49 V6 V49 -20216.24235136714
L6_49 V6 V49 3.041093372725297e-12
C6_49 V6 V49 1.2153478601341987e-19

R6_50 V6 V50 31118.12735172281
L6_50 V6 V50 1.4646110520419218e-12
C6_50 V6 V50 2.9313390828203676e-19

R6_51 V6 V51 15709.475867736084
L6_51 V6 V51 2.6530600820661286e-12
C6_51 V6 V51 3.6394086422317085e-19

R6_52 V6 V52 14181.29122680418
L6_52 V6 V52 1.5329399832909598e-12
C6_52 V6 V52 4.629181828369689e-19

R6_53 V6 V53 17422.485440877288
L6_53 V6 V53 1.766764100082951e-12
C6_53 V6 V53 2.964107777009364e-19

R6_54 V6 V54 4902.195729898361
L6_54 V6 V54 1.3122066758959992e-12
C6_54 V6 V54 4.499081018677978e-19

R6_55 V6 V55 12879.185827962712
L6_55 V6 V55 2.494956055925827e-12
C6_55 V6 V55 2.0318184734286732e-19

R6_56 V6 V56 8696.292890697729
L6_56 V6 V56 1.1357384124844397e-12
C6_56 V6 V56 3.581906367543058e-19

R6_57 V6 V57 494589.8623379971
L6_57 V6 V57 1.8760162352161455e-11
C6_57 V6 V57 -7.546679253075235e-23

R6_58 V6 V58 -43372.45510746148
L6_58 V6 V58 6.553401717057729e-12
C6_58 V6 V58 -1.290985819465217e-19

R6_59 V6 V59 -12351.515512723177
L6_59 V6 V59 -1.3538238711829573e-12
C6_59 V6 V59 -4.431068938096221e-19

R6_60 V6 V60 -8326.988232539177
L6_60 V6 V60 -1.0457024245784871e-12
C6_60 V6 V60 -6.349887490184254e-19

R6_61 V6 V61 -14569.539147522008
L6_61 V6 V61 -1.8031786140737665e-12
C6_61 V6 V61 -2.740141079908612e-19

R6_62 V6 V62 -8311.900616889841
L6_62 V6 V62 -3.1733592138442756e-12
C6_62 V6 V62 -1.4313999847919746e-19

R6_63 V6 V63 43020.6346672737
L6_63 V6 V63 2.9821211685066194e-12
C6_63 V6 V63 2.163101046688611e-19

R6_64 V6 V64 -46494.20174168241
L6_64 V6 V64 2.4745513153008066e-11
C6_64 V6 V64 1.1597032995854235e-19

R6_65 V6 V65 -11019.927568142766
L6_65 V6 V65 -4.843750435428755e-12
C6_65 V6 V65 -1.5724250967361172e-19

R6_66 V6 V66 -27250.31075979363
L6_66 V6 V66 -2.3406078792326845e-12
C6_66 V6 V66 -2.9814792087458807e-19

R6_67 V6 V67 11071.881861559488
L6_67 V6 V67 2.0613663478577565e-12
C6_67 V6 V67 3.0727149868789565e-19

R6_68 V6 V68 15926.247996705186
L6_68 V6 V68 5.11733665094811e-12
C6_68 V6 V68 1.9926743457603995e-19

R6_69 V6 V69 11392.75365802692
L6_69 V6 V69 1.6218009867898971e-12
C6_69 V6 V69 3.0090574907007225e-19

R6_70 V6 V70 38785.84664365685
L6_70 V6 V70 2.7138462359367874e-12
C6_70 V6 V70 1.436300279358152e-19

R6_71 V6 V71 -16176.488339246465
L6_71 V6 V71 -1.2866470663421929e-12
C6_71 V6 V71 -3.792369422243191e-19

R6_72 V6 V72 821715.7007301069
L6_72 V6 V72 -1.9772862357871555e-12
C6_72 V6 V72 -2.5183740828389027e-19

R6_73 V6 V73 -178692.6453286907
L6_73 V6 V73 -2.114442697726978e-11
C6_73 V6 V73 5.478679530890399e-21

R6_74 V6 V74 6558.213032527324
L6_74 V6 V74 7.254355699714243e-13
C6_74 V6 V74 6.2982272219001185e-19

R6_75 V6 V75 -22940.1464963682
L6_75 V6 V75 -2.9201871665075754e-11
C6_75 V6 V75 -8.876186145651888e-20

R6_76 V6 V76 -301103.54984459386
L6_76 V6 V76 1.4848896542365492e-12
C6_76 V6 V76 1.4871306216689829e-19

R6_77 V6 V77 -16734.107495420893
L6_77 V6 V77 -6.313837840047641e-12
C6_77 V6 V77 -1.3921052709320898e-19

R6_78 V6 V78 -8591.208361200654
L6_78 V6 V78 -1.0106701706360052e-12
C6_78 V6 V78 -6.098703549447895e-19

R6_79 V6 V79 1346022.0765987947
L6_79 V6 V79 5.178662685759217e-12
C6_79 V6 V79 1.0002988523380039e-19

R6_80 V6 V80 -14218.580890309044
L6_80 V6 V80 -2.4807707252820223e-12
C6_80 V6 V80 -1.3131620471881041e-19

R6_81 V6 V81 -6973.898598767576
L6_81 V6 V81 -2.9597211705519495e-12
C6_81 V6 V81 -2.567052580142121e-19

R6_82 V6 V82 -5919.072381053761
L6_82 V6 V82 -1.1462774873389197e-12
C6_82 V6 V82 -5.025823433960745e-19

R6_83 V6 V83 11640.820843209907
L6_83 V6 V83 8.5552590539405e-12
C6_83 V6 V83 1.5838434997658917e-19

R6_84 V6 V84 -101560.0552974327
L6_84 V6 V84 -1.6925117511583354e-12
C6_84 V6 V84 -2.208006681726326e-19

R6_85 V6 V85 763089.4355347669
L6_85 V6 V85 -4.006165836768972e-12
C6_85 V6 V85 -1.9905355212033832e-20

R6_86 V6 V86 6276.345671289232
L6_86 V6 V86 1.2521840002915346e-12
C6_86 V6 V86 5.5920239168234805e-19

R6_87 V6 V87 37279.10131065739
L6_87 V6 V87 1.0557809574466596e-11
C6_87 V6 V87 3.629252453754784e-20

R6_88 V6 V88 11594.797194028593
L6_88 V6 V88 1.9909844622283606e-12
C6_88 V6 V88 2.3218988981971405e-19

R6_89 V6 V89 9068.720065042991
L6_89 V6 V89 1.3257904959965012e-12
C6_89 V6 V89 3.3011698648463443e-19

R6_90 V6 V90 5608.129155082897
L6_90 V6 V90 8.423309335854375e-13
C6_90 V6 V90 5.025324452238225e-19

R6_91 V6 V91 -18398.71566904576
L6_91 V6 V91 -1.0791038285967278e-12
C6_91 V6 V91 -3.126107176113671e-19

R6_92 V6 V92 95239.99434531396
L6_92 V6 V92 -2.5550786868071814e-12
C6_92 V6 V92 -4.324751166861492e-20

R6_93 V6 V93 -13089.861948142463
L6_93 V6 V93 -6.816317360719762e-11
C6_93 V6 V93 -5.579840859330304e-20

R6_94 V6 V94 -6023.150306315641
L6_94 V6 V94 -8.945132452609939e-13
C6_94 V6 V94 -5.221451862939066e-19

R6_95 V6 V95 -12639.712506669375
L6_95 V6 V95 -1.6524375420625494e-11
C6_95 V6 V95 -1.1184960009520333e-19

R6_96 V6 V96 -7951.98246362232
L6_96 V6 V96 -6.371602134783398e-12
C6_96 V6 V96 -2.2352622906722e-19

R6_97 V6 V97 -6508.704973474478
L6_97 V6 V97 -1.1955211684571027e-12
C6_97 V6 V97 -3.642352050834592e-19

R6_98 V6 V98 -14419.928909386032
L6_98 V6 V98 -7.809846438880977e-12
C6_98 V6 V98 -1.98396538074556e-19

R6_99 V6 V99 4657.634812187308
L6_99 V6 V99 9.738513619570988e-13
C6_99 V6 V99 5.886635841645787e-19

R6_100 V6 V100 11419.802029352806
L6_100 V6 V100 7.492263156359363e-11
C6_100 V6 V100 8.292264858571185e-20

R6_101 V6 V101 12875.714517142822
L6_101 V6 V101 1.9358725297660008e-12
C6_101 V6 V101 1.7577571356065752e-19

R6_102 V6 V102 4461.257557143646
L6_102 V6 V102 9.774495710053934e-13
C6_102 V6 V102 4.729082885181125e-19

R6_103 V6 V103 14483.437007762437
L6_103 V6 V103 5.221719491434046e-12
C6_103 V6 V103 2.2839562716626847e-19

R6_104 V6 V104 15020.064227463874
L6_104 V6 V104 6.099446468712167e-12
C6_104 V6 V104 2.2761192932419222e-19

R6_105 V6 V105 132557.69538365194
L6_105 V6 V105 1.5311327566077489e-12
C6_105 V6 V105 3.606997044337896e-19

R6_106 V6 V106 -11483.3346971978
L6_106 V6 V106 -3.2093132459233773e-12
C6_106 V6 V106 -6.803247112023015e-20

R6_107 V6 V107 -5691.774772035366
L6_107 V6 V107 -8.400837548671893e-13
C6_107 V6 V107 -6.543468857151894e-19

R6_108 V6 V108 -48243.31697290916
L6_108 V6 V108 2.5221349195077017e-11
C6_108 V6 V108 -7.418237579561941e-20

R6_109 V6 V109 -16470.25350758632
L6_109 V6 V109 -1.437747576279975e-12
C6_109 V6 V109 -3.8121411363723527e-19

R6_110 V6 V110 -8465.959827256223
L6_110 V6 V110 -1.5385919890132435e-11
C6_110 V6 V110 -2.635124340749459e-19

R6_111 V6 V111 76586.20828373992
L6_111 V6 V111 -2.7924433380633004e-12
C6_111 V6 V111 -9.152643932608395e-20

R6_112 V6 V112 39417.97140505666
L6_112 V6 V112 -2.169803626920105e-12
C6_112 V6 V112 -8.021882480838603e-20

R6_113 V6 V113 -6933.974307028424
L6_113 V6 V113 -1.4922053990493093e-12
C6_113 V6 V113 -4.022204782163409e-19

R6_114 V6 V114 14455.043346726648
L6_114 V6 V114 7.279578746722131e-12
C6_114 V6 V114 -1.6525611125782852e-20

R6_115 V6 V115 7226.125552541783
L6_115 V6 V115 6.46665339076236e-13
C6_115 V6 V115 6.254900887524094e-19

R6_116 V6 V116 -148162.08298465962
L6_116 V6 V116 1.8726195905208284e-12
C6_116 V6 V116 1.336201045129757e-19

R6_117 V6 V117 16145.488735679633
L6_117 V6 V117 9.419198188469003e-13
C6_117 V6 V117 5.078075315126555e-19

R6_118 V6 V118 9692.466963713203
L6_118 V6 V118 7.316720872882964e-12
C6_118 V6 V118 3.0411895773422207e-19

R6_119 V6 V119 -70642.6912509051
L6_119 V6 V119 -3.23724755926348e-12
C6_119 V6 V119 -1.1065029687419572e-19

R6_120 V6 V120 14576.4718489529
L6_120 V6 V120 6.224841178046529e-12
C6_120 V6 V120 1.020579781423141e-19

R6_121 V6 V121 21016.646417083084
L6_121 V6 V121 2.479172554565206e-12
C6_121 V6 V121 1.3814332430162743e-19

R6_122 V6 V122 -6352.921185808485
L6_122 V6 V122 -1.9624570241595098e-12
C6_122 V6 V122 -4.71502340985836e-19

R6_123 V6 V123 -30029.304100328147
L6_123 V6 V123 -1.4596269162809036e-12
C6_123 V6 V123 -1.5511250969165618e-19

R6_124 V6 V124 -26099.620115803136
L6_124 V6 V124 -1.5031546766100432e-12
C6_124 V6 V124 -1.2475223708791686e-19

R6_125 V6 V125 -11657.642709685879
L6_125 V6 V125 -1.0268538177926552e-12
C6_125 V6 V125 -3.0115857573535775e-19

R6_126 V6 V126 -16080.597500557422
L6_126 V6 V126 -7.65987717489101e-12
C6_126 V6 V126 -2.6641003233787773e-20

R6_127 V6 V127 -13960.76027935066
L6_127 V6 V127 5.3222355665446264e-12
C6_127 V6 V127 -1.87725881176394e-19

R6_128 V6 V128 -12814.03636494173
L6_128 V6 V128 6.282463883996675e-12
C6_128 V6 V128 -1.961001787304375e-19

R6_129 V6 V129 -4384.56262962717
L6_129 V6 V129 -1.054039130072152e-12
C6_129 V6 V129 -6.719980565441871e-19

R6_130 V6 V130 5592.03328261729
L6_130 V6 V130 7.563069712571659e-13
C6_130 V6 V130 5.135381421668662e-19

R6_131 V6 V131 14484.389770815
L6_131 V6 V131 -4.3666848756199717e-10
C6_131 V6 V131 1.894400744894496e-19

R6_132 V6 V132 7368.888505265269
L6_132 V6 V132 2.615626943303978e-12
C6_132 V6 V132 4.005846917785217e-19

R6_133 V6 V133 3757.8976508960072
L6_133 V6 V133 4.999849734121629e-13
C6_133 V6 V133 8.652753065193011e-19

R6_134 V6 V134 -3891.849877555483
L6_134 V6 V134 -5.34577343433922e-13
C6_134 V6 V134 -1.0746169863140264e-18

R6_135 V6 V135 13218.911476470701
L6_135 V6 V135 2.7045667999400127e-12
C6_135 V6 V135 2.216727239348508e-19

R6_136 V6 V136 37192.00718827516
L6_136 V6 V136 -6.673420909518052e-12
C6_136 V6 V136 4.6599804429422444e-20

R6_137 V6 V137 6498.678245913999
L6_137 V6 V137 1.1878725620646343e-12
C6_137 V6 V137 6.572486650737006e-19

R6_138 V6 V138 14341.586193475998
L6_138 V6 V138 1.2999887676026638e-12
C6_138 V6 V138 5.843071127618717e-19

R6_139 V6 V139 -17284.0558844002
L6_139 V6 V139 2.7282716339743775e-12
C6_139 V6 V139 -9.481446179851474e-20

R6_140 V6 V140 -11810.386283292344
L6_140 V6 V140 3.8259113583487135e-12
C6_140 V6 V140 -1.6700510022657459e-19

R6_141 V6 V141 -2739.390394366619
L6_141 V6 V141 -3.543753280214166e-13
C6_141 V6 V141 -1.5248738753242915e-18

R6_142 V6 V142 7171.221915658679
L6_142 V6 V142 4.77772850020003e-13
C6_142 V6 V142 3.1619492251209864e-19

R6_143 V6 V143 -13406.508151565871
L6_143 V6 V143 -1.0318405765276468e-12
C6_143 V6 V143 -3.63353771703016e-19

R6_144 V6 V144 -19591.292277490014
L6_144 V6 V144 -4.709321765312226e-12
C6_144 V6 V144 -2.1231175467645054e-19

R6_145 V6 V145 -3478.183097592063
L6_145 V6 V145 -1.5877465507921424e-12
C6_145 V6 V145 -6.041776084120658e-19

R6_146 V6 V146 -8487.809014287934
L6_146 V6 V146 -4.394372658559318e-13
C6_146 V6 V146 -1.9697538927235957e-19

R6_147 V6 V147 -13494.834417313165
L6_147 V6 V147 -4.882282168038948e-12
C6_147 V6 V147 -9.342051513519359e-20

R6_148 V6 V148 346029.69066194067
L6_148 V6 V148 -1.3571389098961275e-12
C6_148 V6 V148 2.4651683494716217e-20

R6_149 V6 V149 1400.0737505809625
L6_149 V6 V149 2.3308309212260734e-13
C6_149 V6 V149 2.2117001519134894e-18

R6_150 V6 V150 -5092.378440767197
L6_150 V6 V150 -1.1145388993045703e-12
C6_150 V6 V150 -1.1919777014471936e-18

R6_151 V6 V151 5476.2294418916335
L6_151 V6 V151 1.873243790334267e-12
C6_151 V6 V151 4.386806239789977e-19

R6_152 V6 V152 15834.63667445675
L6_152 V6 V152 2.2715341621347405e-12
C6_152 V6 V152 -2.3046617098393586e-21

R6_153 V6 V153 18651.006601826815
L6_153 V6 V153 3.4130291839679654e-12
C6_153 V6 V153 3.9523178107703865e-19

R6_154 V6 V154 3674.9606994876704
L6_154 V6 V154 8.483470984785861e-13
C6_154 V6 V154 1.1080772348137508e-18

R6_155 V6 V155 -13184.8920179701
L6_155 V6 V155 9.89582143306949e-13
C6_155 V6 V155 6.22837426032455e-20

R6_156 V6 V156 37207.302073837214
L6_156 V6 V156 4.407721669934517e-12
C6_156 V6 V156 2.557500125923719e-19

R6_157 V6 V157 -1868.9075021905953
L6_157 V6 V157 -2.9343656771641783e-13
C6_157 V6 V157 -1.8541486899782798e-18

R6_158 V6 V158 -15997.896980195443
L6_158 V6 V158 9.075545411351786e-13
C6_158 V6 V158 -7.856259065711507e-20

R6_159 V6 V159 9409.051378398322
L6_159 V6 V159 -2.3966713357918285e-12
C6_159 V6 V159 3.0810004649070906e-19

R6_160 V6 V160 413373.10404638335
L6_160 V6 V160 8.27648448058899e-12
C6_160 V6 V160 1.7299524280821096e-19

R6_161 V6 V161 -5732.835258998126
L6_161 V6 V161 -2.9695228048214097e-12
C6_161 V6 V161 -4.551546315804203e-19

R6_162 V6 V162 16661.950426857773
L6_162 V6 V162 3.932857044089707e-12
C6_162 V6 V162 2.281975276762405e-19

R6_163 V6 V163 -14881.140387517276
L6_163 V6 V163 -1.4033178606471505e-12
C6_163 V6 V163 -4.452444768129374e-19

R6_164 V6 V164 17559.948052741714
L6_164 V6 V164 -2.652811218460095e-12
C6_164 V6 V164 -8.571525736365077e-20

R6_165 V6 V165 3760.2565220895954
L6_165 V6 V165 5.657270080500937e-13
C6_165 V6 V165 1.1531841054813778e-18

R6_166 V6 V166 13408.14809436749
L6_166 V6 V166 -1.0495109005593332e-12
C6_166 V6 V166 -2.1665328342361427e-19

R6_167 V6 V167 -55247.123658170596
L6_167 V6 V167 -4.577576639715394e-12
C6_167 V6 V167 -1.1508583161929155e-19

R6_168 V6 V168 -5671.428221069601
L6_168 V6 V168 -2.702981177166908e-12
C6_168 V6 V168 -5.734031601916025e-19

R6_169 V6 V169 17814.817485751017
L6_169 V6 V169 6.073946877353044e-12
C6_169 V6 V169 1.9418903711899784e-19

R6_170 V6 V170 143933.25755174167
L6_170 V6 V170 1.5720607756462636e-12
C6_170 V6 V170 4.820128529177354e-19

R6_171 V6 V171 8795.716466207314
L6_171 V6 V171 5.977112148094477e-13
C6_171 V6 V171 7.686598419981854e-19

R6_172 V6 V172 11135.979566036682
L6_172 V6 V172 1.0367179839611789e-12
C6_172 V6 V172 5.651244911066537e-19

R6_173 V6 V173 -5899.041160534781
L6_173 V6 V173 -1.3975558398512265e-12
C6_173 V6 V173 -3.639713368771804e-19

R6_174 V6 V174 -13977.456914018398
L6_174 V6 V174 9.211528993526335e-13
C6_174 V6 V174 -2.636283207160801e-19

R6_175 V6 V175 6025.251799772689
L6_175 V6 V175 1.5823755975363733e-12
C6_175 V6 V175 2.8743679982950935e-19

R6_176 V6 V176 6003.466444986912
L6_176 V6 V176 1.476558302407599e-12
C6_176 V6 V176 3.210006854435664e-19

R6_177 V6 V177 30664.590439281812
L6_177 V6 V177 -1.4350434578448846e-11
C6_177 V6 V177 8.737664014858584e-20

R6_178 V6 V178 -13532.935040584272
L6_178 V6 V178 -6.411760732198192e-13
C6_178 V6 V178 -4.458559324454892e-19

R6_179 V6 V179 -3222.0263174005513
L6_179 V6 V179 -5.218216022508167e-13
C6_179 V6 V179 -1.0113874206324694e-18

R6_180 V6 V180 -3925.0705869738563
L6_180 V6 V180 -4.972955019099717e-13
C6_180 V6 V180 -7.771562459774493e-19

R6_181 V6 V181 -20884.26054563029
L6_181 V6 V181 6.716976934862671e-11
C6_181 V6 V181 -3.7142993770826913e-19

R6_182 V6 V182 6115.220215035643
L6_182 V6 V182 5.113016225469635e-13
C6_182 V6 V182 6.252554335943365e-19

R6_183 V6 V183 -17232.985119986417
L6_183 V6 V183 -1.275880955540285e-12
C6_183 V6 V183 -1.1775939580084127e-19

R6_184 V6 V184 -20806.252472568645
L6_184 V6 V184 -2.3782701121437144e-12
C6_184 V6 V184 -6.625672656742542e-20

R6_185 V6 V185 -29407.454612075006
L6_185 V6 V185 -3.652955310652904e-12
C6_185 V6 V185 1.8576362354897048e-19

R6_186 V6 V186 59897.5533997379
L6_186 V6 V186 2.0714831596673295e-12
C6_186 V6 V186 -1.535215513887876e-19

R6_187 V6 V187 6059.044636550132
L6_187 V6 V187 6.520392908356081e-13
C6_187 V6 V187 5.487769053187759e-19

R6_188 V6 V188 8186.255090050204
L6_188 V6 V188 5.34508074061877e-13
C6_188 V6 V188 4.588179328643695e-19

R6_189 V6 V189 3998.555811085553
L6_189 V6 V189 1.2396910173004291e-12
C6_189 V6 V189 6.0691416240476895e-19

R6_190 V6 V190 -5622.976721183336
L6_190 V6 V190 -1.0125363540558323e-12
C6_190 V6 V190 -5.920481633639166e-19

R6_191 V6 V191 6150.553446692721
L6_191 V6 V191 7.925647145358101e-13
C6_191 V6 V191 6.148228426394841e-19

R6_192 V6 V192 6606.843177543655
L6_192 V6 V192 1.7722886966144814e-12
C6_192 V6 V192 5.557999091249504e-19

R6_193 V6 V193 -11820.761596871882
L6_193 V6 V193 -3.411289803912075e-12
C6_193 V6 V193 -2.8323687466200875e-19

R6_194 V6 V194 21530.037662198338
L6_194 V6 V194 1.3528041456632946e-12
C6_194 V6 V194 2.648566513369243e-19

R6_195 V6 V195 -3582.110473062673
L6_195 V6 V195 -4.534003198482422e-13
C6_195 V6 V195 -1.0153991526229047e-18

R6_196 V6 V196 -4670.485944678833
L6_196 V6 V196 -4.600907832117153e-13
C6_196 V6 V196 -9.019003480241308e-19

R6_197 V6 V197 -4091.5106945113666
L6_197 V6 V197 -8.527873228150833e-13
C6_197 V6 V197 -6.471434101243214e-19

R6_198 V6 V198 8896.148148297061
L6_198 V6 V198 2.5374289982683433e-12
C6_198 V6 V198 1.3532863886469678e-19

R6_199 V6 V199 -32081.012715512392
L6_199 V6 V199 -1.3382422205980853e-12
C6_199 V6 V199 -3.1411185371905113e-19

R6_200 V6 V200 -6539.380115168305
L6_200 V6 V200 -2.8103587378231415e-12
C6_200 V6 V200 -3.8675652190346754e-19

R7_7 V7 0 1140.156737724878
L7_7 V7 0 1.84916994512883e-13
C7_7 V7 0 2.150891669657797e-18

R7_8 V7 V8 -13101.120491031055
L7_8 V7 V8 -5.777367915520196e-13
C7_8 V7 V8 -6.436534870731887e-19

R7_9 V7 V9 -11404.396971993068
L7_9 V7 V9 -2.5262954550997042e-12
C7_9 V7 V9 1.0029573052074868e-19

R7_10 V7 V10 -27562.47687290382
L7_10 V7 V10 -1.4166931805108757e-11
C7_10 V7 V10 5.3967753876118456e-20

R7_11 V7 V11 -11373.244389594769
L7_11 V7 V11 6.403845845372621e-12
C7_11 V7 V11 4.2155957639924077e-19

R7_12 V7 V12 7253.455320569823
L7_12 V7 V12 4.4610051976654306e-11
C7_12 V7 V12 3.9797069158501054e-19

R7_13 V7 V13 58843.54272343212
L7_13 V7 V13 4.783522815178204e-12
C7_13 V7 V13 7.786165900468317e-20

R7_14 V7 V14 11502.513366033218
L7_14 V7 V14 1.318672856185901e-12
C7_14 V7 V14 5.284917522746298e-19

R7_15 V7 V15 11570.29332019593
L7_15 V7 V15 4.657153534056056e-13
C7_15 V7 V15 1.0551879311933172e-18

R7_16 V7 V16 22620.74546388226
L7_16 V7 V16 6.930227124059137e-13
C7_16 V7 V16 5.357343931282609e-19

R7_17 V7 V17 77624.01947000221
L7_17 V7 V17 8.768698766871484e-12
C7_17 V7 V17 -2.0912330959859403e-20

R7_18 V7 V18 85986.14898039092
L7_18 V7 V18 4.767726907323084e-12
C7_18 V7 V18 -1.6492289859426125e-21

R7_19 V7 V19 29707.013808245087
L7_19 V7 V19 -3.2739264542801818e-12
C7_19 V7 V19 -6.566278702359141e-19

R7_20 V7 V20 -15315.37990632638
L7_20 V7 V20 -7.0943929940997556e-12
C7_20 V7 V20 -2.3000065992785977e-19

R7_21 V7 V21 7293.007148836987
L7_21 V7 V21 1.2836329250773803e-12
C7_21 V7 V21 1.9051276174114061e-19

R7_22 V7 V22 22968.025644834375
L7_22 V7 V22 -7.8103366947414e-12
C7_22 V7 V22 -1.3899518498251673e-19

R7_23 V7 V23 4776.288681694748
L7_23 V7 V23 2.7227581474547367e-12
C7_23 V7 V23 2.5887552112989135e-19

R7_24 V7 V24 175505.26746926375
L7_24 V7 V24 2.198412385373277e-12
C7_24 V7 V24 5.0303064161804524e-20

R7_25 V7 V25 -10642.334510854726
L7_25 V7 V25 -2.3648387356421026e-12
C7_25 V7 V25 -1.3229947791139275e-19

R7_26 V7 V26 -14840.6398478463
L7_26 V7 V26 2.2065309652414718e-11
C7_26 V7 V26 7.26605952012688e-22

R7_27 V7 V27 -3557.1677518644688
L7_27 V7 V27 -1.2270053157394244e-12
C7_27 V7 V27 -4.726638058998035e-19

R7_28 V7 V28 -14911.11410945236
L7_28 V7 V28 -1.0940924591210022e-12
C7_28 V7 V28 -2.5135619554152917e-19

R7_29 V7 V29 -8199.0924028959
L7_29 V7 V29 -1.1258197429560995e-12
C7_29 V7 V29 -3.4686399648457023e-19

R7_30 V7 V30 -21982.732014327285
L7_30 V7 V30 -3.870907051891681e-12
C7_30 V7 V30 -1.0592563523964886e-19

R7_31 V7 V31 -30655.49195597883
L7_31 V7 V31 -1.0518004175396582e-11
C7_31 V7 V31 3.6007274123790885e-19

R7_32 V7 V32 42565.836529248794
L7_32 V7 V32 -2.4624897860547085e-12
C7_32 V7 V32 -8.18406031502938e-20

R7_33 V7 V33 52497.861835756645
L7_33 V7 V33 1.1626861888647947e-12
C7_33 V7 V33 4.0742087390570323e-19

R7_34 V7 V34 33134.79147151996
L7_34 V7 V34 2.2213708905097944e-12
C7_34 V7 V34 4.1174793215225223e-20

R7_35 V7 V35 8661.591151103448
L7_35 V7 V35 1.5501942663779801e-12
C7_35 V7 V35 2.7169884115235e-19

R7_36 V7 V36 13566.018096144531
L7_36 V7 V36 1.1293108876075142e-12
C7_36 V7 V36 3.7897917021680273e-19

R7_37 V7 V37 11209.33021716349
L7_37 V7 V37 1.4601991529952974e-12
C7_37 V7 V37 2.973430041345188e-19

R7_38 V7 V38 14526.041518558719
L7_38 V7 V38 1.4967535528071964e-12
C7_38 V7 V38 3.554593371389426e-19

R7_39 V7 V39 23595.989272144365
L7_39 V7 V39 -2.965671255557071e-12
C7_39 V7 V39 -4.652038292818435e-19

R7_40 V7 V40 -15506.637630658464
L7_40 V7 V40 2.0378428065785686e-11
C7_40 V7 V40 -1.9790541708625001e-19

R7_41 V7 V41 -20420.071939106332
L7_41 V7 V41 -1.9153338701303493e-12
C7_41 V7 V41 -3.5237132701538785e-19

R7_42 V7 V42 -2848875.3661584733
L7_42 V7 V42 -7.801190921449416e-12
C7_42 V7 V42 -1.2328130222714536e-19

R7_43 V7 V43 7979.260570463837
L7_43 V7 V43 1.2280555279299508e-12
C7_43 V7 V43 5.14561226555748e-19

R7_44 V7 V44 67030.17480421363
L7_44 V7 V44 1.0202662787916518e-11
C7_44 V7 V44 1.4678307254322295e-20

R7_45 V7 V45 -10678.349774547265
L7_45 V7 V45 -1.3895256864235862e-12
C7_45 V7 V45 -2.9877744609577166e-19

R7_46 V7 V46 -6936.872171215334
L7_46 V7 V46 -9.030407011586061e-13
C7_46 V7 V46 -6.061540333152657e-19

R7_47 V7 V47 -6394.427163457192
L7_47 V7 V47 -1.4308023500934472e-12
C7_47 V7 V47 -1.3244231693032009e-19

R7_48 V7 V48 -21513.450573047015
L7_48 V7 V48 -9.467352499145564e-13
C7_48 V7 V48 -4.013340871374001e-19

R7_49 V7 V49 -20047.59962108916
L7_49 V7 V49 5.429373743207868e-12
C7_49 V7 V49 3.72842708661237e-20

R7_50 V7 V50 64465.62884979276
L7_50 V7 V50 1.5662604331683361e-12
C7_50 V7 V50 2.841616933248575e-19

R7_51 V7 V51 -23789.719192313158
L7_51 V7 V51 -1.7985029853777677e-12
C7_51 V7 V51 -3.066934223395397e-19

R7_52 V7 V52 33630.65667451577
L7_52 V7 V52 4.584502425111052e-12
C7_52 V7 V52 2.262655480384663e-19

R7_53 V7 V53 23191.742186649313
L7_53 V7 V53 1.88691373377504e-12
C7_53 V7 V53 3.2833569547656476e-19

R7_54 V7 V54 9320.277394503471
L7_54 V7 V54 1.2504732645061758e-12
C7_54 V7 V54 4.1395260636308763e-19

R7_55 V7 V55 8511.591445091195
L7_55 V7 V55 2.0253165036428954e-12
C7_55 V7 V55 3.550380547415306e-19

R7_56 V7 V56 13415.533706325354
L7_56 V7 V56 1.0918250070607747e-12
C7_56 V7 V56 3.9196132228366434e-19

R7_57 V7 V57 -210029.0894996889
L7_57 V7 V57 1.764419435422104e-11
C7_57 V7 V57 -5.289701846551427e-20

R7_58 V7 V58 -20299.529974661487
L7_58 V7 V58 -2.298931915414499e-12
C7_58 V7 V58 -2.52906826039601e-19

R7_59 V7 V59 36959.942437298945
L7_59 V7 V59 2.2802120916251594e-12
C7_59 V7 V59 2.1247854987613665e-20

R7_60 V7 V60 -10603.253705538407
L7_60 V7 V60 -2.575483044571188e-12
C7_60 V7 V60 -5.025298249591655e-19

R7_61 V7 V61 -20924.35674025521
L7_61 V7 V61 -1.7988521905191222e-12
C7_61 V7 V61 -3.012346946841605e-19

R7_62 V7 V62 -20822.337383731836
L7_62 V7 V62 -3.197833315230839e-12
C7_62 V7 V62 -2.4234887368360245e-19

R7_63 V7 V63 80582.17148926947
L7_63 V7 V63 1.6209323686319133e-11
C7_63 V7 V63 6.59930825554693e-20

R7_64 V7 V64 -196729.60084849183
L7_64 V7 V64 -4.180230609128505e-12
C7_64 V7 V64 -1.4906305475164113e-20

R7_65 V7 V65 -13657.53023324492
L7_65 V7 V65 -7.903924979389535e-12
C7_65 V7 V65 -1.2011682458213666e-19

R7_66 V7 V66 -50787.93207174468
L7_66 V7 V66 3.516248103251163e-12
C7_66 V7 V66 3.249139466453598e-20

R7_67 V7 V67 -48101.34031428052
L7_67 V7 V67 -2.9317703969733986e-12
C7_67 V7 V67 -1.933090208020923e-19

R7_68 V7 V68 30923.789947995265
L7_68 V7 V68 -1.5257744220883107e-10
C7_68 V7 V68 1.6052628590603931e-19

R7_69 V7 V69 19385.250737898674
L7_69 V7 V69 1.9616911175948164e-12
C7_69 V7 V69 3.013084182524528e-19

R7_70 V7 V70 20765.24964517838
L7_70 V7 V70 4.386641506643717e-12
C7_70 V7 V70 1.810854939082012e-19

R7_71 V7 V71 -6059.795713469038
L7_71 V7 V71 -2.358132500291639e-12
C7_71 V7 V71 -1.8457681033575805e-19

R7_72 V7 V72 -77913.52419508372
L7_72 V7 V72 -3.0154824654786534e-12
C7_72 V7 V72 -1.8944810024440256e-19

R7_73 V7 V73 -27988.977452566094
L7_73 V7 V73 -4.473771163266771e-12
C7_73 V7 V73 -1.3465087242195095e-19

R7_74 V7 V74 77242.46874707946
L7_74 V7 V74 -3.318019212878337e-11
C7_74 V7 V74 -2.4828508429353372e-20

R7_75 V7 V75 5632.081856515955
L7_75 V7 V75 1.155311505385605e-12
C7_75 V7 V75 5.262423515592139e-19

R7_76 V7 V76 187312.6969008234
L7_76 V7 V76 1.4841007691290343e-12
C7_76 V7 V76 1.2183727908650537e-19

R7_77 V7 V77 -97919.69956533714
L7_77 V7 V77 4.287817685784928e-11
C7_77 V7 V77 -2.3675708577412043e-20

R7_78 V7 V78 85523.6399547144
L7_78 V7 V78 1.5110103614009666e-11
C7_78 V7 V78 1.536646096386837e-19

R7_79 V7 V79 -71582.9994590376
L7_79 V7 V79 -2.0101950737689675e-12
C7_79 V7 V79 -4.014877318184283e-19

R7_80 V7 V80 -68254.54830822338
L7_80 V7 V80 -3.3999644331464565e-12
C7_80 V7 V80 3.667118235167149e-20

R7_81 V7 V81 -15989.962297749576
L7_81 V7 V81 -5.533557240698921e-12
C7_81 V7 V81 -5.773917836570882e-20

R7_82 V7 V82 -12612.724798357249
L7_82 V7 V82 -2.593263641623876e-12
C7_82 V7 V82 -3.4329428438304827e-19

R7_83 V7 V83 136445.02663568963
L7_83 V7 V83 -6.838022480284764e-12
C7_83 V7 V83 1.0863522872843423e-19

R7_84 V7 V84 -125327.17479595241
L7_84 V7 V84 -1.8179696469047931e-12
C7_84 V7 V84 -1.970349784766881e-19

R7_85 V7 V85 -20360.398631025302
L7_85 V7 V85 -2.0599761006192748e-12
C7_85 V7 V85 -2.1847788499262276e-19

R7_86 V7 V86 -24643.591156221006
L7_86 V7 V86 -2.350471152044121e-12
C7_86 V7 V86 -1.8257903168850717e-19

R7_87 V7 V87 8184.830496301858
L7_87 V7 V87 9.477098493899522e-13
C7_87 V7 V87 7.365130854991339e-19

R7_88 V7 V88 12914.874904455057
L7_88 V7 V88 1.989181949449622e-12
C7_88 V7 V88 2.059833867784497e-19

R7_89 V7 V89 12452.361470122682
L7_89 V7 V89 1.6275362720914872e-12
C7_89 V7 V89 3.013902525965061e-19

R7_90 V7 V90 4267.038494330913
L7_90 V7 V90 5.931508640237661e-13
C7_90 V7 V90 8.796720097468328e-19

R7_91 V7 V91 -3303.2795604645285
L7_91 V7 V91 -4.283407046323624e-13
C7_91 V7 V91 -1.459868669481736e-18

R7_92 V7 V92 -32324.660839199318
L7_92 V7 V92 -1.487499671868585e-12
C7_92 V7 V92 -1.0812321646810901e-19

R7_93 V7 V93 521473.04103379644
L7_93 V7 V93 2.974692232256309e-12
C7_93 V7 V93 2.043789098372322e-19

R7_94 V7 V94 -13733.866159798978
L7_94 V7 V94 -3.288137001439311e-12
C7_94 V7 V94 -2.3806133851211247e-19

R7_95 V7 V95 23075.277834151842
L7_95 V7 V95 2.1581397201688134e-12
C7_95 V7 V95 -3.8147701155046335e-20

R7_96 V7 V96 -10810.03685832482
L7_96 V7 V96 5.02309231705809e-12
C7_96 V7 V96 -1.4589582899323762e-19

R7_97 V7 V97 -6404.151691176023
L7_97 V7 V97 -1.0928472321481382e-12
C7_97 V7 V97 -6.4790695789086015e-19

R7_98 V7 V98 -7381.854433949149
L7_98 V7 V98 -9.141121778783249e-13
C7_98 V7 V98 -6.1078476950177045e-19

R7_99 V7 V99 3088.188874046969
L7_99 V7 V99 4.449875088087336e-13
C7_99 V7 V99 1.7077686624424272e-18

R7_100 V7 V100 6641.634215139418
L7_100 V7 V100 2.6789081511435946e-12
C7_100 V7 V100 2.192346661957682e-19

R7_101 V7 V101 22419.137111200263
L7_101 V7 V101 2.412468880556071e-12
C7_101 V7 V101 1.994878813221542e-19

R7_102 V7 V102 9007.911521255646
L7_102 V7 V102 1.5363439292933155e-12
C7_102 V7 V102 3.678504449941973e-19

R7_103 V7 V103 -12496.262401945278
L7_103 V7 V103 -7.132393327484035e-13
C7_103 V7 V103 -8.167688083576915e-19

R7_104 V7 V104 -29319.106519628116
L7_104 V7 V104 -1.9459709577908864e-12
C7_104 V7 V104 -6.797403958290945e-20

R7_105 V7 V105 250221.96777189072
L7_105 V7 V105 2.4325827061675326e-12
C7_105 V7 V105 3.5730680280827145e-19

R7_106 V7 V106 11427.915376919047
L7_106 V7 V106 1.233358984905042e-12
C7_106 V7 V106 5.997756025983588e-19

R7_107 V7 V107 -4994.155155653302
L7_107 V7 V107 -1.5480919398616429e-12
C7_107 V7 V107 -6.005632202789046e-19

R7_108 V7 V108 -32240.133142821665
L7_108 V7 V108 4.151386607615255e-12
C7_108 V7 V108 -7.155148318248487e-21

R7_109 V7 V109 -15562.449590662482
L7_109 V7 V109 -1.7428420232307225e-12
C7_109 V7 V109 -4.769703610002275e-19

R7_110 V7 V110 -11234.603984170095
L7_110 V7 V110 -1.8889390753019138e-12
C7_110 V7 V110 -4.700747417222244e-19

R7_111 V7 V111 -10243.289545170395
L7_111 V7 V111 -2.501223549772953e-11
C7_111 V7 V111 3.775559065221037e-20

R7_112 V7 V112 12636.276410113725
L7_112 V7 V112 -6.758484096437344e-12
C7_112 V7 V112 1.6019859134979065e-19

R7_113 V7 V113 -16302.848001067112
L7_113 V7 V113 -6.310775134946654e-12
C7_113 V7 V113 -1.3116076498275262e-19

R7_114 V7 V114 -13603.169230232832
L7_114 V7 V114 -1.3024219948848752e-12
C7_114 V7 V114 -5.504478700827732e-19

R7_115 V7 V115 4216.142771981562
L7_115 V7 V115 6.09269587156436e-13
C7_115 V7 V115 5.743397016885663e-19

R7_116 V7 V116 -32712.5400282305
L7_116 V7 V116 3.4150063804220994e-12
C7_116 V7 V116 -1.0891838624660693e-19

R7_117 V7 V117 24982.928632139683
L7_117 V7 V117 1.1505384703797275e-12
C7_117 V7 V117 3.6718589446439376e-19

R7_118 V7 V118 8237.97075629689
L7_118 V7 V118 1.1758431070594016e-12
C7_118 V7 V118 7.500006204117339e-19

R7_119 V7 V119 -47926.42430297939
L7_119 V7 V119 -8.846896770929418e-12
C7_119 V7 V119 5.107782754522997e-20

R7_120 V7 V120 10838.137875511726
L7_120 V7 V120 2.640038978921719e-12
C7_120 V7 V120 2.2647942541478116e-19

R7_121 V7 V121 -22878.617610950634
L7_121 V7 V121 -3.5732318764582487e-12
C7_121 V7 V121 -2.176744740267271e-19

R7_122 V7 V122 -18077.16862303784
L7_122 V7 V122 -7.346204154048389e-12
C7_122 V7 V122 -1.7409561491423693e-19

R7_123 V7 V123 -3534.5728324566057
L7_123 V7 V123 -5.245481564667339e-13
C7_123 V7 V123 -1.0708588212268963e-18

R7_124 V7 V124 -11825.836483578409
L7_124 V7 V124 -1.0613899312250177e-12
C7_124 V7 V124 -1.1015511404726476e-19

R7_125 V7 V125 -28660.406656312036
L7_125 V7 V125 -1.6706703892334485e-12
C7_125 V7 V125 -1.1865241624438197e-20

R7_126 V7 V126 -10100.64620354646
L7_126 V7 V126 -9.272292451527552e-13
C7_126 V7 V126 -5.363710116959512e-19

R7_127 V7 V127 6935.94986695508
L7_127 V7 V127 7.44362993784458e-13
C7_127 V7 V127 6.678853084852836e-19

R7_128 V7 V128 -12553.1252343642
L7_128 V7 V128 8.310949355967902e-12
C7_128 V7 V128 -3.5013936143713295e-19

R7_129 V7 V129 -10160.673426313188
L7_129 V7 V129 -1.4392925492613937e-11
C7_129 V7 V129 -3.506520349033296e-19

R7_130 V7 V130 7649.415475719043
L7_130 V7 V130 1.1343145080230108e-12
C7_130 V7 V130 4.594174755706903e-19

R7_131 V7 V131 16348.612909566262
L7_131 V7 V131 -1.741439466208043e-11
C7_131 V7 V131 8.562879292180911e-20

R7_132 V7 V132 5254.011907796652
L7_132 V7 V132 1.2962060932373986e-12
C7_132 V7 V132 7.309355239264189e-19

R7_133 V7 V133 6950.29873277584
L7_133 V7 V133 1.0626015858225155e-12
C7_133 V7 V133 3.7704051555909615e-19

R7_134 V7 V134 -25638.997640213485
L7_134 V7 V134 -3.8518555136130405e-12
C7_134 V7 V134 -1.994178560983764e-19

R7_135 V7 V135 -3609.6079873991403
L7_135 V7 V135 -5.812157628773976e-13
C7_135 V7 V135 -1.3315984467196335e-18

R7_136 V7 V136 88935.27913900962
L7_136 V7 V136 -2.333103311297496e-12
C7_136 V7 V136 7.128872125241366e-20

R7_137 V7 V137 23328.152095778732
L7_137 V7 V137 3.200960560569036e-11
C7_137 V7 V137 3.1810383577762394e-19

R7_138 V7 V138 -14033.664525191956
L7_138 V7 V138 -1.613445077963653e-12
C7_138 V7 V138 -1.9088962437519868e-19

R7_139 V7 V139 2887.511391419848
L7_139 V7 V139 3.5572702260346136e-13
C7_139 V7 V139 1.8855738625694007e-18

R7_140 V7 V140 -51489.268976139945
L7_140 V7 V140 2.6811586916770556e-12
C7_140 V7 V140 -2.4323016864608154e-19

R7_141 V7 V141 -4477.661974887428
L7_141 V7 V141 -6.286533991143589e-13
C7_141 V7 V141 -8.831581856646342e-19

R7_142 V7 V142 34047.974716858575
L7_142 V7 V142 1.533226015176666e-12
C7_142 V7 V142 5.700929374888331e-20

R7_143 V7 V143 -4967.712620760644
L7_143 V7 V143 -1.5006986758435363e-12
C7_143 V7 V143 -5.791342534228681e-19

R7_144 V7 V144 -6822.85893599473
L7_144 V7 V144 -1.0573708552053853e-11
C7_144 V7 V144 -8.491882004646345e-20

R7_145 V7 V145 -6827.20947292399
L7_145 V7 V145 -9.295568429016037e-12
C7_145 V7 V145 -3.729278641712424e-19

R7_146 V7 V146 -107226.22739571852
L7_146 V7 V146 -5.79149275187486e-12
C7_146 V7 V146 2.0578038940054816e-19

R7_147 V7 V147 21853.687849491773
L7_147 V7 V147 -5.675243759460023e-13
C7_147 V7 V147 -9.728103909086506e-19

R7_148 V7 V148 4814.388048514558
L7_148 V7 V148 -1.8598924136960214e-12
C7_148 V7 V148 8.826959586517887e-20

R7_149 V7 V149 2552.3938136819356
L7_149 V7 V149 4.024808654651458e-13
C7_149 V7 V149 1.3618860261795751e-18

R7_150 V7 V150 -11449.710708204313
L7_150 V7 V150 -1.4937892172677174e-12
C7_150 V7 V150 -5.156107885782973e-19

R7_151 V7 V151 -4871.234565172002
L7_151 V7 V151 1.0614119912967906e-11
C7_151 V7 V151 3.8131085073561913e-19

R7_152 V7 V152 -12172.699554371617
L7_152 V7 V152 7.846707719210906e-12
C7_152 V7 V152 -1.2981603019052427e-19

R7_153 V7 V153 -1276110.3686016023
L7_153 V7 V153 -2.2916630228554e-11
C7_153 V7 V153 7.399367932839969e-20

R7_154 V7 V154 34560.41947547212
L7_154 V7 V154 2.3693898658691286e-12
C7_154 V7 V154 2.6811288644414316e-19

R7_155 V7 V155 1261.1235863592944
L7_155 V7 V155 3.964591104537667e-13
C7_155 V7 V155 1.2273816183849235e-18

R7_156 V7 V156 26658.957327101492
L7_156 V7 V156 4.304160589208386e-12
C7_156 V7 V156 7.70172906442645e-20

R7_157 V7 V157 -4619.297512758095
L7_157 V7 V157 -5.257327736271105e-13
C7_157 V7 V157 -9.048314438564158e-19

R7_158 V7 V158 16573.942385932307
L7_158 V7 V158 2.776612747625592e-12
C7_158 V7 V158 1.5247406168775959e-19

R7_159 V7 V159 -2848.214585131297
L7_159 V7 V159 -1.3616786015326689e-12
C7_159 V7 V159 -7.552262211003129e-19

R7_160 V7 V160 -15680.375218208479
L7_160 V7 V160 7.266318033937249e-12
C7_160 V7 V160 1.722986275439232e-19

R7_161 V7 V161 -12974.843885442488
L7_161 V7 V161 4.5634385860741965e-12
C7_161 V7 V161 -7.091966511949132e-20

R7_162 V7 V162 16827.082227350304
L7_162 V7 V162 1.6966842316828639e-12
C7_162 V7 V162 2.8481548423075867e-19

R7_163 V7 V163 19346.20903959988
L7_163 V7 V163 -1.0170695029205536e-12
C7_163 V7 V163 3.4439195738336017e-19

R7_164 V7 V164 7313.188378749561
L7_164 V7 V164 -2.189060850267017e-12
C7_164 V7 V164 3.9534777421277726e-20

R7_165 V7 V165 13197.374109175189
L7_165 V7 V165 4.190730143826743e-12
C7_165 V7 V165 3.25213531219692e-19

R7_166 V7 V166 -47330.007786772
L7_166 V7 V166 -1.4035544858066247e-12
C7_166 V7 V166 -2.619662764341491e-19

R7_167 V7 V167 -51472.46024026314
L7_167 V7 V167 2.811475275491384e-12
C7_167 V7 V167 -1.1393508315899874e-19

R7_168 V7 V168 -15242.806114504876
L7_168 V7 V168 5.753135063980452e-12
C7_168 V7 V168 -1.3772407727007056e-19

R7_169 V7 V169 -17426.60515410219
L7_169 V7 V169 -3.7171175984058845e-12
C7_169 V7 V169 -1.6410920394397763e-19

R7_170 V7 V170 -251558.35613070056
L7_170 V7 V170 3.821169631713518e-12
C7_170 V7 V170 2.73365131367166e-19

R7_171 V7 V171 8118.399324793204
L7_171 V7 V171 1.7474629850878408e-12
C7_171 V7 V171 1.1212260008600186e-19

R7_172 V7 V172 -18805.134141268307
L7_172 V7 V172 7.765735744558284e-12
C7_172 V7 V172 3.656611109671706e-20

R7_173 V7 V173 86800.50339065585
L7_173 V7 V173 1.8839104801308116e-12
C7_173 V7 V173 1.6747713131782957e-19

R7_174 V7 V174 35516.37934668439
L7_174 V7 V174 1.4388083139453713e-12
C7_174 V7 V174 -1.447774296319381e-19

R7_175 V7 V175 15412.64623746221
L7_175 V7 V175 1.3361469424701959e-12
C7_175 V7 V175 6.88307832832789e-19

R7_176 V7 V176 5992.614067938257
L7_176 V7 V176 2.493458191340875e-12
C7_176 V7 V176 1.5938485121775265e-19

R7_177 V7 V177 -27299.768321004412
L7_177 V7 V177 -2.109872806828573e-12
C7_177 V7 V177 -9.928879646397969e-20

R7_178 V7 V178 -14455.22611318199
L7_178 V7 V178 -1.163036666878474e-12
C7_178 V7 V178 -1.924196998181657e-19

R7_179 V7 V179 22037.22467821004
L7_179 V7 V179 -9.276461046373374e-13
C7_179 V7 V179 -6.599680360133235e-19

R7_180 V7 V180 -6599.2209722453945
L7_180 V7 V180 -1.0771460234372998e-12
C7_180 V7 V180 -3.3183443663342434e-19

R7_181 V7 V181 -74599.73034593707
L7_181 V7 V181 6.052282580343302e-12
C7_181 V7 V181 -2.193117475805564e-19

R7_182 V7 V182 11824.050537079607
L7_182 V7 V182 1.2301898089801006e-12
C7_182 V7 V182 3.1152909570841835e-19

R7_183 V7 V183 -5467.890580094463
L7_183 V7 V183 -1.4351160656280313e-12
C7_183 V7 V183 -4.072674888272814e-20

R7_184 V7 V184 -18307.12291678034
L7_184 V7 V184 -1.862297224768191e-12
C7_184 V7 V184 -1.300748672426953e-19

R7_185 V7 V185 162557.86191503232
L7_185 V7 V185 9.975332825264283e-12
C7_185 V7 V185 2.2500690412482346e-19

R7_186 V7 V186 -38500.614537635665
L7_186 V7 V186 -5.5374887598984565e-12
C7_186 V7 V186 -3.1029667638640183e-19

R7_187 V7 V187 6795.934464793965
L7_187 V7 V187 6.446217949511374e-13
C7_187 V7 V187 6.160603117851604e-19

R7_188 V7 V188 7451.590396928038
L7_188 V7 V188 6.903842623933325e-13
C7_188 V7 V188 3.9536418704725854e-19

R7_189 V7 V189 20988.628196604335
L7_189 V7 V189 -9.220049529801653e-12
C7_189 V7 V189 4.283697732804198e-20

R7_190 V7 V190 -21159.810408302474
L7_190 V7 V190 -5.273721677431279e-12
C7_190 V7 V190 -1.5360344391292542e-19

R7_191 V7 V191 -25888.869709110855
L7_191 V7 V191 5.38765085685388e-12
C7_191 V7 V191 -4.124557173859475e-19

R7_192 V7 V192 173479.39209599842
L7_192 V7 V192 6.568179967487409e-12
C7_192 V7 V192 5.421931465377778e-20

R7_193 V7 V193 -35766.56359580013
L7_193 V7 V193 1.735202507444752e-11
C7_193 V7 V193 -6.981004247788414e-20

R7_194 V7 V194 -172647.15187344572
L7_194 V7 V194 -6.32969168418555e-12
C7_194 V7 V194 -8.329660157529473e-20

R7_195 V7 V195 24187.2471028054
L7_195 V7 V195 -1.9280506965509836e-12
C7_195 V7 V195 5.510036721756985e-19

R7_196 V7 V196 -4720.788080764853
L7_196 V7 V196 -8.131624490443506e-13
C7_196 V7 V196 -6.515518937816735e-19

R7_197 V7 V197 -6759.646782072732
L7_197 V7 V197 -4.312306540081504e-12
C7_197 V7 V197 -2.5475180380438183e-19

R7_198 V7 V198 16282.317463165955
L7_198 V7 V198 4.3736317039298806e-12
C7_198 V7 V198 1.116894949575335e-19

R7_199 V7 V199 6254.917436226318
L7_199 V7 V199 1.05950852261801e-10
C7_199 V7 V199 1.1522359312535268e-19

R7_200 V7 V200 -17240.567670217108
L7_200 V7 V200 3.584176991683794e-12
C7_200 V7 V200 9.931130965442465e-20

R8_8 V8 0 441.67804479299633
L8_8 V8 0 1.3130728957151281e-13
C8_8 V8 0 5.991408017979055e-18

R8_9 V8 V9 -95690.00453826731
L8_9 V8 V9 -2.769531174489916e-12
C8_9 V8 V9 1.3921230017181007e-19

R8_10 V8 V10 150933.8858988788
L8_10 V8 V10 -1.0220083890512085e-11
C8_10 V8 V10 1.215311537216857e-21

R8_11 V8 V11 -200334.4019556899
L8_11 V8 V11 1.9750109911271643e-11
C8_11 V8 V11 1.1065158845808014e-19

R8_12 V8 V12 -6035.545450360764
L8_12 V8 V12 8.112697190569357e-11
C8_12 V8 V12 5.513371949647942e-19

R8_13 V8 V13 50688.84398890453
L8_13 V8 V13 4.329403653955506e-12
C8_13 V8 V13 2.048868433738595e-19

R8_14 V8 V14 7935.1493591044755
L8_14 V8 V14 1.248077332760583e-12
C8_14 V8 V14 7.04590560233978e-19

R8_15 V8 V15 7746.856855875894
L8_15 V8 V15 1.1429421414849497e-12
C8_15 V8 V15 7.34160181044493e-19

R8_16 V8 V16 5439.294995299441
L8_16 V8 V16 3.7917848395574165e-13
C8_16 V8 V16 1.4107513502386743e-18

R8_17 V8 V17 -39257.96006966103
L8_17 V8 V17 8.400694366809232e-12
C8_17 V8 V17 -1.2528674671514062e-19

R8_18 V8 V18 -18280.781769016074
L8_18 V8 V18 5.3633203459870734e-12
C8_18 V8 V18 -1.2584491340478022e-19

R8_19 V8 V19 -15247.060343452198
L8_19 V8 V19 -7.791317010713524e-12
C8_19 V8 V19 -3.6726774568309694e-19

R8_20 V8 V20 44978.19327846417
L8_20 V8 V20 -3.5766897263129037e-12
C8_20 V8 V20 -1.0043008011355808e-18

R8_21 V8 V21 13586.709031277544
L8_21 V8 V21 1.2496764167194387e-12
C8_21 V8 V21 1.848941036389632e-19

R8_22 V8 V22 95851.3427661058
L8_22 V8 V22 -1.2074143976490321e-11
C8_22 V8 V22 -1.217962685932531e-19

R8_23 V8 V23 15490.256671519775
L8_23 V8 V23 3.0663732928522793e-12
C8_23 V8 V23 1.9804650367130405e-19

R8_24 V8 V24 3455.4248508803953
L8_24 V8 V24 1.8091512049827497e-12
C8_24 V8 V24 3.80575703998073e-19

R8_25 V8 V25 -16494.788013606576
L8_25 V8 V25 -2.12610998482228e-12
C8_25 V8 V25 -1.8728498004286369e-19

R8_26 V8 V26 -12545.493032732451
L8_26 V8 V26 -2.41661209002353e-11
C8_26 V8 V26 -1.7215394627526734e-19

R8_27 V8 V27 -7594.225210186004
L8_27 V8 V27 -2.361354255277702e-12
C8_27 V8 V27 -4.254862334442423e-19

R8_28 V8 V28 -2115.106375015227
L8_28 V8 V28 -7.188465523689798e-13
C8_28 V8 V28 -9.27902975707176e-19

R8_29 V8 V29 -11492.772992285572
L8_29 V8 V29 -1.0956606344392053e-12
C8_29 V8 V29 -4.339705940384824e-19

R8_30 V8 V30 -46399.59187633526
L8_30 V8 V30 -3.4393677895750614e-12
C8_30 V8 V30 -1.5811614721047742e-19

R8_31 V8 V31 -21487.423659262957
L8_31 V8 V31 -3.681620138343727e-12
C8_31 V8 V31 -1.320212312574573e-19

R8_32 V8 V32 -43060.43342096502
L8_32 V8 V32 -3.682980934545831e-12
C8_32 V8 V32 6.953494719320362e-19

R8_33 V8 V33 15342.91187536815
L8_33 V8 V33 1.1788216631057068e-12
C8_33 V8 V33 4.204689206947431e-19

R8_34 V8 V34 25624.087409578162
L8_34 V8 V34 2.3574527145920724e-12
C8_34 V8 V34 -4.74641790899214e-20

R8_35 V8 V35 18060.62973828103
L8_35 V8 V35 1.4078235457987016e-12
C8_35 V8 V35 1.8899197395659884e-19

R8_36 V8 V36 3173.259008224089
L8_36 V8 V36 1.075592100556892e-12
C8_36 V8 V36 8.345562459168414e-19

R8_37 V8 V37 12472.049835438738
L8_37 V8 V37 1.3809542107690132e-12
C8_37 V8 V37 3.3881070383157375e-19

R8_38 V8 V38 13080.563353472502
L8_38 V8 V38 1.4448992711961336e-12
C8_38 V8 V38 4.667054875535239e-19

R8_39 V8 V39 -419615.9153632546
L8_39 V8 V39 5.452836800461009e-12
C8_39 V8 V39 -9.573993239557643e-20

R8_40 V8 V40 9102.995663032556
L8_40 V8 V40 -3.619254955350213e-12
C8_40 V8 V40 -4.740848759896902e-19

R8_41 V8 V41 -12010.210400605167
L8_41 V8 V41 -1.7969915191855155e-12
C8_41 V8 V41 -4.95079902002826e-19

R8_42 V8 V42 -14909.95583705973
L8_42 V8 V42 -5.00206538799734e-12
C8_42 V8 V42 -3.583138209609137e-19

R8_43 V8 V43 -59793.46557136067
L8_43 V8 V43 1.0707606441872996e-11
C8_43 V8 V43 -6.721919639043337e-20

R8_44 V8 V44 6698.999008535819
L8_44 V8 V44 1.5818240348627205e-12
C8_44 V8 V44 6.017810406496833e-19

R8_45 V8 V45 -9492.64077130884
L8_45 V8 V45 -1.3132739622563985e-12
C8_45 V8 V45 -3.9888211957594053e-19

R8_46 V8 V46 -5259.167530805251
L8_46 V8 V46 -8.82546750149003e-13
C8_46 V8 V46 -7.706327421741692e-19

R8_47 V8 V47 -8122.629365755387
L8_47 V8 V47 -1.4463629422801136e-12
C8_47 V8 V47 -3.9585099899975157e-19

R8_48 V8 V48 -2665.586716609114
L8_48 V8 V48 -7.877211018352233e-13
C8_48 V8 V48 -5.33090429490359e-19

R8_49 V8 V49 -39835.00804661599
L8_49 V8 V49 5.5496894615885714e-12
C8_49 V8 V49 -3.735975718392198e-20

R8_50 V8 V50 55383.231431291475
L8_50 V8 V50 1.637240078994275e-12
C8_50 V8 V50 2.396241578274306e-19

R8_51 V8 V51 -25230.043847888675
L8_51 V8 V51 3.4485066162817553e-12
C8_51 V8 V51 4.595516784591127e-20

R8_52 V8 V52 12526.664221295048
L8_52 V8 V52 -4.6542609679539485e-12
C8_52 V8 V52 1.135746513129715e-19

R8_53 V8 V53 16539.846637006973
L8_53 V8 V53 1.9824249833684344e-12
C8_53 V8 V53 3.7175260677958134e-19

R8_54 V8 V54 7352.073935533105
L8_54 V8 V54 1.2565541015327054e-12
C8_54 V8 V54 4.942673538543475e-19

R8_55 V8 V55 16835.13050700646
L8_55 V8 V55 2.0904937686981335e-12
C8_55 V8 V55 2.6461180620586867e-19

R8_56 V8 V56 3251.5637116214693
L8_56 V8 V56 1.1017072874650795e-12
C8_56 V8 V56 9.280515186894442e-19

R8_57 V8 V57 -39519.00933093618
L8_57 V8 V57 1.6421542102941443e-11
C8_57 V8 V57 -2.210602066625649e-19

R8_58 V8 V58 -8483.59203635235
L8_58 V8 V58 -2.0472609554077725e-12
C8_58 V8 V58 -4.493434219627756e-19

R8_59 V8 V59 -8469.3469101526
L8_59 V8 V59 -2.2106758226717984e-12
C8_59 V8 V59 -6.546773186965753e-19

R8_60 V8 V60 15408.80396239074
L8_60 V8 V60 2.892227154203664e-12
C8_60 V8 V60 -5.830548494385673e-20

R8_61 V8 V61 -18820.436100253257
L8_61 V8 V61 -1.713295132565496e-12
C8_61 V8 V61 -2.900674200596318e-19

R8_62 V8 V62 -17600.401852623618
L8_62 V8 V62 -2.9210697998168188e-12
C8_62 V8 V62 -3.490696450055668e-19

R8_63 V8 V63 30569.83846422382
L8_63 V8 V63 4.867974908995707e-12
C8_63 V8 V63 1.8897608395547275e-19

R8_64 V8 V64 -17756.48923004183
L8_64 V8 V64 -2.1428522941968296e-12
C8_64 V8 V64 -6.044895542606799e-20

R8_65 V8 V65 -11794.009854858215
L8_65 V8 V65 -6.813369482853468e-12
C8_65 V8 V65 -2.371640288329366e-19

R8_66 V8 V66 -33043.397298131575
L8_66 V8 V66 3.5351228372372857e-12
C8_66 V8 V66 -1.3962077295676373e-20

R8_67 V8 V67 24326.725239428844
L8_67 V8 V67 1.946332054668608e-12
C8_67 V8 V67 2.7023195238164294e-19

R8_68 V8 V68 -10311.933701275777
L8_68 V8 V68 -1.4029502925901015e-12
C8_68 V8 V68 -3.0294389825270965e-19

R8_69 V8 V69 8731.203389913791
L8_69 V8 V69 1.9592008453104854e-12
C8_69 V8 V69 4.860211531762653e-19

R8_70 V8 V70 9061.019924403889
L8_70 V8 V70 4.152960299400637e-12
C8_70 V8 V70 3.706086132671159e-19

R8_71 V8 V71 -17545.44383611744
L8_71 V8 V71 -1.3547437470386935e-12
C8_71 V8 V71 -3.1555170535139374e-19

R8_72 V8 V72 -8801.850534199442
L8_72 V8 V72 1.9973650920325392e-11
C8_72 V8 V72 1.2020720439403151e-19

R8_73 V8 V73 -18499.98989571336
L8_73 V8 V73 -4.986814913149028e-12
C8_73 V8 V73 -2.7125546662301874e-19

R8_74 V8 V74 -119928.90801084238
L8_74 V8 V74 -2.3447163622153168e-11
C8_74 V8 V74 -1.6350121135907295e-19

R8_75 V8 V75 -14637.317744764217
L8_75 V8 V75 6.102069543439785e-11
C8_75 V8 V75 -2.1737936839990236e-19

R8_76 V8 V76 2815.028684682052
L8_76 V8 V76 6.822894469016236e-13
C8_76 V8 V76 9.602403900047386e-19

R8_77 V8 V77 -37378.71901343379
L8_77 V8 V77 2.187999029128258e-11
C8_77 V8 V77 -1.1957417806175997e-19

R8_78 V8 V78 -138803.3820154522
L8_78 V8 V78 2.4891145846443826e-11
C8_78 V8 V78 2.7074038571348963e-19

R8_79 V8 V79 17437.986295177685
L8_79 V8 V79 2.4466578296100556e-12
C8_79 V8 V79 2.616497758336444e-19

R8_80 V8 V80 -15052.722680011091
L8_80 V8 V80 -9.27484430333551e-13
C8_80 V8 V80 -7.123025189273115e-19

R8_81 V8 V81 -10956.974470308192
L8_81 V8 V81 -3.3391625335146183e-12
C8_81 V8 V81 -2.3773458205646063e-19

R8_82 V8 V82 -10455.395640319104
L8_82 V8 V82 -2.823828170118694e-12
C8_82 V8 V82 -4.718687978718697e-19

R8_83 V8 V83 -24147.78446121518
L8_83 V8 V83 7.410084596181234e-12
C8_83 V8 V83 -1.3600281336327765e-19

R8_84 V8 V84 -6505.927731133433
L8_84 V8 V84 -1.2420913748100415e-12
C8_84 V8 V84 -2.1999113633019755e-19

R8_85 V8 V85 -20087.08043264996
L8_85 V8 V85 -2.3215657273146114e-12
C8_85 V8 V85 -2.1102675607043598e-19

R8_86 V8 V86 -10255.092620390567
L8_86 V8 V86 -2.8199528038708098e-12
C8_86 V8 V86 -3.3238318238461483e-19

R8_87 V8 V87 29793.62043873208
L8_87 V8 V87 6.5950315295460284e-12
C8_87 V8 V87 1.917804134345364e-19

R8_88 V8 V88 6017.188063769878
L8_88 V8 V88 6.973891694838149e-13
C8_88 V8 V88 1.0636489455886644e-18

R8_89 V8 V89 8137.894108329241
L8_89 V8 V89 1.4022140723392791e-12
C8_89 V8 V89 4.355475858293643e-19

R8_90 V8 V90 3821.676302319968
L8_90 V8 V90 6.191487789719648e-13
C8_90 V8 V90 9.75099119296294e-19

R8_91 V8 V91 -6548.769040039107
L8_91 V8 V91 -1.1669579963002768e-12
C8_91 V8 V91 -5.725650212872233e-19

R8_92 V8 V92 -4996.373969909014
L8_92 V8 V92 -4.818890670551187e-13
C8_92 V8 V92 -1.1806714080907793e-18

R8_93 V8 V93 -73049.6712591114
L8_93 V8 V93 3.231687681805599e-12
C8_93 V8 V93 1.1730237323447473e-19

R8_94 V8 V94 -9895.869633567001
L8_94 V8 V94 -3.1883965935992486e-12
C8_94 V8 V94 -3.8039874767271656e-19

R8_95 V8 V95 -485939.0214068957
L8_95 V8 V95 1.1875836845171853e-11
C8_95 V8 V95 -9.970233968456134e-20

R8_96 V8 V96 10124.144293134965
L8_96 V8 V96 1.3187526799358283e-12
C8_96 V8 V96 -1.6441830521096993e-19

R8_97 V8 V97 -5386.830595559575
L8_97 V8 V97 -1.0764287666761257e-12
C8_97 V8 V97 -1.073775801024878e-18

R8_98 V8 V98 -5204.106703811789
L8_98 V8 V98 -9.121931701448028e-13
C8_98 V8 V98 -7.956186650893183e-19

R8_99 V8 V99 7487.118809964353
L8_99 V8 V99 7.80351473967401e-13
C8_99 V8 V99 5.6738471991498025e-19

R8_100 V8 V100 5012.2075868903
L8_100 V8 V100 8.959900473529128e-13
C8_100 V8 V100 1.7007375515593149e-18

R8_101 V8 V101 204405.7629562981
L8_101 V8 V101 2.324317981972925e-12
C8_101 V8 V101 2.0750797301692665e-19

R8_102 V8 V102 8319.469920014279
L8_102 V8 V102 1.4550974700149475e-12
C8_102 V8 V102 4.735087468071938e-19

R8_103 V8 V103 -13085.472913131605
L8_103 V8 V103 -3.2720132806191027e-12
C8_103 V8 V103 -1.7580868322287035e-19

R8_104 V8 V104 -6941.53824227047
L8_104 V8 V104 -6.835476848586722e-13
C8_104 V8 V104 -1.0511750049578147e-18

R8_105 V8 V105 18458.96047447741
L8_105 V8 V105 2.366883516132056e-12
C8_105 V8 V105 4.4496336831710245e-19

R8_106 V8 V106 11035.259962318367
L8_106 V8 V106 1.6548753700750663e-12
C8_106 V8 V106 6.66443035627251e-19

R8_107 V8 V107 -7759.038406920654
L8_107 V8 V107 -1.4138482776123693e-12
C8_107 V8 V107 -4.807305361358926e-19

R8_108 V8 V108 -53588.43653901919
L8_108 V8 V108 1.2754427287248583e-12
C8_108 V8 V108 -2.497567556672649e-20

R8_109 V8 V109 -11384.313385145935
L8_109 V8 V109 -1.7829746635178935e-12
C8_109 V8 V109 -7.384041046752556e-19

R8_110 V8 V110 -79536.54431740909
L8_110 V8 V110 -3.2821836928887793e-12
C8_110 V8 V110 -2.973855151365227e-19

R8_111 V8 V111 37423.05423687033
L8_111 V8 V111 -1.1549770519788797e-11
C8_111 V8 V111 2.0968597057250386e-19

R8_112 V8 V112 -3553.49399465397
L8_112 V8 V112 -1.154490254040478e-12
C8_112 V8 V112 -5.170020156881576e-19

R8_113 V8 V113 -20984.721942833203
L8_113 V8 V113 -4.30158544605649e-12
C8_113 V8 V113 -1.0537913550063995e-19

R8_114 V8 V114 -11393.299431134563
L8_114 V8 V114 -1.2722320125377121e-12
C8_114 V8 V114 -6.675803930825721e-19

R8_115 V8 V115 5486.167203095197
L8_115 V8 V115 1.336955263348021e-12
C8_115 V8 V115 2.9423139742989564e-19

R8_116 V8 V116 3860.880965588726
L8_116 V8 V116 1.0863460321971766e-12
C8_116 V8 V116 3.6725854803763215e-19

R8_117 V8 V117 9264.893907350319
L8_117 V8 V117 1.1711429749804347e-12
C8_117 V8 V117 4.705123539968479e-19

R8_118 V8 V118 10606.814071454104
L8_118 V8 V118 1.6993503382148462e-12
C8_118 V8 V118 8.067617326563455e-19

R8_119 V8 V119 22961.53282794245
L8_119 V8 V119 7.421558322697915e-12
C8_119 V8 V119 4.0079097131626294e-19

R8_120 V8 V120 10857.91167508878
L8_120 V8 V120 1.441452402441425e-12
C8_120 V8 V120 1.0687309195161105e-18

R8_121 V8 V121 -16621.589734270954
L8_121 V8 V121 -4.225229164184063e-12
C8_121 V8 V121 -3.2670004686850457e-19

R8_122 V8 V122 170134.6408664816
L8_122 V8 V122 -1.7421484505124685e-10
C8_122 V8 V122 5.712108328547205e-20

R8_123 V8 V123 -7379.6455848800615
L8_123 V8 V123 -1.4207446362317592e-12
C8_123 V8 V123 -3.253701125841247e-19

R8_124 V8 V124 -2229.017636397958
L8_124 V8 V124 -3.8767663803126356e-13
C8_124 V8 V124 -2.1155700600572778e-18

R8_125 V8 V125 -13982.578212596509
L8_125 V8 V125 -1.443908357978273e-12
C8_125 V8 V125 -3.307370968362496e-20

R8_126 V8 V126 -11555.81656388633
L8_126 V8 V126 -9.613262495491364e-13
C8_126 V8 V126 -5.039134923995057e-19

R8_127 V8 V127 -62124.657216546555
L8_127 V8 V127 -2.203903693042173e-12
C8_127 V8 V127 -5.26509041578909e-19

R8_128 V8 V128 5784.990717131424
L8_128 V8 V128 7.648173640436651e-13
C8_128 V8 V128 3.5628612460494137e-19

R8_129 V8 V129 -31474.452144800347
L8_129 V8 V129 -6.070070604613236e-11
C8_129 V8 V129 -4.235259057196751e-19

R8_130 V8 V130 5672.596713704025
L8_130 V8 V130 1.18327056134508e-12
C8_130 V8 V130 5.579045634738385e-19

R8_131 V8 V131 19388.175668188378
L8_131 V8 V131 1.5320426829273199e-12
C8_131 V8 V131 6.944184328801726e-19

R8_132 V8 V132 8507.367586915696
L8_132 V8 V132 1.8368227337917148e-12
C8_132 V8 V132 9.85902297929314e-19

R8_133 V8 V133 4902.42318034596
L8_133 V8 V133 1.0108061905807547e-12
C8_133 V8 V133 7.127682469523378e-19

R8_134 V8 V134 22776.362670917926
L8_134 V8 V134 -6.761798920002709e-12
C8_134 V8 V134 3.120105623550462e-19

R8_135 V8 V135 7978.460218253111
L8_135 V8 V135 9.461075864076466e-12
C8_135 V8 V135 3.319768871911687e-19

R8_136 V8 V136 -2913.453844313258
L8_136 V8 V136 -4.983187578314857e-13
C8_136 V8 V136 -1.6991553768141601e-18

R8_137 V8 V137 151343.66632327816
L8_137 V8 V137 -6.434302437541361e-12
C8_137 V8 V137 1.0431414137157916e-19

R8_138 V8 V138 -13308.546209156759
L8_138 V8 V138 -1.4594199679210613e-12
C8_138 V8 V138 -4.795010568056909e-19

R8_139 V8 V139 109389.9249153612
L8_139 V8 V139 -9.474191709976228e-12
C8_139 V8 V139 -3.240342385945045e-19

R8_140 V8 V140 3046.8614347882335
L8_140 V8 V140 4.676468561154441e-13
C8_140 V8 V140 1.940974083120335e-18

R8_141 V8 V141 -3654.8019272869997
L8_141 V8 V141 -6.330400753358568e-13
C8_141 V8 V141 -9.567257298996264e-19

R8_142 V8 V142 157165.41262600198
L8_142 V8 V142 1.7695236514601402e-12
C8_142 V8 V142 -2.056123148135423e-20

R8_143 V8 V143 -7399.8992870967395
L8_143 V8 V143 -2.0318362790091516e-12
C8_143 V8 V143 -1.5122914038248475e-19

R8_144 V8 V144 8629.465666146394
L8_144 V8 V144 -8.566549777231942e-12
C8_144 V8 V144 -3.0806095004342e-19

R8_145 V8 V145 -52143.43225940718
L8_145 V8 V145 1.959884419933141e-11
C8_145 V8 V145 -1.8152977294673415e-19

R8_146 V8 V146 21578.77848705899
L8_146 V8 V146 6.078288293167195e-11
C8_146 V8 V146 2.995170355290907e-19

R8_147 V8 V147 46091.12774651814
L8_147 V8 V147 -2.221314085805205e-12
C8_147 V8 V147 -2.4920161945241346e-19

R8_148 V8 V148 -1632.65435924077
L8_148 V8 V148 -4.072680691559134e-13
C8_148 V8 V148 -1.2781227725028005e-18

R8_149 V8 V149 4026.0664366331994
L8_149 V8 V149 4.619113674940587e-13
C8_149 V8 V149 1.003779232835629e-18

R8_150 V8 V150 -4468.641659737262
L8_150 V8 V150 -1.1514817095808324e-12
C8_150 V8 V150 -8.052516938960858e-19

R8_151 V8 V151 45650.63467328661
L8_151 V8 V151 2.269345289427116e-12
C8_151 V8 V151 7.542937130842199e-20

R8_152 V8 V152 3468.7460449256414
L8_152 V8 V152 1.2609178884430788e-12
C8_152 V8 V152 3.9259319683999543e-19

R8_153 V8 V153 6028.210253205415
L8_153 V8 V153 2.874288166695067e-12
C8_153 V8 V153 2.9033685485521335e-19

R8_154 V8 V154 5484.62337499496
L8_154 V8 V154 1.2776407510733571e-12
C8_154 V8 V154 3.0792532955434446e-19

R8_155 V8 V155 7017.848030754717
L8_155 V8 V155 1.1039155914694547e-12
C8_155 V8 V155 2.5047673659533107e-19

R8_156 V8 V156 -25557.73672014062
L8_156 V8 V156 1.076836196352553e-12
C8_156 V8 V156 9.280748982449832e-19

R8_157 V8 V157 -2310.4076307234445
L8_157 V8 V157 -4.756359028162203e-13
C8_157 V8 V157 -1.3478510749321452e-18

R8_158 V8 V158 -8004.471020795032
L8_158 V8 V158 5.818562760149068e-12
C8_158 V8 V158 6.92330193650402e-20

R8_159 V8 V159 -5831.733253934491
L8_159 V8 V159 -7.319452652634329e-12
C8_159 V8 V159 1.027777744871756e-20

R8_160 V8 V160 5875.229159447724
L8_160 V8 V160 4.327295669760156e-12
C8_160 V8 V160 -3.5039856366410443e-19

R8_161 V8 V161 71291.27261593558
L8_161 V8 V161 2.104674416804929e-12
C8_161 V8 V161 1.938945069794187e-20

R8_162 V8 V162 26773.16706167936
L8_162 V8 V162 1.6851141130876278e-12
C8_162 V8 V162 1.523836569466806e-19

R8_163 V8 V163 -11570.807153324267
L8_163 V8 V163 -3.5925007077903227e-12
C8_163 V8 V163 -2.3121367411566894e-19

R8_164 V8 V164 -2746.765952623183
L8_164 V8 V164 -9.079120613726855e-13
C8_164 V8 V164 2.477251429940931e-19

R8_165 V8 V165 -24132.830896401156
L8_165 V8 V165 9.960564847024465e-12
C8_165 V8 V165 1.9800071573524767e-19

R8_166 V8 V166 -7916.190467324465
L8_166 V8 V166 -1.3274940394728972e-12
C8_166 V8 V166 -5.324012380612637e-19

R8_167 V8 V167 -8732.983875055239
L8_167 V8 V167 -3.4141674488881586e-11
C8_167 V8 V167 -3.2132321620325174e-20

R8_168 V8 V168 3017.766379460476
L8_168 V8 V168 1.4302375578642894e-12
C8_168 V8 V168 -1.13308560772065e-19

R8_169 V8 V169 -9764.028209191289
L8_169 V8 V169 -6.424365655553597e-12
C8_169 V8 V169 -4.463509856177289e-19

R8_170 V8 V170 150792.3350420677
L8_170 V8 V170 2.1559641994425227e-12
C8_170 V8 V170 2.6301878095002355e-19

R8_171 V8 V171 8007.442963879308
L8_171 V8 V171 1.1617492499782697e-12
C8_171 V8 V171 1.4207001726194562e-19

R8_172 V8 V172 12930.524347236773
L8_172 V8 V172 -4.159946003756907e-12
C8_172 V8 V172 1.5200219684897608e-19

R8_173 V8 V173 10319.539456920502
L8_173 V8 V173 1.9065403866755153e-12
C8_173 V8 V173 3.0050325511349337e-19

R8_174 V8 V174 11502.673396023858
L8_174 V8 V174 1.671236927160539e-12
C8_174 V8 V174 -1.0670757995545051e-19

R8_175 V8 V175 12650.053480564624
L8_175 V8 V175 5.825996822350278e-12
C8_175 V8 V175 2.3358210783200203e-19

R8_176 V8 V176 -26624.777441992577
L8_176 V8 V176 1.474361146079119e-12
C8_176 V8 V176 8.95569086390566e-19

R8_177 V8 V177 -6873.427464629617
L8_177 V8 V177 -2.3574220658815885e-12
C8_177 V8 V177 -1.9047530521104778e-19

R8_178 V8 V178 -11491.098109872575
L8_178 V8 V178 -1.0962382478044995e-12
C8_178 V8 V178 -1.2834561219612563e-19

R8_179 V8 V179 -6179.966192812196
L8_179 V8 V179 -9.60583839511395e-13
C8_179 V8 V179 -4.525429031383968e-19

R8_180 V8 V180 -13288.408980824956
L8_180 V8 V180 -9.218828266425585e-13
C8_180 V8 V180 -9.148486612952704e-19

R8_181 V8 V181 599493.7016490739
L8_181 V8 V181 2.4913513957827493e-11
C8_181 V8 V181 -2.0971875513442277e-19

R8_182 V8 V182 6734.077171153678
L8_182 V8 V182 1.4691041470348433e-12
C8_182 V8 V182 1.8235141846319884e-19

R8_183 V8 V183 -12319.974453896308
L8_183 V8 V183 -1.7185572098890073e-12
C8_183 V8 V183 -1.909656707764814e-19

R8_184 V8 V184 -14957.765509391156
L8_184 V8 V184 -1.467055776679601e-12
C8_184 V8 V184 2.0348042008534517e-19

R8_185 V8 V185 11946.403071984329
L8_185 V8 V185 1.4860194852315914e-11
C8_185 V8 V185 2.4255370666851413e-19

R8_186 V8 V186 -13292.704587017713
L8_186 V8 V186 -3.029041721510694e-12
C8_186 V8 V186 -9.855269479865602e-20

R8_187 V8 V187 5736.713326525499
L8_187 V8 V187 1.6686985251684818e-12
C8_187 V8 V187 5.268056867146427e-19

R8_188 V8 V188 2965.96969287963
L8_188 V8 V188 4.140722026122573e-13
C8_188 V8 V188 4.365905569402747e-19

R8_189 V8 V189 -34717.5008544309
L8_189 V8 V189 -1.3505656819870284e-11
C8_189 V8 V189 3.049407879064391e-20

R8_190 V8 V190 -7617.908987227725
L8_190 V8 V190 -7.1008751386506e-12
C8_190 V8 V190 -3.2630461377359427e-19

R8_191 V8 V191 8472.277786495219
L8_191 V8 V191 8.320996007137637e-13
C8_191 V8 V191 1.2940333665556327e-19

R8_192 V8 V192 -14560.406275557969
L8_192 V8 V192 -9.556753155579962e-13
C8_192 V8 V192 -4.983009943972065e-19

R8_193 V8 V193 20852.306120531128
L8_193 V8 V193 3.3041043027808117e-11
C8_193 V8 V193 -1.0643533238154253e-19

R8_194 V8 V194 -13028.70061196265
L8_194 V8 V194 -3.622976576369541e-12
C8_194 V8 V194 -4.795325326336336e-19

R8_195 V8 V195 -3248.5863235707775
L8_195 V8 V195 -5.62937414815394e-13
C8_195 V8 V195 -9.029662568434824e-19

R8_196 V8 V196 -12836.265464099068
L8_196 V8 V196 1.9002164780004766e-12
C8_196 V8 V196 9.259354413607546e-19

R8_197 V8 V197 -36946.699580604036
L8_197 V8 V197 -4.064563213665055e-12
C8_197 V8 V197 -4.092705050191098e-20

R8_198 V8 V198 -7347.988426427007
L8_198 V8 V198 1.1271328456662445e-11
C8_198 V8 V198 -2.2862672811723376e-19

R8_199 V8 V199 -2879.1749268634803
L8_199 V8 V199 -3.74811868816929e-11
C8_199 V8 V199 -2.331380441697562e-19

R8_200 V8 V200 4024.0418849558423
L8_200 V8 V200 -2.9279396218484916e-11
C8_200 V8 V200 2.858044790600239e-20

R9_9 V9 0 49.43404697720155
L9_9 V9 0 2.415271893611173e-13
C9_9 V9 0 -4.776969280889368e-19

R9_10 V9 V10 -729.1119066815212
L9_10 V9 V10 -3.515006353031899e-12
C9_10 V9 V10 -1.048213894395463e-19

R9_11 V9 V11 -962.3346886827239
L9_11 V9 V11 -4.780780549801041e-12
C9_11 V9 V11 -8.744075152106967e-20

R9_12 V9 V12 -730.2485277294394
L9_12 V9 V12 -3.632631908649036e-12
C9_12 V9 V12 -1.0229424760395363e-19

R9_13 V9 V13 292.72551407818594
L9_13 V9 V13 -2.8396965091223858e-12
C9_13 V9 V13 3.2017456518149517e-19

R9_14 V9 V14 3987.3903639373284
L9_14 V9 V14 4.919581988527352e-11
C9_14 V9 V14 9.772797661615013e-20

R9_15 V9 V15 5556.131936214847
L9_15 V9 V15 1.6211838221292756e-11
C9_15 V9 V15 5.240859808726405e-20

R9_16 V9 V16 3041.2943387904397
L9_16 V9 V16 1.0045760892258451e-11
C9_16 V9 V16 3.496441839549124e-20

R9_17 V9 V17 1148.3179604338382
L9_17 V9 V17 1.0753998966000885e-12
C9_17 V9 V17 2.2741147496562244e-19

R9_18 V9 V18 -9688.92072942849
L9_18 V9 V18 3.6368214871630005e-12
C9_18 V9 V18 2.459031524361601e-20

R9_19 V9 V19 5037.8330660415695
L9_19 V9 V19 4.229690360392429e-12
C9_19 V9 V19 7.808520788252947e-20

R9_20 V9 V20 3229.553834628137
L9_20 V9 V20 3.036206596917383e-12
C9_20 V9 V20 1.2107337348968769e-19

R9_21 V9 V21 148.22623596472943
L9_21 V9 V21 1.4948340459695705e-12
C9_21 V9 V21 -2.738411558892966e-19

R9_22 V9 V22 681.4464303937673
L9_22 V9 V22 5.73632305985576e-12
C9_22 V9 V22 -2.3505314415474448e-20

R9_23 V9 V23 1146.9937738892932
L9_23 V9 V23 8.496560122809046e-12
C9_23 V9 V23 -9.233485480533614e-20

R9_24 V9 V24 844.9818834734012
L9_24 V9 V24 6.526016200965222e-12
C9_24 V9 V24 -1.3045656956600554e-19

R9_25 V9 V25 -201.41108250902928
L9_25 V9 V25 -1.0993671808884471e-12
C9_25 V9 V25 1.526904908863874e-19

R9_26 V9 V26 -1243.8373960218362
L9_26 V9 V26 -3.7535421461132425e-12
C9_26 V9 V26 -3.1598180090216435e-20

R9_27 V9 V27 -2636.0630905762946
L9_27 V9 V27 -3.343405976574389e-12
C9_27 V9 V27 6.513674953799648e-20

R9_28 V9 V28 -1566.773986938294
L9_28 V9 V28 -2.0560692975609115e-12
C9_28 V9 V28 1.121764052901629e-19

R9_29 V9 V29 -193.7288732744302
L9_29 V9 V29 -2.090701657904671e-12
C9_29 V9 V29 4.248268453112759e-20

R9_30 V9 V30 -2241.5981368126204
L9_30 V9 V30 -1.0104220001325538e-11
C9_30 V9 V30 4.3493864910898654e-20

R9_31 V9 V31 -2150.263712011827
L9_31 V9 V31 -1.558120939975906e-11
C9_31 V9 V31 2.1264603969706812e-20

R9_32 V9 V32 -1378.8591962411467
L9_32 V9 V32 -9.241835190822384e-12
C9_32 V9 V32 1.6059697619143467e-20

R9_33 V9 V33 -469.5914109553382
L9_33 V9 V33 -2.3286148422189576e-12
C9_33 V9 V33 -7.688885766193917e-20

R9_34 V9 V34 8285.106530608731
L9_34 V9 V34 -2.5058104666542922e-11
C9_34 V9 V34 2.701731753352099e-20

R9_35 V9 V35 2092.8445705923446
L9_35 V9 V35 7.241093092842005e-11
C9_35 V9 V35 -2.929778243791933e-20

R9_36 V9 V36 1308.6882911243636
L9_36 V9 V36 1.4425460699997464e-11
C9_36 V9 V36 -2.7749710912082494e-20

R9_37 V9 V37 484.94315412084734
L9_37 V9 V37 1.3179045120703464e-12
C9_37 V9 V37 -1.0810291594298617e-19

R9_38 V9 V38 3089.0527307775133
L9_38 V9 V38 4.443204675589893e-12
C9_38 V9 V38 -1.1079504346151798e-19

R9_39 V9 V39 2183.9085225843987
L9_39 V9 V39 3.871792352550002e-12
C9_39 V9 V39 -4.258290915560464e-21

R9_40 V9 V40 1415.603561176078
L9_40 V9 V40 2.655696553631829e-12
C9_40 V9 V40 -4.663094641383943e-22

R9_41 V9 V41 2083.006767154557
L9_41 V9 V41 -6.107127317615078e-12
C9_41 V9 V41 1.1392674163342203e-20

R9_42 V9 V42 2519.284072856005
L9_42 V9 V42 -1.4308237085050855e-10
C9_42 V9 V42 4.80524727543159e-22

R9_43 V9 V43 1710.3141162135344
L9_43 V9 V43 2.741371640134569e-11
C9_43 V9 V43 -3.771011168184528e-20

R9_44 V9 V44 1373.2559713802405
L9_44 V9 V44 -1.1676336014153856e-10
C9_44 V9 V44 -4.9502748053628704e-20

R9_45 V9 V45 -379.92399739400184
L9_45 V9 V45 -1.6725374970703177e-12
C9_45 V9 V45 2.6289261198898747e-20

R9_46 V9 V46 560892.6790298707
L9_46 V9 V46 2.7924594028562852e-11
C9_46 V9 V46 5.964345892119478e-20

R9_47 V9 V47 -1256422.7695644887
L9_47 V9 V47 -9.643312630799034e-12
C9_47 V9 V47 3.5960098158020306e-20

R9_48 V9 V48 -3502.3652436912603
L9_48 V9 V48 -4.095107105809665e-12
C9_48 V9 V48 5.1325389501782185e-20

R9_49 V9 V49 -348.8180768046324
L9_49 V9 V49 4.915881176032369e-12
C9_49 V9 V49 1.9726117360785305e-19

R9_50 V9 V50 4786.59940622865
L9_50 V9 V50 -2.201151329271715e-11
C9_50 V9 V50 1.571820204539527e-20

R9_51 V9 V51 12583.344629387913
L9_51 V9 V51 -1.3376070625420824e-11
C9_51 V9 V51 7.966825579083901e-20

R9_52 V9 V52 2834.815842341711
L9_52 V9 V52 1.1519017714769869e-10
C9_52 V9 V52 1.0240396335848346e-19

R9_53 V9 V53 -725.2241077416555
L9_53 V9 V53 -2.7030468613929178e-12
C9_53 V9 V53 -1.4387932670320092e-19

R9_54 V9 V54 -2390.5299881477767
L9_54 V9 V54 -1.7049666554452295e-11
C9_54 V9 V54 -1.760305485738201e-20

R9_55 V9 V55 -1985.2465779150607
L9_55 V9 V55 -7.913382671389961e-12
C9_55 V9 V55 -3.6064987628308165e-20

R9_56 V9 V56 -3285.4319367310395
L9_56 V9 V56 -2.056524348886143e-11
C9_56 V9 V56 -4.890936379273615e-20

R9_57 V9 V57 -36043.55331341941
L9_57 V9 V57 3.423935677736227e-12
C9_57 V9 V57 -2.6666315452514896e-19

R9_58 V9 V58 1818.4945710349702
L9_58 V9 V58 7.066025402948442e-12
C9_58 V9 V58 -7.16594586638223e-20

R9_59 V9 V59 1069.086197467746
L9_59 V9 V59 3.4249758158840636e-12
C9_59 V9 V59 -5.502633102248409e-20

R9_60 V9 V60 752.9819352145785
L9_60 V9 V60 2.6413305839634086e-12
C9_60 V9 V60 -9.86948490076236e-20

R9_61 V9 V61 1633.2978625983496
L9_61 V9 V61 -1.2001686966043165e-11
C9_61 V9 V61 2.538883148812976e-19

R9_62 V9 V62 18357.47429965928
L9_62 V9 V62 2.247974861972392e-11
C9_62 V9 V62 -2.5731975901456348e-20

R9_63 V9 V63 19681.284221798516
L9_63 V9 V63 9.892411276254075e-12
C9_63 V9 V63 -5.895768074351456e-20

R9_64 V9 V64 -8422.204000109177
L9_64 V9 V64 3.2946511565108865e-11
C9_64 V9 V64 -2.726067595619641e-20

R9_65 V9 V65 -455.7393608194747
L9_65 V9 V65 -2.681417823175469e-12
C9_65 V9 V65 9.205942454349361e-20

R9_66 V9 V66 4041.083255201012
L9_66 V9 V66 2.121604673641611e-11
C9_66 V9 V66 7.212292040189504e-20

R9_67 V9 V67 4745.015609357967
L9_67 V9 V67 -1.5717780481499097e-11
C9_67 V9 V67 1.0479233438349713e-19

R9_68 V9 V68 10838.441679000138
L9_68 V9 V68 -5.149320279884517e-12
C9_68 V9 V68 1.758299621350612e-19

R9_69 V9 V69 -778.9128653588799
L9_69 V9 V69 -4.975176862136845e-11
C9_69 V9 V69 6.85767564462424e-20

R9_70 V9 V70 7241.920353758574
L9_70 V9 V70 -8.643076889129788e-12
C9_70 V9 V70 1.510198172769112e-20

R9_71 V9 V71 25847.7003798838
L9_71 V9 V71 -5.312547760937305e-12
C9_71 V9 V71 5.090203588886107e-20

R9_72 V9 V72 17815.652095478268
L9_72 V9 V72 -6.710744187129634e-12
C9_72 V9 V72 3.814482552507536e-20

R9_73 V9 V73 -1718.8398236401301
L9_73 V9 V73 -2.362656132307145e-12
C9_73 V9 V73 -3.139366585592524e-19

R9_74 V9 V74 -3696.5379438969776
L9_74 V9 V74 -3.926014832859611e-11
C9_74 V9 V74 -1.2041087990485524e-19

R9_75 V9 V75 -4163.4050131886415
L9_75 V9 V75 -2.2809534184896008e-10
C9_75 V9 V75 -1.4017966418475662e-19

R9_76 V9 V76 10149.374131291843
L9_76 V9 V76 8.401559141738508e-12
C9_76 V9 V76 -1.9661386582783764e-19

R9_77 V9 V77 2041.1390316322838
L9_77 V9 V77 1.654159310630001e-12
C9_77 V9 V77 -1.9400469488961035e-20

R9_78 V9 V78 -3692.863597821943
L9_78 V9 V78 -2.9262524719164405e-10
C9_78 V9 V78 -4.5259165632972094e-21

R9_79 V9 V79 10886.927229194685
L9_79 V9 V79 5.7579030755956485e-12
C9_79 V9 V79 4.029220751776928e-20

R9_80 V9 V80 19782.97591829768
L9_80 V9 V80 6.398654991325749e-12
C9_80 V9 V80 8.470506047245045e-20

R9_81 V9 V81 -247.2830608164334
L9_81 V9 V81 -2.623434947267587e-12
C9_81 V9 V81 2.3132907395393023e-19

R9_82 V9 V82 1522.8079758699876
L9_82 V9 V82 7.273156780089411e-12
C9_82 V9 V82 1.0301042398969034e-19

R9_83 V9 V83 910.8552916486437
L9_83 V9 V83 6.140472835737451e-12
C9_83 V9 V83 4.501146172538599e-20

R9_84 V9 V84 943.1262362591223
L9_84 V9 V84 6.652858049159984e-12
C9_84 V9 V84 1.0291351313364456e-19

R9_85 V9 V85 27159.01248990207
L9_85 V9 V85 -3.1796007861554744e-12
C9_85 V9 V85 -1.0302863770054172e-19

R9_86 V9 V86 666.6719507027486
L9_86 V9 V86 4.6612241214331217e-11
C9_86 V9 V86 8.2279015565913e-21

R9_87 V9 V87 2536.333006414601
L9_87 V9 V87 -1.985369430422997e-11
C9_87 V9 V87 -2.9198386456770624e-20

R9_88 V9 V88 2176.840949313791
L9_88 V9 V88 -6.835620764034405e-12
C9_88 V9 V88 -4.508218119230848e-20

R9_89 V9 V89 -1997.0215185593725
L9_89 V9 V89 -2.90947172854152e-12
C9_89 V9 V89 1.0483311749973469e-19

R9_90 V9 V90 -961.2760839334958
L9_90 V9 V90 -7.582664532463774e-12
C9_90 V9 V90 -1.187833116672876e-19

R9_91 V9 V91 -1479.9001871959845
L9_91 V9 V91 -3.686905793208991e-12
C9_91 V9 V91 6.948639806558078e-20

R9_92 V9 V92 -3883.39646903631
L9_92 V9 V92 -8.083716844169808e-12
C9_92 V9 V92 3.528716991873664e-20

R9_93 V9 V93 -466.19927903790955
L9_93 V9 V93 1.9241828747121545e-12
C9_93 V9 V93 -3.724053713371719e-20

R9_94 V9 V94 -1282.6990937684614
L9_94 V9 V94 2.2944972481067905e-11
C9_94 V9 V94 3.386370896615867e-20

R9_95 V9 V95 -5856.982201246701
L9_95 V9 V95 5.522789795024133e-12
C9_95 V9 V95 -2.754995919077454e-20

R9_96 V9 V96 -2784.8017223029597
L9_96 V9 V96 3.9853729307580544e-12
C9_96 V9 V96 -2.4683306530278885e-20

R9_97 V9 V97 -592.5761405445828
L9_97 V9 V97 -3.883489933839663e-12
C9_97 V9 V97 -2.8582260580205783e-19

R9_98 V9 V98 447.58992078500887
L9_98 V9 V98 1.2268683428946774e-11
C9_98 V9 V98 5.831085925503058e-20

R9_99 V9 V99 478.9707055591826
L9_99 V9 V99 5.6354848124124845e-12
C9_99 V9 V99 -3.849713149346565e-20

R9_100 V9 V100 463.69075891175305
L9_100 V9 V100 6.699962236815812e-12
C9_100 V9 V100 -1.3453676673130373e-20

R9_101 V9 V101 1173.686442179661
L9_101 V9 V101 -3.193408613274345e-12
C9_101 V9 V101 2.1419027615867066e-19

R9_102 V9 V102 9365.217022486178
L9_102 V9 V102 1.6181133050721052e-11
C9_102 V9 V102 -6.862683883971166e-20

R9_103 V9 V103 -16805.05186728041
L9_103 V9 V103 -5.4669412452178256e-11
C9_103 V9 V103 -6.899425583382399e-21

R9_104 V9 V104 3674.872508948065
L9_104 V9 V104 -2.853247587460325e-10
C9_104 V9 V104 2.1642017434857424e-20

R9_105 V9 V105 -199.1585917402352
L9_105 V9 V105 -1.090268771745086e-11
C9_105 V9 V105 4.673658343889801e-20

R9_106 V9 V106 3662.9109684311766
L9_106 V9 V106 -3.36137791073439e-11
C9_106 V9 V106 -1.2662257430023292e-20

R9_107 V9 V107 -6853.606360548167
L9_107 V9 V107 -9.896883994347969e-12
C9_107 V9 V107 4.557330538492875e-20

R9_108 V9 V108 -2309.8254272191684
L9_108 V9 V108 -4.498045525412672e-12
C9_108 V9 V108 1.9314262144070754e-20

R9_109 V9 V109 1059.394180428586
L9_109 V9 V109 -4.7054801964964474e-12
C9_109 V9 V109 -2.5769835217475767e-20

R9_110 V9 V110 -44982.875560119515
L9_110 V9 V110 6.332412003253831e-11
C9_110 V9 V110 5.1121414591583324e-20

R9_111 V9 V111 7485.324661268121
L9_111 V9 V111 -1.24465807394957e-11
C9_111 V9 V111 5.195296916400015e-20

R9_112 V9 V112 2776.3366962114064
L9_112 V9 V112 1.9648573596213324e-11
C9_112 V9 V112 2.448960604527066e-20

R9_113 V9 V113 -1550.6169964428816
L9_113 V9 V113 3.67570664675032e-12
C9_113 V9 V113 -4.576322348217973e-21

R9_114 V9 V114 2979.928264120799
L9_114 V9 V114 1.911325106791331e-11
C9_114 V9 V114 -2.0285221494691002e-20

R9_115 V9 V115 2039.3123511711967
L9_115 V9 V115 5.935652004049047e-12
C9_115 V9 V115 -1.0237473930976597e-19

R9_116 V9 V116 3646.4063493861195
L9_116 V9 V116 5.460826167210817e-12
C9_116 V9 V116 -7.976515455766055e-20

R9_117 V9 V117 -469.4273514101902
L9_117 V9 V117 7.246073864252253e-12
C9_117 V9 V117 -2.562889200799539e-19

R9_118 V9 V118 -12421.09911993647
L9_118 V9 V118 -2.9736974858749415e-11
C9_118 V9 V118 -6.848878888823245e-21

R9_119 V9 V119 2617.9901288578726
L9_119 V9 V119 -1.2423014945713744e-11
C9_119 V9 V119 6.901746511774827e-21

R9_120 V9 V120 1389.34857449031
L9_120 V9 V120 -1.201147357245051e-11
C9_120 V9 V120 -1.7814864456303202e-20

R9_121 V9 V121 24875.003575684183
L9_121 V9 V121 -1.5283828378721844e-12
C9_121 V9 V121 2.8849101567133944e-19

R9_122 V9 V122 1968.3234709272542
L9_122 V9 V122 -1.8891437136442778e-11
C9_122 V9 V122 2.596347682352549e-21

R9_123 V9 V123 -2604.680665053065
L9_123 V9 V123 -9.44658706919593e-11
C9_123 V9 V123 2.1570746216394853e-20

R9_124 V9 V124 -1963.9752167287688
L9_124 V9 V124 -4.037431335651393e-11
C9_124 V9 V124 1.0000896717787641e-19

R9_125 V9 V125 -323.60268139347306
L9_125 V9 V125 -2.886538541623758e-12
C9_125 V9 V125 1.0721448958717682e-19

R9_126 V9 V126 6403.227744146809
L9_126 V9 V126 -1.9092252440771057e-11
C9_126 V9 V126 6.19403719691007e-20

R9_127 V9 V127 7656.348955230087
L9_127 V9 V127 1.7675768379855975e-11
C9_127 V9 V127 1.915385416885784e-20

R9_128 V9 V128 -2718.1932258329884
L9_128 V9 V128 -4.642454457376934e-11
C9_128 V9 V128 1.032406371766915e-20

R9_129 V9 V129 2699.312640692348
L9_129 V9 V129 4.4365443175789056e-12
C9_129 V9 V129 -2.229356167239166e-19

R9_130 V9 V130 -4000.0356096753376
L9_130 V9 V130 5.2557792182459205e-12
C9_130 V9 V130 -4.649833555980648e-20

R9_131 V9 V131 18294.062839164613
L9_131 V9 V131 -3.371167489752367e-11
C9_131 V9 V131 -1.613511093305055e-20

R9_132 V9 V132 1044.8861424760441
L9_132 V9 V132 1.523875169078056e-11
C9_132 V9 V132 -6.794650600951644e-20

R9_133 V9 V133 511.456496486001
L9_133 V9 V133 1.885188101578062e-12
C9_133 V9 V133 6.347598836479553e-20

R9_134 V9 V134 788.7231482509125
L9_134 V9 V134 3.713065931675074e-11
C9_134 V9 V134 -2.319049216983436e-20

R9_135 V9 V135 -5523.926385817456
L9_135 V9 V135 1.7843470753905794e-11
C9_135 V9 V135 -5.740152883769496e-21

R9_136 V9 V136 -1713.535941202711
L9_136 V9 V136 1.8261243375936266e-11
C9_136 V9 V136 1.3354647273525428e-20

R9_137 V9 V137 -354.4598685912266
L9_137 V9 V137 3.857374927558418e-12
C9_137 V9 V137 -6.819586627193884e-20

R9_138 V9 V138 -573.9023016103627
L9_138 V9 V138 -1.2066231335303465e-11
C9_138 V9 V138 4.6407518198074986e-20

R9_139 V9 V139 1526.051303691344
L9_139 V9 V139 -8.33366293754271e-12
C9_139 V9 V139 7.047371730085629e-21

R9_140 V9 V140 1859.3177273168437
L9_140 V9 V140 -1.94213216918067e-11
C9_140 V9 V140 -5.2276372183434206e-20

R9_141 V9 V141 680.1648423987941
L9_141 V9 V141 -1.0937472169507687e-12
C9_141 V9 V141 4.4646914616669144e-20

R9_142 V9 V142 750.1404985047365
L9_142 V9 V142 -5.517087957757378e-11
C9_142 V9 V142 -7.474777798209111e-22

R9_143 V9 V143 2338.3539781326494
L9_143 V9 V143 4.244037290261238e-12
C9_143 V9 V143 -2.6856265856044266e-20

R9_144 V9 V144 882.1342846168732
L9_144 V9 V144 2.0694923452697283e-11
C9_144 V9 V144 6.035018945696124e-20

R9_145 V9 V145 -301.0009323334427
L9_145 V9 V145 -2.7486441557942813e-12
C9_145 V9 V145 1.6653132387630967e-19

R9_146 V9 V146 1174.6073291029745
L9_146 V9 V146 1.8901909557448596e-11
C9_146 V9 V146 -2.962297388970707e-20

R9_147 V9 V147 -2772.592994745258
L9_147 V9 V147 -6.672834501236991e-12
C9_147 V9 V147 1.0715751110395838e-19

R9_148 V9 V148 -571.9521402552315
L9_148 V9 V148 -5.791683979409622e-12
C9_148 V9 V148 5.572985579293795e-20

R9_149 V9 V149 187.74923319366607
L9_149 V9 V149 2.0282476472743416e-12
C9_149 V9 V149 -1.1819864288275527e-19

R9_150 V9 V150 -590.2214766223029
L9_150 V9 V150 -9.284395333108618e-12
C9_150 V9 V150 4.652754988402518e-20

R9_151 V9 V151 -681.5689631098834
L9_151 V9 V151 -2.523833550962873e-12
C9_151 V9 V151 -1.4044688398999476e-20

R9_152 V9 V152 1149.3536194438707
L9_152 V9 V152 -2.3665776606668054e-11
C9_152 V9 V152 -2.5685556970963882e-20

R9_153 V9 V153 -258.2602365589074
L9_153 V9 V153 3.166161109508843e-12
C9_153 V9 V153 -1.7586666122785066e-19

R9_154 V9 V154 2174.8409856778535
L9_154 V9 V154 1.0095788516840794e-11
C9_154 V9 V154 -5.0382902328675156e-20

R9_155 V9 V155 377.5883716420832
L9_155 V9 V155 6.752745694143113e-12
C9_155 V9 V155 1.858009637209209e-20

R9_156 V9 V156 -5448.926856949902
L9_156 V9 V156 1.0656649147444017e-11
C9_156 V9 V156 -9.303115127883575e-20

R9_157 V9 V157 -284.9222084901185
L9_157 V9 V157 -7.179384473332604e-12
C9_157 V9 V157 1.3039676073572326e-20

R9_158 V9 V158 1442.6722174203765
L9_158 V9 V158 1.0905717920158528e-11
C9_158 V9 V158 -1.2827331210866867e-20

R9_159 V9 V159 -2503.957049965423
L9_159 V9 V159 2.4416588730249953e-12
C9_159 V9 V159 -9.403127194141536e-20

R9_160 V9 V160 1046.6908072984647
L9_160 V9 V160 3.1353955754428607e-12
C9_160 V9 V160 1.777303030072916e-21

R9_161 V9 V161 -1178.6867123040283
L9_161 V9 V161 -1.0530378826909376e-11
C9_161 V9 V161 2.0847797160538355e-19

R9_162 V9 V162 3747.209956720273
L9_162 V9 V162 8.680248703459965e-12
C9_162 V9 V162 -7.064346071295154e-20

R9_163 V9 V163 684.1684883520146
L9_163 V9 V163 3.982515926115617e-12
C9_163 V9 V163 -2.324945696267868e-20

R9_164 V9 V164 4441.646960530592
L9_164 V9 V164 -5.357810019046501e-10
C9_164 V9 V164 6.987975728898294e-21

R9_165 V9 V165 -367.29635979673606
L9_165 V9 V165 -9.706463550815272e-13
C9_165 V9 V165 -6.73313081764133e-20

R9_166 V9 V166 785.5303576660077
L9_166 V9 V166 -2.1449794530971344e-12
C9_166 V9 V166 8.827167149041356e-20

R9_167 V9 V167 -3620.308029970192
L9_167 V9 V167 -2.4049903019495698e-12
C9_167 V9 V167 7.262932878436784e-20

R9_168 V9 V168 528.2535287613169
L9_168 V9 V168 -2.8399306206325497e-12
C9_168 V9 V168 1.3096248635057954e-19

R9_169 V9 V169 -5868.557685774833
L9_169 V9 V169 3.1929217618352936e-12
C9_169 V9 V169 -7.184591325492254e-20

R9_170 V9 V170 -347.7517252213915
L9_170 V9 V170 1.2369917056988654e-11
C9_170 V9 V170 2.4606155922690113e-20

R9_171 V9 V171 -475.7548038026928
L9_171 V9 V171 -4.312670330308692e-12
C9_171 V9 V171 5.769468225222123e-20

R9_172 V9 V172 -545.0305434383021
L9_172 V9 V172 1.0035152099111452e-10
C9_172 V9 V172 -2.3641306051723673e-20

R9_173 V9 V173 -390.587990995173
L9_173 V9 V173 1.3692147367808168e-12
C9_173 V9 V173 -9.885318413463032e-20

R9_174 V9 V174 456.0193335855871
L9_174 V9 V174 1.582519071776642e-12
C9_174 V9 V174 -1.735717984449797e-19

R9_175 V9 V175 432.18431131618996
L9_175 V9 V175 1.9214910216934573e-12
C9_175 V9 V175 -1.4509057729409578e-19

R9_176 V9 V176 544.9950148379602
L9_176 V9 V176 1.6176613245506014e-12
C9_176 V9 V176 -1.7735845801167784e-19

R9_177 V9 V177 839.5475099069993
L9_177 V9 V177 -2.0309231180627454e-12
C9_177 V9 V177 1.0278063947171872e-19

R9_178 V9 V178 -2857.966558815135
L9_178 V9 V178 -6.859511459737372e-12
C9_178 V9 V178 4.8318621696963314e-20

R9_179 V9 V179 6723.520127520687
L9_179 V9 V179 5.215506561403217e-10
C9_179 V9 V179 4.180079710089717e-20

R9_180 V9 V180 -1682.3009668699483
L9_180 V9 V180 -4.212954476710886e-12
C9_180 V9 V180 8.357188391813184e-20

R9_181 V9 V181 435.39511659946055
L9_181 V9 V181 5.427826557791531e-12
C9_181 V9 V181 1.7659278933160943e-19

R9_182 V9 V182 -992.6929669654787
L9_182 V9 V182 -4.784542661911428e-12
C9_182 V9 V182 9.925647505050511e-21

R9_183 V9 V183 -994.0428146646316
L9_183 V9 V183 -4.508350984577911e-11
C9_183 V9 V183 9.679471872690831e-23

R9_184 V9 V184 -1033.167563585797
L9_184 V9 V184 -4.501994315428542e-12
C9_184 V9 V184 3.3827911514126585e-20

R9_185 V9 V185 -168.23651476164943
L9_185 V9 V185 -3.2127008542056576e-12
C9_185 V9 V185 -1.8262791169045904e-19

R9_186 V9 V186 453.264873037939
L9_186 V9 V186 -2.192324936870375e-12
C9_186 V9 V186 8.292621356737982e-20

R9_187 V9 V187 2424.8592758360915
L9_187 V9 V187 -2.7623968838531528e-12
C9_187 V9 V187 2.0396292526861424e-20

R9_188 V9 V188 1754.1832981417017
L9_188 V9 V188 -3.0033731950218556e-12
C9_188 V9 V188 3.0712781909796664e-20

R9_189 V9 V189 177.63439506731322
L9_189 V9 V189 4.902783435442238e-12
C9_189 V9 V189 -2.40155946287471e-20

R9_190 V9 V190 -2420.996000762706
L9_190 V9 V190 3.6094160295255123e-12
C9_190 V9 V190 -2.111425777066162e-20

R9_191 V9 V191 -592.9599705851997
L9_191 V9 V191 -3.109485096262786e-11
C9_191 V9 V191 1.7442766997883405e-20

R9_192 V9 V192 -844.0687064081092
L9_192 V9 V192 2.5681079541893056e-12
C9_192 V9 V192 -4.072043259287341e-20

R9_193 V9 V193 1817.6413510449631
L9_193 V9 V193 1.7792382962931632e-12
C9_193 V9 V193 -1.0044362566768904e-20

R9_194 V9 V194 -519.8503549257923
L9_194 V9 V194 1.8408822309621844e-12
C9_194 V9 V194 -1.2047284431942723e-19

R9_195 V9 V195 6234.635862102777
L9_195 V9 V195 5.7245372561055536e-12
C9_195 V9 V195 -1.9233427761809252e-20

R9_196 V9 V196 123360.80215009724
L9_196 V9 V196 3.6599124473024724e-12
C9_196 V9 V196 -9.152074330388163e-20

R9_197 V9 V197 -304.12626707840013
L9_197 V9 V197 -4.322661945579166e-12
C9_197 V9 V197 1.2181155974139048e-19

R9_198 V9 V198 640.6404341781799
L9_198 V9 V198 -4.014201583273578e-12
C9_198 V9 V198 2.1124654445162635e-20

R9_199 V9 V199 401.930755040641
L9_199 V9 V199 1.1889212335729066e-11
C9_199 V9 V199 -6.583850845251844e-20

R9_200 V9 V200 444.59779613066235
L9_200 V9 V200 -3.4302623669386598e-12
C9_200 V9 V200 9.330892882197228e-20

R10_10 V10 0 100.06149897077361
L10_10 V10 0 1.2223725916360974e-12
C10_10 V10 0 -6.602213601377321e-19

R10_11 V10 V11 -2027.6805382123514
L10_11 V10 V11 -5.574055233549134e-12
C10_11 V10 V11 -1.0954241723442e-19

R10_12 V10 V12 -1885.9710297434226
L10_12 V10 V12 -5.343018824725683e-12
C10_12 V10 V12 -9.894162353842841e-20

R10_13 V10 V13 1856.8913402017856
L10_13 V10 V13 -1.7334412337849647e-11
C10_13 V10 V13 9.007308531068723e-20

R10_14 V10 V14 663.8243289451442
L10_14 V10 V14 -5.329984688205103e-12
C10_14 V10 V14 2.5838729571977784e-19

R10_15 V10 V15 3711.61656189095
L10_15 V10 V15 1.8196808143181524e-11
C10_15 V10 V15 9.917020927507909e-20

R10_16 V10 V16 3333.789953012465
L10_16 V10 V16 1.3119833248886904e-11
C10_16 V10 V16 8.779617042649503e-20

R10_17 V10 V17 53216.10395865616
L10_17 V10 V17 3.5994747077261445e-12
C10_17 V10 V17 2.629115266793051e-20

R10_18 V10 V18 1672.219517081667
L10_18 V10 V18 1.2113348197344487e-12
C10_18 V10 V18 4.1557865287567025e-19

R10_19 V10 V19 5306.445463995549
L10_19 V10 V19 4.205024150199552e-12
C10_19 V10 V19 1.2061027770779423e-19

R10_20 V10 V20 3789.5670335465243
L10_20 V10 V20 3.3348771457377055e-12
C10_20 V10 V20 1.5923174805372498e-19

R10_21 V10 V21 840.5074918801
L10_21 V10 V21 3.587381098390105e-12
C10_21 V10 V21 -5.651779862714671e-20

R10_22 V10 V22 558.9134502708393
L10_22 V10 V22 -4.49884063937614e-12
C10_22 V10 V22 -4.0368699458770425e-19

R10_23 V10 V23 2800.4034285936164
L10_23 V10 V23 -1.0154746342050108e-11
C10_23 V10 V23 -1.1480981254625678e-19

R10_24 V10 V24 2498.0581595989033
L10_24 V10 V24 -8.037479580678484e-12
C10_24 V10 V24 -1.5343004371311598e-19

R10_25 V10 V25 -1059.2296478545552
L10_25 V10 V25 -2.0524307329166064e-12
C10_25 V10 V25 -2.811536636071258e-20

R10_26 V10 V26 -933.0780237512525
L10_26 V10 V26 -3.1451187565248176e-12
C10_26 V10 V26 -1.2737701522699717e-20

R10_27 V10 V27 -4220.278724257759
L10_27 V10 V27 -6.001418745217475e-12
C10_27 V10 V27 -1.4306784051406767e-20

R10_28 V10 V28 -3382.057005248801
L10_28 V10 V28 -4.0665361212063235e-12
C10_28 V10 V28 -2.98498813128822e-21

R10_29 V10 V29 -1369.4357657323385
L10_29 V10 V29 -9.592003696115196e-12
C10_29 V10 V29 1.9190690814970964e-20

R10_30 V10 V30 -539.0873192883762
L10_30 V10 V30 9.117304540593882e-12
C10_30 V10 V30 2.3028005137632924e-19

R10_31 V10 V31 -2134.3007520496612
L10_31 V10 V31 8.976221414705283e-12
C10_31 V10 V31 6.582113057758555e-20

R10_32 V10 V32 -1798.3666352078487
L10_32 V10 V32 7.748495137828352e-12
C10_32 V10 V32 9.124993334393421e-20

R10_33 V10 V33 -3009.0061764117163
L10_33 V10 V33 -9.087787181660548e-12
C10_33 V10 V33 4.247376194224432e-20

R10_34 V10 V34 1876.2052478253706
L10_34 V10 V34 -3.991872324990358e-12
C10_34 V10 V34 -9.491299811366795e-20

R10_35 V10 V35 2905.2104466025016
L10_35 V10 V35 -4.2998248823439816e-10
C10_35 V10 V35 -1.2857375563101824e-20

R10_36 V10 V36 1763.2265239851358
L10_36 V10 V36 3.782750614577807e-11
C10_36 V10 V36 1.5506237139153986e-20

R10_37 V10 V37 3860.4434445620846
L10_37 V10 V37 6.394795833896997e-12
C10_37 V10 V37 -6.962915611545462e-20

R10_38 V10 V38 1471.4381410528838
L10_38 V10 V38 -7.108606888163433e-12
C10_38 V10 V38 -2.0520626024995122e-19

R10_39 V10 V39 2564.5822746925155
L10_39 V10 V39 -1.0784539192808807e-11
C10_39 V10 V39 -5.653812472190508e-20

R10_40 V10 V40 1815.5559953689738
L10_40 V10 V40 -1.0662434593728787e-11
C10_40 V10 V40 -6.43052482287309e-20

R10_41 V10 V41 -8051.838514886902
L10_41 V10 V41 1.0547471056031626e-11
C10_41 V10 V41 -4.16343629216213e-21

R10_42 V10 V42 1452.087530895531
L10_42 V10 V42 -8.50884766541243e-12
C10_42 V10 V42 5.342057759022186e-20

R10_43 V10 V43 9113.283980521815
L10_43 V10 V43 9.094237968768078e-12
C10_43 V10 V43 3.6921854195427964e-22

R10_44 V10 V44 12416.79122505578
L10_44 V10 V44 7.710472389392024e-12
C10_44 V10 V44 8.604232702585253e-21

R10_45 V10 V45 -2182.3487368426627
L10_45 V10 V45 -5.2261534625585875e-12
C10_45 V10 V45 -1.7874284697234727e-20

R10_46 V10 V46 -1045.8321659824073
L10_46 V10 V46 1.3825414221879305e-12
C10_46 V10 V46 3.092631852209633e-19

R10_47 V10 V47 -5696.918642018627
L10_47 V10 V47 8.34885209744024e-12
C10_47 V10 V47 5.2455591781030966e-20

R10_48 V10 V48 -2695.3597700745927
L10_48 V10 V48 9.276669856079035e-12
C10_48 V10 V48 7.006952669374593e-20

R10_49 V10 V49 -3176.466740299203
L10_49 V10 V49 -2.0095437341137744e-11
C10_49 V10 V49 5.0236664077661835e-20

R10_50 V10 V50 -1414.7997322636736
L10_50 V10 V50 -2.9277901315671202e-12
C10_50 V10 V50 -1.7054529758433978e-19

R10_51 V10 V51 -12436.45353518095
L10_51 V10 V51 -3.449445376896821e-12
C10_51 V10 V51 -7.466008031231546e-20

R10_52 V10 V52 11257.793536888837
L10_52 V10 V52 -2.721069010685876e-12
C10_52 V10 V52 -9.640824208264152e-20

R10_53 V10 V53 -2807.7496476055335
L10_53 V10 V53 -2.3470577208611882e-11
C10_53 V10 V53 8.483934261045605e-20

R10_54 V10 V54 2355.954931247085
L10_54 V10 V54 -2.161133761066881e-12
C10_54 V10 V54 -2.4080728485730113e-19

R10_55 V10 V55 19218.559524134227
L10_55 V10 V55 5.157705242666048e-10
C10_55 V10 V55 3.684038469756627e-20

R10_56 V10 V56 2862.8441296776273
L10_56 V10 V56 -3.8589448104646636e-11
C10_56 V10 V56 4.341921609285693e-20

R10_57 V10 V57 -20564.199626146295
L10_57 V10 V57 7.740110709793143e-12
C10_57 V10 V57 -1.6387905245956183e-19

R10_58 V10 V58 -5334.645525210812
L10_58 V10 V58 3.048350199138453e-12
C10_58 V10 V58 2.8892500032715096e-19

R10_59 V10 V59 3942.928327724938
L10_59 V10 V59 2.89934623750296e-12
C10_59 V10 V59 7.086074738258917e-20

R10_60 V10 V60 2663.067674665038
L10_60 V10 V60 2.0104250825264145e-12
C10_60 V10 V60 1.0820806488483524e-19

R10_61 V10 V61 21935.622442813343
L10_61 V10 V61 -8.081709936669687e-12
C10_61 V10 V61 7.41821517652868e-21

R10_62 V10 V62 1532.2961242139927
L10_62 V10 V62 1.1788052176235307e-11
C10_62 V10 V62 -9.635344686335011e-21

R10_63 V10 V63 -24023.67150300002
L10_63 V10 V63 -9.635293227262161e-12
C10_63 V10 V63 -1.3141011688124215e-19

R10_64 V10 V64 -4402.513193293331
L10_64 V10 V64 -5.686237697363203e-12
C10_64 V10 V64 -1.5242969171207355e-19

R10_65 V10 V65 -2777.5989420815677
L10_65 V10 V65 5.7275770479220145e-12
C10_65 V10 V65 1.5483758698180395e-19

R10_66 V10 V66 -1356.1641934447916
L10_66 V10 V66 -2.3798449712970584e-11
C10_66 V10 V66 -1.4106654319262695e-19

R10_67 V10 V67 100792.04102807374
L10_67 V10 V67 -2.328757214007861e-11
C10_67 V10 V67 1.7180027839821477e-20

R10_68 V10 V68 -7409.830312814827
L10_68 V10 V68 -1.7099696785150092e-11
C10_68 V10 V68 4.253140206988007e-20

R10_69 V10 V69 -31753.450150866003
L10_69 V10 V69 -3.192031456343187e-12
C10_69 V10 V69 -1.8032068312547338e-20

R10_70 V10 V70 -1645.8924313107282
L10_70 V10 V70 2.1911584762785867e-11
C10_70 V10 V70 1.9431709743887234e-19

R10_71 V10 V71 -7944.335742539032
L10_71 V10 V71 2.193774205763952e-11
C10_71 V10 V71 9.248373031921592e-20

R10_72 V10 V72 -9651.643092189548
L10_72 V10 V72 1.0438685179845399e-11
C10_72 V10 V72 1.23494281577527e-19

R10_73 V10 V73 -1747.3262147704945
L10_73 V10 V73 -5.1364925313368165e-12
C10_73 V10 V73 -1.2117571815845744e-19

R10_74 V10 V74 1194.914978740495
L10_74 V10 V74 -3.377011640629936e-12
C10_74 V10 V74 -1.0574178048902823e-19

R10_75 V10 V75 -12316.778989709233
L10_75 V10 V75 -4.4892181606487796e-11
C10_75 V10 V75 -6.324557535828342e-20

R10_76 V10 V76 2835.532582167596
L10_76 V10 V76 -7.860329505939787e-12
C10_76 V10 V76 -1.1098825560633756e-19

R10_77 V10 V77 5002.300543080952
L10_77 V10 V77 2.0885151960088206e-12
C10_77 V10 V77 3.3864819892362936e-20

R10_78 V10 V78 -3529.96599855057
L10_78 V10 V78 3.3421090826398673e-12
C10_78 V10 V78 8.114469102934179e-20

R10_79 V10 V79 3465.614704885099
L10_79 V10 V79 -8.33915681487661e-11
C10_79 V10 V79 8.507552649684977e-21

R10_80 V10 V80 13227.358806547936
L10_80 V10 V80 2.0414878611006703e-11
C10_80 V10 V80 2.1124110994244925e-20

R10_81 V10 V81 -1336.4592284908297
L10_81 V10 V81 -7.0499354440371296e-12
C10_81 V10 V81 8.263244259982325e-20

R10_82 V10 V82 -9700.93360883862
L10_82 V10 V82 5.507898887751059e-12
C10_82 V10 V82 8.094148170600694e-21

R10_83 V10 V83 8058.257143537287
L10_83 V10 V83 6.81872586418502e-12
C10_83 V10 V83 1.4097145447219242e-20

R10_84 V10 V84 365925.6974612286
L10_84 V10 V84 3.2615983090926754e-12
C10_84 V10 V84 8.814670285972887e-20

R10_85 V10 V85 5626.545672968934
L10_85 V10 V85 -1.3174602273146748e-11
C10_85 V10 V85 -1.8079623564348824e-20

R10_86 V10 V86 -1104.3229335171352
L10_86 V10 V86 -3.2061633196747744e-12
C10_86 V10 V86 -1.2644726978702438e-19

R10_87 V10 V87 62725.49478626455
L10_87 V10 V87 7.821218809978868e-11
C10_87 V10 V87 -2.3415546425793885e-20

R10_88 V10 V88 13085.810622422594
L10_88 V10 V88 -8.838134220048767e-12
C10_88 V10 V88 -5.281397956921443e-20

R10_89 V10 V89 -7961.944756651836
L10_89 V10 V89 -3.2726497705121777e-12
C10_89 V10 V89 -2.0992840963905773e-20

R10_90 V10 V90 1096.5354242000924
L10_90 V10 V90 -5.436565403700846e-12
C10_90 V10 V90 9.827511790221367e-20

R10_91 V10 V91 -7697.546964194203
L10_91 V10 V91 -7.893084429711495e-12
C10_91 V10 V91 5.631665091059937e-20

R10_92 V10 V92 14432.24323315523
L10_92 V10 V92 -4.317506998760858e-12
C10_92 V10 V92 2.2702252603392983e-20

R10_93 V10 V93 -1880.658591637961
L10_93 V10 V93 4.68265157592256e-12
C10_93 V10 V93 -3.7171166530817376e-22

R10_94 V10 V94 1494.0556670807503
L10_94 V10 V94 1.920204283805363e-12
C10_94 V10 V94 4.654846189947912e-22

R10_95 V10 V95 18418.851826813203
L10_95 V10 V95 6.047797752854387e-12
C10_95 V10 V95 -1.1373335837228254e-20

R10_96 V10 V96 6644.371036835108
L10_96 V10 V96 3.484549235706433e-12
C10_96 V10 V96 5.980382295482959e-21

R10_97 V10 V97 4251.43100649777
L10_97 V10 V97 4.259629111377464e-12
C10_97 V10 V97 -3.328004125152942e-20

R10_98 V10 V98 -894.7614883595091
L10_98 V10 V98 -5.263829031013565e-12
C10_98 V10 V98 2.7450680658114506e-21

R10_99 V10 V99 1110.1689629941663
L10_99 V10 V99 1.1747409114515608e-10
C10_99 V10 V99 -5.434681844303933e-20

R10_100 V10 V100 1475.4417595569244
L10_100 V10 V100 6.4223886962939705e-12
C10_100 V10 V100 2.777690445436202e-21

R10_101 V10 V101 -3572.5048257934086
L10_101 V10 V101 -3.6732470707029646e-12
C10_101 V10 V101 3.700104261635302e-20

R10_102 V10 V102 1332.3013428656295
L10_102 V10 V102 -2.4866919278777647e-12
C10_102 V10 V102 -7.216352421135267e-20

R10_103 V10 V103 -1859.5153879078557
L10_103 V10 V103 -4.093276653100841e-12
C10_103 V10 V103 -1.7616589031546652e-20

R10_104 V10 V104 -1724.40945866931
L10_104 V10 V104 -4.008068845782701e-12
C10_104 V10 V104 -9.276025398914365e-21

R10_105 V10 V105 -1044.770075020557
L10_105 V10 V105 -3.280373268862866e-12
C10_105 V10 V105 -3.518496303334687e-20

R10_106 V10 V106 -527.3353434165687
L10_106 V10 V106 2.1432033366348457e-12
C10_106 V10 V106 1.0032995141017671e-20

R10_107 V10 V107 -4257.491446385612
L10_107 V10 V107 4.1316157673514584e-12
C10_107 V10 V107 4.996864513816532e-20

R10_108 V10 V108 -21185.981901350613
L10_108 V10 V108 -4.1498096139053544e-11
C10_108 V10 V108 -1.3433685472269256e-20

R10_109 V10 V109 1306.6916592144846
L10_109 V10 V109 1.3699210721771392e-11
C10_109 V10 V109 2.795896453509317e-20

R10_110 V10 V110 609.7538281111822
L10_110 V10 V110 -2.115064277493813e-11
C10_110 V10 V110 1.7453701955049356e-19

R10_111 V10 V111 -450844.76776792505
L10_111 V10 V111 1.3522722137338917e-11
C10_111 V10 V111 1.1591866730416083e-20

R10_112 V10 V112 6037.362224237085
L10_112 V10 V112 2.9885061058711185e-11
C10_112 V10 V112 -2.8475860045036898e-21

R10_113 V10 V113 -1844.10353762568
L10_113 V10 V113 2.530181825867839e-12
C10_113 V10 V113 6.29768971315025e-20

R10_114 V10 V114 702.540598053551
L10_114 V10 V114 -2.2299127431641153e-12
C10_114 V10 V114 -1.8534483605056422e-19

R10_115 V10 V115 1323.2371320467946
L10_115 V10 V115 -3.6119976149375888e-12
C10_115 V10 V115 -6.956913736964985e-20

R10_116 V10 V116 2200.4895870743308
L10_116 V10 V116 -2.335720542775446e-09
C10_116 V10 V116 -1.596848489388519e-20

R10_117 V10 V117 -11403.097190455155
L10_117 V10 V117 -3.620512624036773e-11
C10_117 V10 V117 -1.1944890557547387e-19

R10_118 V10 V118 -344.39233690936237
L10_118 V10 V118 7.690479217899019e-12
C10_118 V10 V118 -9.329204641337865e-22

R10_119 V10 V119 -1901.4116121900465
L10_119 V10 V119 9.437996450662475e-12
C10_119 V10 V119 1.5031534486601524e-20

R10_120 V10 V120 -2959.7020792074995
L10_120 V10 V120 2.7185187439519988e-11
C10_120 V10 V120 -5.4351629753132745e-21

R10_121 V10 V121 -7667.351496720459
L10_121 V10 V121 -1.5352006215521132e-12
C10_121 V10 V121 3.652220964951989e-20

R10_122 V10 V122 6717.145061695807
L10_122 V10 V122 2.584290846610219e-12
C10_122 V10 V122 1.6457242989326028e-19

R10_123 V10 V123 -1461.4727652592176
L10_123 V10 V123 -4.6801799292758296e-11
C10_123 V10 V123 3.5259295761264025e-21

R10_124 V10 V124 -1399.22338284783
L10_124 V10 V124 -5.6576800384219415e-12
C10_124 V10 V124 3.495657396987287e-21

R10_125 V10 V125 -864.8415702055617
L10_125 V10 V125 -3.7687353899379416e-11
C10_125 V10 V125 7.063379616366324e-20

R10_126 V10 V126 679.6289076534584
L10_126 V10 V126 -2.4751070174219523e-12
C10_126 V10 V126 -8.993533740976021e-20

R10_127 V10 V127 822.4812746553876
L10_127 V10 V127 -4.059192219225375e-11
C10_127 V10 V127 1.492518180227319e-20

R10_128 V10 V128 927.4683763669261
L10_128 V10 V128 2.128242236940433e-11
C10_128 V10 V128 1.6771277135996377e-20

R10_129 V10 V129 1059.2016826915253
L10_129 V10 V129 1.5638049717119943e-12
C10_129 V10 V129 9.908073851205688e-21

R10_130 V10 V130 10540.013937041022
L10_130 V10 V130 -6.754598916736452e-12
C10_130 V10 V130 -4.550471643843381e-20

R10_131 V10 V131 -1087.2279049376687
L10_131 V10 V131 9.11132535874987e-12
C10_131 V10 V131 4.086572784357738e-21

R10_132 V10 V132 -1080.0939265060376
L10_132 V10 V132 1.0715422052427717e-11
C10_132 V10 V132 -6.683907348589876e-21

R10_133 V10 V133 1539.0151970543177
L10_133 V10 V133 -3.1299913056017968e-12
C10_133 V10 V133 -7.253169233312124e-20

R10_134 V10 V134 -550.9220090109789
L10_134 V10 V134 1.842319910175023e-12
C10_134 V10 V134 1.303465060916711e-19

R10_135 V10 V135 -1395.7929527617298
L10_135 V10 V135 -4.3429995302063734e-12
C10_135 V10 V135 -3.09639030042076e-20

R10_136 V10 V136 -840.9697693167071
L10_136 V10 V136 -7.05634846086282e-12
C10_136 V10 V136 -3.055515696982754e-20

R10_137 V10 V137 -467.1504401557167
L10_137 V10 V137 -3.3923479023281097e-12
C10_137 V10 V137 -7.03405561379225e-20

R10_138 V10 V138 1248.1862297190767
L10_138 V10 V138 -2.0487936495681563e-12
C10_138 V10 V138 -7.990197506197173e-20

R10_139 V10 V139 653.0499120113823
L10_139 V10 V139 -1.8307359813694108e-11
C10_139 V10 V139 6.7060227717626744e-21

R10_140 V10 V140 637.0569061354349
L10_140 V10 V140 -6.359200953932658e-11
C10_140 V10 V140 3.734827450003312e-21

R10_141 V10 V141 4673.845014830525
L10_141 V10 V141 2.832525022726297e-12
C10_141 V10 V141 1.3850440697338578e-19

R10_142 V10 V142 299.99172967565755
L10_142 V10 V142 -2.516255978141745e-12
C10_142 V10 V142 1.2011198884817392e-20

R10_143 V10 V143 -1503.3119031168874
L10_143 V10 V143 2.638225611812732e-12
C10_143 V10 V143 3.13420400059407e-20

R10_144 V10 V144 1625.9811748111765
L10_144 V10 V144 7.59829521824471e-12
C10_144 V10 V144 5.002572434775212e-20

R10_145 V10 V145 780.5742476487168
L10_145 V10 V145 6.9484406954314304e-12
C10_145 V10 V145 9.89201162689292e-20

R10_146 V10 V146 -236.8456010164591
L10_146 V10 V146 9.610614893203176e-13
C10_146 V10 V146 -1.487953918737087e-20

R10_147 V10 V147 1869.3613403267218
L10_147 V10 V147 -6.9106066488659e-12
C10_147 V10 V147 2.597628875395957e-20

R10_148 V10 V148 -420.229244229063
L10_148 V10 V148 -1.3648586082164733e-11
C10_148 V10 V148 -1.7091075850973337e-20

R10_149 V10 V149 12752.244893230163
L10_149 V10 V149 -1.1427588436407809e-12
C10_149 V10 V149 -2.0520156777397502e-19

R10_150 V10 V150 -557.7886803937649
L10_150 V10 V150 -2.966280542286217e-12
C10_150 V10 V150 8.873521471876392e-20

R10_151 V10 V151 -2823.0548688524077
L10_151 V10 V151 -3.5060231775452596e-12
C10_151 V10 V151 -4.9306993577630804e-20

R10_152 V10 V152 312.67832796527097
L10_152 V10 V152 -2.6304166579071526e-11
C10_152 V10 V152 -3.0855735445222265e-21

R10_153 V10 V153 -486.19593646390575
L10_153 V10 V153 -4.279901821696841e-11
C10_153 V10 V153 -8.301356232844835e-20

R10_154 V10 V154 513.0356257338395
L10_154 V10 V154 -2.358129425279041e-12
C10_154 V10 V154 -1.0179138304756866e-19

R10_155 V10 V155 412.11296822229826
L10_155 V10 V155 -3.4409920242331446e-10
C10_155 V10 V155 2.901809385105481e-20

R10_156 V10 V156 -272.24933783211253
L10_156 V10 V156 2.2457416386728243e-11
C10_156 V10 V156 -1.794685888313531e-20

R10_157 V10 V157 13158.714537096175
L10_157 V10 V157 1.1832983966871466e-12
C10_157 V10 V157 1.3823743844915934e-19

R10_158 V10 V158 1089.8902756690259
L10_158 V10 V158 2.896825628094593e-12
C10_158 V10 V158 4.589653257632256e-20

R10_159 V10 V159 -287.111908524819
L10_159 V10 V159 4.6396041517706105e-12
C10_159 V10 V159 -6.946692885108973e-20

R10_160 V10 V160 -2126.5592696793797
L10_160 V10 V160 1.2495885012067681e-11
C10_160 V10 V160 -3.133310219435136e-20

R10_161 V10 V161 737.3860188900261
L10_161 V10 V161 1.885112063730308e-11
C10_161 V10 V161 1.087696005239344e-19

R10_162 V10 V162 -868.9967308807759
L10_162 V10 V162 5.968925966514125e-12
C10_162 V10 V162 -9.366244137302439e-20

R10_163 V10 V163 607.7726921824288
L10_163 V10 V163 3.74998517013392e-12
C10_163 V10 V163 3.2647627216672955e-20

R10_164 V10 V164 1001.1598507830547
L10_164 V10 V164 -1.4810159843890834e-09
C10_164 V10 V164 6.792094991616242e-21

R10_165 V10 V165 -463.45469328906574
L10_165 V10 V165 -1.182537907988224e-12
C10_165 V10 V165 -1.223390410635132e-19

R10_166 V10 V166 -397.4354847970847
L10_166 V10 V166 -1.261742104460407e-12
C10_166 V10 V166 5.095621702552783e-20

R10_167 V10 V167 -5268.833148860183
L10_167 V10 V167 2.13355699317798e-11
C10_167 V10 V167 3.1310957427713855e-20

R10_168 V10 V168 511.2174631586399
L10_168 V10 V168 4.0422115171263845e-12
C10_168 V10 V168 9.883636837103804e-20

R10_169 V10 V169 -776.3345966999174
L10_169 V10 V169 1.4265008667147112e-11
C10_169 V10 V169 -6.183179134771995e-20

R10_170 V10 V170 443.5397564563051
L10_170 V10 V170 4.288727115070243e-12
C10_170 V10 V170 -3.5640607323287356e-20

R10_171 V10 V171 -1783.1329672843135
L10_171 V10 V171 -1.7059703665351664e-12
C10_171 V10 V171 -5.575079095021911e-20

R10_172 V10 V172 -580.1856924514796
L10_172 V10 V172 -2.4702282994161416e-12
C10_172 V10 V172 -5.808588229995256e-20

R10_173 V10 V173 1190.6032303572858
L10_173 V10 V173 1.6408723480968951e-12
C10_173 V10 V173 2.6007516991917423e-20

R10_174 V10 V174 418.2918996792813
L10_174 V10 V174 1.507115834043697e-12
C10_174 V10 V174 -4.776442808919249e-20

R10_175 V10 V175 8225.351153543763
L10_175 V10 V175 9.112997159821611e-12
C10_175 V10 V175 -7.185953811737766e-20

R10_176 V10 V176 44566.89555437295
L10_176 V10 V176 1.0887430122532037e-11
C10_176 V10 V176 -7.450802719038015e-20

R10_177 V10 V177 -1383.8647082757266
L10_177 V10 V177 -7.2280203674512975e-12
C10_177 V10 V177 2.1948298110134802e-20

R10_178 V10 V178 -325.4264092334231
L10_178 V10 V178 -5.372346115970471e-12
C10_178 V10 V178 8.437777310580149e-20

R10_179 V10 V179 1381.4656422200342
L10_179 V10 V179 1.996251838462949e-12
C10_179 V10 V179 1.1369133425892025e-19

R10_180 V10 V180 8291.749695930603
L10_180 V10 V180 2.1155787411852373e-12
C10_180 V10 V180 8.965985446549034e-20

R10_181 V10 V181 2083.6819797525104
L10_181 V10 V181 -4.9947308185237194e-11
C10_181 V10 V181 6.34061988327021e-20

R10_182 V10 V182 6297.996677178672
L10_182 V10 V182 -1.384142982209568e-12
C10_182 V10 V182 -5.967783113112903e-20

R10_183 V10 V183 -747.4428965414289
L10_183 V10 V183 5.6475931445211655e-12
C10_183 V10 V183 1.1881631153998657e-20

R10_184 V10 V184 -1352.9029911898817
L10_184 V10 V184 -2.0220902540455193e-11
C10_184 V10 V184 2.985397640914005e-20

R10_185 V10 V185 -2733.735051676846
L10_185 V10 V185 -8.28362479303625e-12
C10_185 V10 V185 -5.417888003926397e-20

R10_186 V10 V186 617.7887747590011
L10_186 V10 V186 -4.967862057275981e-12
C10_186 V10 V186 1.2787956343398747e-20

R10_187 V10 V187 1540.1801934000002
L10_187 V10 V187 -1.8984722307277602e-12
C10_187 V10 V187 -4.45832580433191e-20

R10_188 V10 V188 505.032737127527
L10_188 V10 V188 -1.9393844426929513e-12
C10_188 V10 V188 -4.1215770901536614e-20

R10_189 V10 V189 -3170.4557388401163
L10_189 V10 V189 -1.4642994681020904e-11
C10_189 V10 V189 -5.595685390524258e-20

R10_190 V10 V190 -670.7431004915449
L10_190 V10 V190 2.1147812061726312e-12
C10_190 V10 V190 6.982147765268896e-20

R10_191 V10 V191 2899.275685412224
L10_191 V10 V191 -2.9619799370146678e-12
C10_191 V10 V191 -5.843851068425595e-20

R10_192 V10 V192 -1540.5757725098567
L10_192 V10 V192 -1.6126962433866165e-11
C10_192 V10 V192 -7.267439560326423e-20

R10_193 V10 V193 1475.4420291251274
L10_193 V10 V193 2.9593174940128923e-12
C10_193 V10 V193 1.539140910455273e-20

R10_194 V10 V194 2067.397012661717
L10_194 V10 V194 3.27617064151567e-11
C10_194 V10 V194 -8.425799852225446e-20

R10_195 V10 V195 -1068.8888454303706
L10_195 V10 V195 1.4363003286867883e-12
C10_195 V10 V195 9.063816170924926e-20

R10_196 V10 V196 -785.5316033500711
L10_196 V10 V196 1.0723145941848455e-12
C10_196 V10 V196 7.82678582152687e-20

R10_197 V10 V197 2860.5756221189317
L10_197 V10 V197 5.074901205370894e-12
C10_197 V10 V197 1.0059367665935767e-19

R10_198 V10 V198 1142.745921360767
L10_198 V10 V198 -2.674883189402776e-12
C10_198 V10 V198 -1.451579217720967e-20

R10_199 V10 V199 -24423.69323722894
L10_199 V10 V199 3.389105699512015e-12
C10_199 V10 V199 1.7332851776622145e-20

R10_200 V10 V200 743.7400879265518
L10_200 V10 V200 -1.4612842417556826e-11
C10_200 V10 V200 7.165971101439245e-20

R11_11 V11 0 178.3950892629741
L11_11 V11 0 8.858209253530768e-13
C11_11 V11 0 -7.703316358960585e-19

R11_12 V11 V12 -1275.480702326382
L11_12 V11 V12 -5.2709173871277954e-12
C11_12 V11 V12 -1.4701360465117082e-19

R11_13 V11 V13 2656.733225791219
L11_13 V11 V13 -1.580820971929422e-11
C11_13 V11 V13 5.622030490816419e-20

R11_14 V11 V14 3766.6057058704723
L11_14 V11 V14 1.0149369206595127e-10
C11_14 V11 V14 -6.52646344663938e-20

R11_15 V11 V15 643.4270008490296
L11_15 V11 V15 -6.680342999973925e-12
C11_15 V11 V15 8.249344803186978e-20

R11_16 V11 V16 2505.261636828839
L11_16 V11 V16 -2.0369753659086755e-11
C11_16 V11 V16 -1.1861135113603832e-20

R11_17 V11 V17 24338.545201141704
L11_17 V11 V17 4.871745423622669e-12
C11_17 V11 V17 2.804899529205743e-20

R11_18 V11 V18 -10817.551883722888
L11_18 V11 V18 8.022776849990772e-12
C11_18 V11 V18 8.517246416107089e-20

R11_19 V11 V19 809.9598214630072
L11_19 V11 V19 1.4615647799039152e-12
C11_19 V11 V19 4.2710013429782515e-19

R11_20 V11 V20 2052.023326606944
L11_20 V11 V20 3.413488465465804e-12
C11_20 V11 V20 1.8712921457689946e-19

R11_21 V11 V21 1187.1354582178826
L11_21 V11 V21 5.395956351833725e-12
C11_21 V11 V21 -7.927554718233166e-20

R11_22 V11 V22 1792.0507208605964
L11_22 V11 V22 3.981693991852263e-11
C11_22 V11 V22 -2.817782117973155e-20

R11_23 V11 V23 853.2716811847644
L11_23 V11 V23 -2.4763588681396644e-12
C11_23 V11 V23 -4.3135430076360636e-19

R11_24 V11 V24 2093.937796564266
L11_24 V11 V24 -6.986926350637858e-12
C11_24 V11 V24 -1.5324582420413876e-19

R11_25 V11 V25 -1428.1733058337184
L11_25 V11 V25 -2.891676702562753e-12
C11_25 V11 V25 -1.0504265535964198e-20

R11_26 V11 V26 -1983.752133237071
L11_26 V11 V26 -4.584179298660481e-12
C11_26 V11 V26 -5.94371936980745e-20

R11_27 V11 V27 -1498.6413665017217
L11_27 V11 V27 -6.031561344957595e-12
C11_27 V11 V27 1.4405360918330106e-19

R11_28 V11 V28 -2430.5867785589653
L11_28 V11 V28 -5.456510071915424e-12
C11_28 V11 V28 4.0450160610542106e-20

R11_29 V11 V29 -2042.8652156426938
L11_29 V11 V29 -1.757209956432271e-11
C11_29 V11 V29 8.634080687296849e-20

R11_30 V11 V30 -4614.703978081343
L11_30 V11 V30 1.600372667743578e-11
C11_30 V11 V30 6.021155294793117e-20

R11_31 V11 V31 -472.34006849578753
L11_31 V11 V31 3.1644247723972216e-12
C11_31 V11 V31 1.5786106105607973e-19

R11_32 V11 V32 -1361.0074727451074
L11_32 V11 V32 7.560882286304863e-12
C11_32 V11 V32 9.733309526470182e-20

R11_33 V11 V33 -7620.656708784151
L11_33 V11 V33 -1.4155388279848794e-11
C11_33 V11 V33 -4.492604170933088e-20

R11_34 V11 V34 6409.039329865749
L11_34 V11 V34 4.176763798111208e-11
C11_34 V11 V34 5.904564571245184e-20

R11_35 V11 V35 1347.3973651793917
L11_35 V11 V35 -3.698281577678807e-12
C11_35 V11 V35 -2.8170829237313147e-19

R11_36 V11 V36 1912.2758358168658
L11_36 V11 V36 2.514633721685349e-10
C11_36 V11 V36 -6.874839635121675e-20

R11_37 V11 V37 4125.342830763523
L11_37 V11 V37 7.301565924497515e-12
C11_37 V11 V37 -1.0291762843175418e-19

R11_38 V11 V38 10838.857522832734
L11_38 V11 V38 -9.968336932450905e-12
C11_38 V11 V38 -1.6055310900943667e-19

R11_39 V11 V39 595.0907642598455
L11_39 V11 V39 1.6256336299955153e-11
C11_39 V11 V39 1.8090892257339012e-20

R11_40 V11 V40 1011.6568956451524
L11_40 V11 V40 3.808984398613636e-11
C11_40 V11 V40 -1.1985668935990403e-20

R11_41 V11 V41 -6388.377597428726
L11_41 V11 V41 1.1582531766027219e-11
C11_41 V11 V41 6.110631168187411e-20

R11_42 V11 V42 -6672.214265907094
L11_42 V11 V42 7.631283366859669e-11
C11_42 V11 V42 -3.771133152396604e-21

R11_43 V11 V43 2725.147295756671
L11_43 V11 V43 -1.0337512848920987e-11
C11_43 V11 V43 8.256267173357405e-21

R11_44 V11 V44 -7782.23554966879
L11_44 V11 V44 1.7873331089901876e-10
C11_44 V11 V44 1.5492378959606774e-20

R11_45 V11 V45 -3106.3869960829434
L11_45 V11 V45 -6.260093880568545e-12
C11_45 V11 V45 3.0970225610993083e-20

R11_46 V11 V46 -5858.929756870442
L11_46 V11 V46 4.660445793110075e-12
C11_46 V11 V46 2.091959295440299e-19

R11_47 V11 V47 -733.7167934184239
L11_47 V11 V47 8.70656679071957e-12
C11_47 V11 V47 9.460783276212727e-20

R11_48 V11 V48 -1872.2916905137604
L11_48 V11 V48 2.7437509329858022e-11
C11_48 V11 V48 1.0876188578851064e-19

R11_49 V11 V49 -6850.502961364341
L11_49 V11 V49 -3.9598771733393203e-10
C11_49 V11 V49 3.421180175411802e-20

R11_50 V11 V50 -18691.340354720975
L11_50 V11 V50 -5.226532194847e-12
C11_50 V11 V50 -1.186851963476227e-19

R11_51 V11 V51 -1438.6773314450745
L11_51 V11 V51 1.0944779750038132e-11
C11_51 V11 V51 8.330122349167064e-20

R11_52 V11 V52 22777.050173658747
L11_52 V11 V52 -9.731197155031258e-12
C11_52 V11 V52 -7.420700504618113e-20

R11_53 V11 V53 -2807.246664679625
L11_53 V11 V53 -1.8597235251703747e-11
C11_53 V11 V53 1.6171041826643873e-21

R11_54 V11 V54 -8969.551171320549
L11_54 V11 V54 -1.455314457528736e-11
C11_54 V11 V54 -5.911878964643263e-20

R11_55 V11 V55 3303.541805517935
L11_55 V11 V55 -2.6689139982671153e-12
C11_55 V11 V55 -2.993012349292347e-19

R11_56 V11 V56 3872.675454593428
L11_56 V11 V56 -1.8960059989941643e-11
C11_56 V11 V56 -4.8039927990127745e-20

R11_57 V11 V57 10882.250835137664
L11_57 V11 V57 1.3738219006507062e-11
C11_57 V11 V57 -1.2163603671237107e-19

R11_58 V11 V58 -3578.1261985292394
L11_58 V11 V58 1.1208190256010344e-11
C11_58 V11 V58 4.9561416318167414e-20

R11_59 V11 V59 982.3672506746082
L11_59 V11 V59 8.777438343805479e-12
C11_59 V11 V59 7.879353076154148e-20

R11_60 V11 V60 1737.2641681985801
L11_60 V11 V60 6.439444873736799e-12
C11_60 V11 V60 1.0183400587352733e-19

R11_61 V11 V61 261322.04880628642
L11_61 V11 V61 -5.359423964155123e-11
C11_61 V11 V61 7.787404695251889e-20

R11_62 V11 V62 2861.447050693735
L11_62 V11 V62 -1.0799511393716321e-09
C11_62 V11 V62 -2.411188565228804e-20

R11_63 V11 V63 -19302.88769170977
L11_63 V11 V63 2.6761252940899528e-12
C11_63 V11 V63 1.992229002373136e-19

R11_64 V11 V64 -4125.61201094077
L11_64 V11 V64 4.4972647119762677e-11
C11_64 V11 V64 -4.381209440500294e-20

R11_65 V11 V65 -5035.79296885796
L11_65 V11 V65 1.2264627606791341e-11
C11_65 V11 V65 1.1197163631541865e-19

R11_66 V11 V66 -10546.048072718126
L11_66 V11 V66 1.4353543448123085e-11
C11_66 V11 V66 6.162852540024821e-20

R11_67 V11 V67 -1462.6142584973009
L11_67 V11 V67 -6.700767331835177e-12
C11_67 V11 V67 -1.4654221971603054e-19

R11_68 V11 V68 -2962.5399989840953
L11_68 V11 V68 7.835909371224243e-11
C11_68 V11 V68 -5.8599054931661044e-21

R11_69 V11 V69 -5073.145512085517
L11_69 V11 V69 -3.714205162053486e-12
C11_69 V11 V69 -9.946947338639272e-20

R11_70 V11 V70 -6874.056180479657
L11_70 V11 V70 -3.5701435157029684e-11
C11_70 V11 V70 1.2531197970897758e-20

R11_71 V11 V71 -1425.0087235335643
L11_71 V11 V71 -4.2941827349744045e-12
C11_71 V11 V71 1.8084783864414223e-20

R11_72 V11 V72 -3591.2662374966294
L11_72 V11 V72 -4.624777579129241e-11
C11_72 V11 V72 8.789370123995743e-20

R11_73 V11 V73 -2693.4968671771867
L11_73 V11 V73 -2.1484107912410054e-11
C11_73 V11 V73 -2.6911394136819024e-20

R11_74 V11 V74 7057.268467849599
L11_74 V11 V74 -7.149909016423656e-12
C11_74 V11 V74 -1.107163082196492e-19

R11_75 V11 V75 1184.534280585515
L11_75 V11 V75 6.497699580738794e-12
C11_75 V11 V75 4.254840082800138e-20

R11_76 V11 V76 1707.8816799420815
L11_76 V11 V76 -8.245580185278767e-12
C11_76 V11 V76 -8.330875435289953e-20

R11_77 V11 V77 2668.1274346744103
L11_77 V11 V77 3.766039739458369e-12
C11_77 V11 V77 2.6836961424801826e-20

R11_78 V11 V78 -4673.466453268845
L11_78 V11 V78 -3.558219435277672e-10
C11_78 V11 V78 2.4978217409264234e-20

R11_79 V11 V79 1311.7616739910266
L11_79 V11 V79 1.0256637874445069e-11
C11_79 V11 V79 6.158363974488718e-20

R11_80 V11 V80 3148.8925045187225
L11_80 V11 V80 1.9205680105528195e-11
C11_80 V11 V80 4.861523966776609e-21

R11_81 V11 V81 -2504.3883594653253
L11_81 V11 V81 -7.427925705459197e-12
C11_81 V11 V81 6.430323869277139e-20

R11_82 V11 V82 4474.669243154758
L11_82 V11 V82 6.264804824563748e-12
C11_82 V11 V82 1.2910142716377733e-19

R11_83 V11 V83 -2724.9347860982284
L11_83 V11 V83 -7.68732825258493e-12
C11_83 V11 V83 -1.2751743989460404e-19

R11_84 V11 V84 -5650.4469163630665
L11_84 V11 V84 5.275937934544472e-12
C11_84 V11 V84 8.089211910666771e-20

R11_85 V11 V85 32478.24239195398
L11_85 V11 V85 -9.979699608822956e-11
C11_85 V11 V85 1.923983479917382e-20

R11_86 V11 V86 -2976.4170460726145
L11_86 V11 V86 -1.2887100613572076e-09
C11_86 V11 V86 -3.1298698814824563e-20

R11_87 V11 V87 -1015.7704319893126
L11_87 V11 V87 3.379437088554928e-11
C11_87 V11 V87 -7.213146452963297e-20

R11_88 V11 V88 -6171.023218861609
L11_88 V11 V88 -7.05359670880707e-12
C11_88 V11 V88 -6.181469357981767e-20

R11_89 V11 V89 -3253.672642029312
L11_89 V11 V89 -5.530554651860501e-12
C11_89 V11 V89 -7.92602411937435e-20

R11_90 V11 V90 -8607.801555729311
L11_90 V11 V90 -4.5366753095296325e-12
C11_90 V11 V90 -1.9019081623681556e-19

R11_91 V11 V91 10435.548169324427
L11_91 V11 V91 1.5909785634121118e-11
C11_91 V11 V91 2.742136536251615e-19

R11_92 V11 V92 -18283.168629510743
L11_92 V11 V92 -7.122329823495982e-11
C11_92 V11 V92 1.943865932287512e-20

R11_93 V11 V93 -3074.869459427824
L11_93 V11 V93 1.5058888639519874e-11
C11_93 V11 V93 -1.2406242013309604e-20

R11_94 V11 V94 3530.0738275854105
L11_94 V11 V94 9.69098592312176e-12
C11_94 V11 V94 7.91017567541486e-20

R11_95 V11 V95 499.8831690001567
L11_95 V11 V95 1.7161294840119694e-11
C11_95 V11 V95 -1.2858014885553502e-20

R11_96 V11 V96 1349.9936076764661
L11_96 V11 V96 8.515814536053855e-12
C11_96 V11 V96 4.103873322498635e-20

R11_97 V11 V97 1769.091700613507
L11_97 V11 V97 4.486329632395633e-12
C11_97 V11 V97 9.790534213493175e-20

R11_98 V11 V98 -9610.40208884161
L11_98 V11 V98 7.631761912406481e-12
C11_98 V11 V98 1.279461286505735e-19

R11_99 V11 V99 -552.7729337217881
L11_99 V11 V99 -1.5863662604203953e-11
C11_99 V11 V99 -3.0088567337680166e-19

R11_100 V11 V100 -16579.641856482103
L11_100 V11 V100 4.599181493997328e-11
C11_100 V11 V100 -4.165935216527035e-20

R11_101 V11 V101 -3657.435937566866
L11_101 V11 V101 -6.3156500347683286e-12
C11_101 V11 V101 -3.4062260908746165e-20

R11_102 V11 V102 12032.968049181309
L11_102 V11 V102 -7.349903353245994e-12
C11_102 V11 V102 -9.815588947569644e-20

R11_103 V11 V103 48508.27570557499
L11_103 V11 V103 -1.3992507097578577e-11
C11_103 V11 V103 4.6247246391818025e-20

R11_104 V11 V104 -2627.2745919017566
L11_104 V11 V104 -8.597638335858707e-11
C11_104 V11 V104 2.0504403406279694e-21

R11_105 V11 V105 -935.5072792155978
L11_105 V11 V105 -4.808902467757188e-12
C11_105 V11 V105 -7.828695673217575e-20

R11_106 V11 V106 -1251.8408927467126
L11_106 V11 V106 -4.744178816614143e-11
C11_106 V11 V106 -1.1777654403141138e-19

R11_107 V11 V107 1479.4094793300615
L11_107 V11 V107 -1.2955897745539228e-10
C11_107 V11 V107 2.0083351454345827e-19

R11_108 V11 V108 -39690.84682357505
L11_108 V11 V108 -9.523157891032157e-12
C11_108 V11 V108 -1.1248535249065334e-20

R11_109 V11 V109 2533.9147122164936
L11_109 V11 V109 2.180290142790596e-11
C11_109 V11 V109 1.154780442917125e-19

R11_110 V11 V110 1387.4895948217834
L11_110 V11 V110 1.6145154234170952e-11
C11_110 V11 V110 1.2909093103677266e-19

R11_111 V11 V111 -484.0683558495426
L11_111 V11 V111 3.6117848533666685e-12
C11_111 V11 V111 6.292353475400728e-20

R11_112 V11 V112 -2090.489512642698
L11_112 V11 V112 1.5135939290372914e-11
C11_112 V11 V112 -2.810001433912563e-20

R11_113 V11 V113 4994.545171838048
L11_113 V11 V113 5.157650397695737e-12
C11_113 V11 V113 6.278620909893211e-20

R11_114 V11 V114 1142.6206562344914
L11_114 V11 V114 2.2430183015826753e-11
C11_114 V11 V114 8.40707721406583e-20

R11_115 V11 V115 479.3029989872937
L11_115 V11 V115 -3.022787002738254e-12
C11_115 V11 V115 -2.397147019108229e-19

R11_116 V11 V116 964.9171785524256
L11_116 V11 V116 -4.3544182690073225e-11
C11_116 V11 V116 1.9331758627020596e-20

R11_117 V11 V117 3116.4221774820335
L11_117 V11 V117 1.9071780661321512e-11
C11_117 V11 V117 -1.4393542218024478e-19

R11_118 V11 V118 -739.8515885529682
L11_118 V11 V118 -1.3023706089597066e-11
C11_118 V11 V118 -1.3540463672074937e-19

R11_119 V11 V119 -738.1300095551919
L11_119 V11 V119 -1.2824772169586652e-11
C11_119 V11 V119 1.9308811326354284e-20

R11_120 V11 V120 -1501.8540223404573
L11_120 V11 V120 -1.237249945757186e-11
C11_120 V11 V120 -4.9556523371327335e-20

R11_121 V11 V121 -2310.6725382313593
L11_121 V11 V121 -2.644376312386165e-12
C11_121 V11 V121 5.592993263255421e-20

R11_122 V11 V122 36325.63668930185
L11_122 V11 V122 6.443412313769703e-11
C11_122 V11 V122 6.150201669860955e-20

R11_123 V11 V123 -1021.2349233340876
L11_123 V11 V123 2.160430499934279e-12
C11_123 V11 V123 2.549869093577038e-19

R11_124 V11 V124 -1310.8752451810265
L11_124 V11 V124 7.402983264912698e-12
C11_124 V11 V124 2.3447615864668196e-20

R11_125 V11 V125 -623.9645567824692
L11_125 V11 V125 -7.75013286411842e-12
C11_125 V11 V125 3.954354942268655e-20

R11_126 V11 V126 2284.9007759043934
L11_126 V11 V126 9.562851053684928e-12
C11_126 V11 V126 7.290437587234942e-20

R11_127 V11 V127 524.7616306397506
L11_127 V11 V127 -7.558966842966652e-12
C11_127 V11 V127 -1.243406220747803e-19

R11_128 V11 V128 883.8295586019451
L11_128 V11 V128 3.196407523890034e-11
C11_128 V11 V128 6.752199851200093e-20

R11_129 V11 V129 602.3968940329733
L11_129 V11 V129 2.6688963835305545e-12
C11_129 V11 V129 8.888695271302609e-20

R11_130 V11 V130 1746.769727531115
L11_130 V11 V130 -1.9439703183900683e-11
C11_130 V11 V130 -9.389497393055308e-20

R11_131 V11 V131 -1033.182980727864
L11_131 V11 V131 -7.83683936792582e-12
C11_131 V11 V131 -5.482448326586661e-20

R11_132 V11 V132 -1213.474835618974
L11_132 V11 V132 -5.0245392347602925e-12
C11_132 V11 V132 -1.3601474432715364e-19

R11_133 V11 V133 1086.6086088254035
L11_133 V11 V133 -6.99785753344655e-11
C11_133 V11 V133 -1.1876934511587442e-19

R11_134 V11 V134 -4374.433609679651
L11_134 V11 V134 7.691247217500464e-11
C11_134 V11 V134 1.122806505663121e-19

R11_135 V11 V135 -1479.8846090078932
L11_135 V11 V135 3.939955358743573e-12
C11_135 V11 V135 2.1498730236062277e-19

R11_136 V11 V136 -1342.9865800783045
L11_136 V11 V136 2.119139700832515e-11
C11_136 V11 V136 -2.953672389736339e-20

R11_137 V11 V137 -526.7305784119051
L11_137 V11 V137 -7.89783628820192e-12
C11_137 V11 V137 -1.1322554305243334e-19

R11_138 V11 V138 5686.728366884047
L11_138 V11 V138 2.2938233999770673e-11
C11_138 V11 V138 -1.8252824801250982e-20

R11_139 V11 V139 1045.7736913096126
L11_139 V11 V139 -1.6347842512552155e-12
C11_139 V11 V139 -2.919548200099731e-19

R11_140 V11 V140 698.2322992247958
L11_140 V11 V140 -1.4756053721156026e-11
C11_140 V11 V140 5.445524459931494e-20

R11_141 V11 V141 -1199.8032723907377
L11_141 V11 V141 2.2018348583078107e-10
C11_141 V11 V141 2.5125331387865055e-19

R11_142 V11 V142 1634.005234826859
L11_142 V11 V142 3.7395641760433424e-11
C11_142 V11 V142 -3.256363255631117e-20

R11_143 V11 V143 -1173.1352917508402
L11_143 V11 V143 2.7143209452712696e-12
C11_143 V11 V143 1.199781028237191e-19

R11_144 V11 V144 -1770.0252569321647
L11_144 V11 V144 1.5036421839335326e-11
C11_144 V11 V144 4.0341472217804725e-20

R11_145 V11 V145 539.8840019911911
L11_145 V11 V145 1.4230198884459e-11
C11_145 V11 V145 1.3440924905737453e-19

R11_146 V11 V146 -1874.6751494057967
L11_146 V11 V146 1.3396566028808118e-11
C11_146 V11 V146 -2.3946213132272518e-20

R11_147 V11 V147 286.09821052328505
L11_147 V11 V147 3.024196358685914e-12
C11_147 V11 V147 1.5429633205553628e-19

R11_148 V11 V148 2016.4674511669605
L11_148 V11 V148 3.193237181730619e-11
C11_148 V11 V148 -2.889372382090842e-20

R11_149 V11 V149 6802.667440719739
L11_149 V11 V149 -4.678777495391461e-12
C11_149 V11 V149 -3.8977289882912516e-19

R11_150 V11 V150 -570.4194153996576
L11_150 V11 V150 -5.824767898299371e-12
C11_150 V11 V150 1.8518702085325875e-19

R11_151 V11 V151 -139.4509432805917
L11_151 V11 V151 -2.434971453601322e-12
C11_151 V11 V151 -8.750005777499884e-20

R11_152 V11 V152 -2029.6229710670414
L11_152 V11 V152 -2.9925463486412994e-10
C11_152 V11 V152 2.48781562593258e-20

R11_153 V11 V153 -1035.1606941948858
L11_153 V11 V153 -1.7879606128476926e-11
C11_153 V11 V153 -6.370973906915287e-20

R11_154 V11 V154 22562.84505009412
L11_154 V11 V154 -1.7012564581413043e-11
C11_154 V11 V154 -1.3232233975356776e-19

R11_155 V11 V155 80.86790296919494
L11_155 V11 V155 -2.671921333189058e-12
C11_155 V11 V155 -1.9107948209917184e-19

R11_156 V11 V156 -1497.6710946062906
L11_156 V11 V156 -2.8812490029794284e-11
C11_156 V11 V156 -3.064452212334982e-20

R11_157 V11 V157 -1694.1765717909177
L11_157 V11 V157 5.227914320293498e-12
C11_157 V11 V157 2.756131223243743e-19

R11_158 V11 V158 32078.842756537902
L11_158 V11 V158 6.821028350308218e-12
C11_158 V11 V158 -1.7471164865535368e-20

R11_159 V11 V159 -293.2834741434609
L11_159 V11 V159 1.457690957965312e-12
C11_159 V11 V159 7.594455427838873e-20

R11_160 V11 V160 2474.9010325278487
L11_160 V11 V160 2.771202258306984e-11
C11_160 V11 V160 -5.1933086458315125e-20

R11_161 V11 V161 2685.2566951335643
L11_161 V11 V161 -3.334564606948934e-11
C11_161 V11 V161 8.285727885037484e-20

R11_162 V11 V162 -8149.353893120372
L11_162 V11 V162 2.542811302178641e-10
C11_162 V11 V162 -8.063419187510518e-20

R11_163 V11 V163 -400.2560270218565
L11_163 V11 V163 5.579967639277041e-12
C11_163 V11 V163 -3.169302663170858e-20

R11_164 V11 V164 -783.9801577126046
L11_164 V11 V164 8.163145329069745e-12
C11_164 V11 V164 5.183719123162398e-21

R11_165 V11 V165 -1459.3283878874804
L11_165 V11 V165 -4.789369220518031e-12
C11_165 V11 V165 -1.5587976305711182e-19

R11_166 V11 V166 -2875.0004190825093
L11_166 V11 V166 -4.24455258962141e-12
C11_166 V11 V166 6.42162663235233e-20

R11_167 V11 V167 -806.269918879631
L11_167 V11 V167 -1.4108632741125644e-12
C11_167 V11 V167 4.416415173818357e-20

R11_168 V11 V168 532.9027344994362
L11_168 V11 V168 -1.2211639655173235e-11
C11_168 V11 V168 8.271065356794425e-20

R11_169 V11 V169 -1149.5988687349559
L11_169 V11 V169 6.960740126940973e-12
C11_169 V11 V169 5.464966383513231e-21

R11_170 V11 V170 -1447.300154528532
L11_170 V11 V170 9.342821755410948e-12
C11_170 V11 V170 -6.855274918725727e-20

R11_171 V11 V171 208.908402071552
L11_171 V11 V171 3.750798819882048e-11
C11_171 V11 V171 -6.942123142698887e-20

R11_172 V11 V172 5343.091812086087
L11_172 V11 V172 -2.2593243317183208e-11
C11_172 V11 V172 -4.840972081015719e-20

R11_173 V11 V173 1821.2007077834267
L11_173 V11 V173 1.1785504290672401e-11
C11_173 V11 V173 -2.083810873295013e-20

R11_174 V11 V174 584.1117213726105
L11_174 V11 V174 7.791750918055077e-12
C11_174 V11 V174 9.775041873932475e-21

R11_175 V11 V175 -377.66869794752745
L11_175 V11 V175 2.38237077257941e-12
C11_175 V11 V175 -1.5388793081245315e-19

R11_176 V11 V176 6539.267540113705
L11_176 V11 V176 5.681827489374606e-12
C11_176 V11 V176 -7.544954546515733e-20

R11_177 V11 V177 -1004.533546314938
L11_177 V11 V177 -4.0894596790694475e-11
C11_177 V11 V177 2.74295124067848e-20

R11_178 V11 V178 -991.210810113076
L11_178 V11 V178 -9.74698919188407e-11
C11_178 V11 V178 7.741902776469345e-20

R11_179 V11 V179 415.79191474988323
L11_179 V11 V179 -1.3072381286409404e-11
C11_179 V11 V179 1.9981450336208872e-19

R11_180 V11 V180 -1293.9065907083102
L11_180 V11 V180 -2.1023448173949802e-10
C11_180 V11 V180 1.2130871940140706e-19

R11_181 V11 V181 1300.3767430156938
L11_181 V11 V181 -2.7018656428645437e-11
C11_181 V11 V181 8.549851402042597e-20

R11_182 V11 V182 1139.00217016539
L11_182 V11 V182 -6.299779258984453e-12
C11_182 V11 V182 -9.724109694066591e-20

R11_183 V11 V183 -382.84408676921737
L11_183 V11 V183 1.2881785951572143e-11
C11_183 V11 V183 1.067440060571118e-20

R11_184 V11 V184 -2877.513761011533
L11_184 V11 V184 -1.2835842885993144e-10
C11_184 V11 V184 4.1222950185043634e-20

R11_185 V11 V185 -7952.542274639821
L11_185 V11 V185 -7.323421165331278e-12
C11_185 V11 V185 -7.453893790562709e-20

R11_186 V11 V186 2196.4633686373295
L11_186 V11 V186 -7.939027040970283e-12
C11_186 V11 V186 7.879071748489249e-20

R11_187 V11 V187 3825.2205733828714
L11_187 V11 V187 -7.649136120336972e-12
C11_187 V11 V187 -1.4638541722732485e-19

R11_188 V11 V188 481.4880043979528
L11_188 V11 V188 -4.450893359951062e-12
C11_188 V11 V188 -9.782889032593197e-20

R11_189 V11 V189 -1939.53842847859
L11_189 V11 V189 7.44983836143849e-12
C11_189 V11 V189 -5.2563439649109865e-20

R11_190 V11 V190 -1215.9472521108876
L11_190 V11 V190 7.669683935918103e-12
C11_190 V11 V190 6.832093933350474e-20

R11_191 V11 V191 874.8011561351746
L11_191 V11 V191 -8.002203961815923e-12
C11_191 V11 V191 2.7739655047460466e-20

R11_192 V11 V192 -2741.844754970039
L11_192 V11 V192 1.1074631766518503e-11
C11_192 V11 V192 -5.949005900907615e-20

R11_193 V11 V193 4087.29488444149
L11_193 V11 V193 6.062062130822989e-12
C11_193 V11 V193 2.796334887363933e-20

R11_194 V11 V194 2432.4486363704154
L11_194 V11 V194 5.812367273554445e-12
C11_194 V11 V194 -3.1094483392558435e-20

R11_195 V11 V195 -916.3965195889652
L11_195 V11 V195 9.951023839664663e-12
C11_195 V11 V195 -2.387279324912983e-20

R11_196 V11 V196 -377.5603311546146
L11_196 V11 V196 3.167842387340713e-12
C11_196 V11 V196 1.6789719186430482e-19

R11_197 V11 V197 -3712.2348749485855
L11_197 V11 V197 -1.1378305768631477e-11
C11_197 V11 V197 1.1571144215220953e-19

R11_198 V11 V198 -1746.9429079029576
L11_198 V11 V198 -6.896468986582821e-12
C11_198 V11 V198 -2.515936417669745e-20

R11_199 V11 V199 7647.735822278432
L11_199 V11 V199 1.9079456418829978e-11
C11_199 V11 V199 -1.7303196248884005e-21

R11_200 V11 V200 960.1048550245422
L11_200 V11 V200 -5.6418522752487874e-12
C11_200 V11 V200 2.969500805964801e-20

R12_12 V12 0 92.21775950338021
L12_12 V12 0 6.777667928277401e-13
C12_12 V12 0 -1.5189752541082696e-18

R12_13 V12 V13 2000.097624687518
L12_13 V12 V13 -1.3728407720215151e-11
C12_13 V12 V13 3.70567951470915e-20

R12_14 V12 V14 4066.1458637032893
L12_14 V12 V14 1.785782731128801e-11
C12_14 V12 V14 -8.633477273158489e-20

R12_15 V12 V15 2169.8301874413205
L12_15 V12 V15 -1.39681536108552e-10
C12_15 V12 V15 -1.1921895385350741e-19

R12_16 V12 V16 631.0827472266991
L12_16 V12 V16 -1.3648768483508558e-11
C12_16 V12 V16 1.8160677200233843e-20

R12_17 V12 V17 10063.544105699004
L12_17 V12 V17 3.933886585896053e-12
C12_17 V12 V17 6.324624890454647e-20

R12_18 V12 V18 -23142.76401743284
L12_18 V12 V18 7.613564826274169e-12
C12_18 V12 V18 1.0687989505704824e-19

R12_19 V12 V19 3257.0200578050662
L12_19 V12 V19 4.824958729754335e-12
C12_19 V12 V19 2.338797650607744e-19

R12_20 V12 V20 688.8573076036488
L12_20 V12 V20 1.3127198670647633e-12
C12_20 V12 V20 5.633739035850851e-19

R12_21 V12 V21 854.2407717850027
L12_21 V12 V21 3.932656611681915e-12
C12_21 V12 V21 -8.880925861533654e-20

R12_22 V12 V22 1657.1737445141023
L12_22 V12 V22 6.24658941705669e-11
C12_22 V12 V22 -2.935608182553925e-20

R12_23 V12 V23 2472.2609959529955
L12_23 V12 V23 -1.129116551107717e-11
C12_23 V12 V23 -1.7062843404366922e-19

R12_24 V12 V24 862.1604379478124
L12_24 V12 V24 -2.167403922273884e-12
C12_24 V12 V24 -5.093808968605689e-19

R12_25 V12 V25 -1078.6582603663137
L12_25 V12 V25 -2.3126166536173052e-12
C12_25 V12 V25 -1.7972234406552983e-20

R12_26 V12 V26 -2000.604643619087
L12_26 V12 V26 -4.09126700087874e-12
C12_26 V12 V26 -5.1797326933193567e-20

R12_27 V12 V27 -2854.172470029678
L12_27 V12 V27 -5.465277821171117e-12
C12_27 V12 V27 9.150949396350947e-20

R12_28 V12 V28 -1324.381115094358
L12_28 V12 V28 -3.2436234794763257e-12
C12_28 V12 V28 2.233372351867941e-19

R12_29 V12 V29 -1384.119955660715
L12_29 V12 V29 -8.90842435715426e-12
C12_29 V12 V29 1.169594198826423e-19

R12_30 V12 V30 -4244.852177355226
L12_30 V12 V30 1.4687472753565772e-11
C12_30 V12 V30 8.781940290677058e-20

R12_31 V12 V31 -1590.992307336645
L12_31 V12 V31 1.1376364390416995e-11
C12_31 V12 V31 3.550649402289701e-20

R12_32 V12 V32 -445.7434871197026
L12_32 V12 V32 2.746391855132273e-12
C12_32 V12 V32 1.2445922528842637e-19

R12_33 V12 V33 -7359.796806579078
L12_33 V12 V33 -2.5329914289746693e-11
C12_33 V12 V33 -5.178853193850986e-20

R12_34 V12 V34 3228.2639845770586
L12_34 V12 V34 1.6142871048864843e-11
C12_34 V12 V34 8.267361301028119e-20

R12_35 V12 V35 3723.7158259485236
L12_35 V12 V35 1.6408707944580328e-10
C12_35 V12 V35 -6.305571872348865e-20

R12_36 V12 V36 819.507346454771
L12_36 V12 V36 -6.899249661479217e-12
C12_36 V12 V36 -3.342611961302407e-19

R12_37 V12 V37 2603.945833947752
L12_37 V12 V37 5.220743946619072e-12
C12_37 V12 V37 -1.1798880862280358e-19

R12_38 V12 V38 5921.290143807158
L12_38 V12 V38 -1.1186684214299e-11
C12_38 V12 V38 -2.071155177629316e-19

R12_39 V12 V39 1537.2733548698295
L12_39 V12 V39 -3.1553219680055345e-09
C12_39 V12 V39 2.798703534728519e-20

R12_40 V12 V40 486.4315715158596
L12_40 V12 V40 2.0844624126157687e-11
C12_40 V12 V40 1.0020497374870881e-20

R12_41 V12 V41 -6132.313757617965
L12_41 V12 V41 1.2568718791860821e-11
C12_41 V12 V41 9.35229750334889e-20

R12_42 V12 V42 -8139.9498132607405
L12_42 V12 V42 3.6393288684215105e-11
C12_42 V12 V42 4.9743679973954015e-20

R12_43 V12 V43 -4682.076427683396
L12_43 V12 V43 5.0288681176048613e-11
C12_43 V12 V43 -4.900615032677405e-20

R12_44 V12 V44 4406.8073352240535
L12_44 V12 V44 -2.5164594431454864e-11
C12_44 V12 V44 7.805752754900607e-21

R12_45 V12 V45 -2106.3161345109847
L12_45 V12 V45 -4.293664496960568e-12
C12_45 V12 V45 5.129029501335999e-20

R12_46 V12 V46 -4117.007755217314
L12_46 V12 V46 5.6754183713080634e-12
C12_46 V12 V46 2.654359760421034e-19

R12_47 V12 V47 -2314.2787625725596
L12_47 V12 V47 2.994188687409992e-11
C12_47 V12 V47 9.897509088342053e-20

R12_48 V12 V48 -543.5183937789785
L12_48 V12 V48 2.5377634937641046e-11
C12_48 V12 V48 1.996607638727229e-19

R12_49 V12 V49 -5433.034323216402
L12_49 V12 V49 1.22942165934573e-10
C12_49 V12 V49 5.309157662447482e-20

R12_50 V12 V50 17038.956128682938
L12_50 V12 V50 -5.320540846274715e-12
C12_50 V12 V50 -1.310444318745386e-19

R12_51 V12 V51 -6120.073522344336
L12_51 V12 V51 -7.72980120595442e-12
C12_51 V12 V51 4.435428181821369e-21

R12_52 V12 V52 -5423.503790255776
L12_52 V12 V52 8.500443073609142e-11
C12_52 V12 V52 -6.238979485701807e-20

R12_53 V12 V53 -2685.960710795255
L12_53 V12 V53 -3.44835193790246e-11
C12_53 V12 V53 -4.3226279493810125e-21

R12_54 V12 V54 333845.9086467005
L12_54 V12 V54 -2.6531793818225134e-11
C12_54 V12 V54 -7.908444773964907e-20

R12_55 V12 V55 -9428.34567469189
L12_55 V12 V55 -4.2733632574066745e-11
C12_55 V12 V55 -4.6459599374295624e-20

R12_56 V12 V56 1093.6925142637435
L12_56 V12 V56 -2.7956922103188332e-12
C12_56 V12 V56 -3.666713518793945e-19

R12_57 V12 V57 7359.888342705846
L12_57 V12 V57 1.2164300717414277e-11
C12_57 V12 V57 -9.851735469036427e-20

R12_58 V12 V58 -3179.303216969477
L12_58 V12 V58 9.145274043618873e-12
C12_58 V12 V58 1.0332689148464492e-19

R12_59 V12 V59 2608.99984925841
L12_59 V12 V59 9.714317193206752e-12
C12_59 V12 V59 9.30643721385946e-20

R12_60 V12 V60 782.8047541096859
L12_60 V12 V60 3.962123265856295e-12
C12_60 V12 V60 1.2224693467638998e-19

R12_61 V12 V61 -38767.3763523143
L12_61 V12 V61 -1.7235992290487362e-11
C12_61 V12 V61 7.775036765877186e-20

R12_62 V12 V62 2860.6250917513776
L12_62 V12 V62 -6.424828160876903e-11
C12_62 V12 V62 1.6825549142163922e-21

R12_63 V12 V63 -7647.622874668667
L12_63 V12 V63 -1.4809528425021312e-10
C12_63 V12 V63 -1.0179580529810318e-19

R12_64 V12 V64 -2577.073866786734
L12_64 V12 V64 2.9583348220108212e-12
C12_64 V12 V64 2.321413081742345e-19

R12_65 V12 V65 -3458.7368465977215
L12_65 V12 V65 1.0970889579939584e-11
C12_65 V12 V65 1.5707108376423078e-19

R12_66 V12 V66 -406965.0993646029
L12_66 V12 V66 1.1541769951360914e-11
C12_66 V12 V66 6.389214718737035e-20

R12_67 V12 V67 156998.60788619568
L12_67 V12 V67 1.8861677979810853e-11
C12_67 V12 V67 3.330899030917398e-20

R12_68 V12 V68 -1120.9358597480655
L12_68 V12 V68 -7.540989512833646e-12
C12_68 V12 V68 -1.0239637985147143e-19

R12_69 V12 V69 -6870.192556888588
L12_69 V12 V69 -3.6942737268933315e-12
C12_69 V12 V69 -1.5703736157177662e-19

R12_70 V12 V70 -6763.206501804248
L12_70 V12 V70 -7.181753099200811e-11
C12_70 V12 V70 -2.6456426429905117e-20

R12_71 V12 V71 -7542.574373414701
L12_71 V12 V71 -4.5043417728120056e-11
C12_71 V12 V71 1.0958801529981923e-19

R12_72 V12 V72 -1377.6183908093074
L12_72 V12 V72 -4.059246680210428e-12
C12_72 V12 V72 -5.0781787823260085e-20

R12_73 V12 V73 -2963.7082318191838
L12_73 V12 V73 -1.399224747509288e-11
C12_73 V12 V73 -1.2725012460388916e-20

R12_74 V12 V74 5163.3883969638355
L12_74 V12 V74 -6.529481836653198e-12
C12_74 V12 V74 -8.030325898141845e-20

R12_75 V12 V75 -6594.839700577099
L12_75 V12 V75 -9.43435802885046e-12
C12_75 V12 V75 -8.512849162709032e-20

R12_76 V12 V76 591.2407298098587
L12_76 V12 V76 8.395211365122839e-12
C12_76 V12 V76 -4.7281832481014404e-20

R12_77 V12 V77 2886.755511953429
L12_77 V12 V77 3.279443089199408e-12
C12_77 V12 V77 6.086007258595789e-20

R12_78 V12 V78 -2488.773793744748
L12_78 V12 V78 -4.286408933672165e-11
C12_78 V12 V78 -2.5365859387016752e-20

R12_79 V12 V79 2259.648928124042
L12_79 V12 V79 9.557054964059057e-11
C12_79 V12 V79 1.8127636514539243e-20

R12_80 V12 V80 6002.697480594795
L12_80 V12 V80 6.867699965687209e-12
C12_80 V12 V80 7.89636912978686e-20

R12_81 V12 V81 -1369.6253070995622
L12_81 V12 V81 -6.029678770852325e-12
C12_81 V12 V81 9.082901012233849e-20

R12_82 V12 V82 3659.5378150432052
L12_82 V12 V82 5.752413642336562e-12
C12_82 V12 V82 1.7887082588646823e-19

R12_83 V12 V83 -6755.077935400086
L12_83 V12 V83 7.789726812188688e-12
C12_83 V12 V83 3.03883974208175e-20

R12_84 V12 V84 -2163.023958979904
L12_84 V12 V84 -1.2006362263088633e-11
C12_84 V12 V84 3.048852684189164e-20

R12_85 V12 V85 16485.182894943402
L12_85 V12 V85 -2.5497966131729635e-11
C12_85 V12 V85 2.97090310561213e-20

R12_86 V12 V86 -6731.899038944266
L12_86 V12 V86 -1.6857725908890724e-10
C12_86 V12 V86 2.898257116602002e-20

R12_87 V12 V87 -6735.144310317764
L12_87 V12 V87 -1.606582768523808e-11
C12_87 V12 V87 -1.2284636010933338e-19

R12_88 V12 V88 -1119.1228893956043
L12_88 V12 V88 -1.9489987649450497e-11
C12_88 V12 V88 -1.7000006331122173e-19

R12_89 V12 V89 -4789.295716547185
L12_89 V12 V89 -5.29121077269403e-12
C12_89 V12 V89 -1.1658087697027753e-19

R12_90 V12 V90 -7361.663457538229
L12_90 V12 V90 -4.8804197525557475e-12
C12_90 V12 V90 -2.7960296549839844e-19

R12_91 V12 V91 -2074.124779155929
L12_91 V12 V91 -2.4331988330468037e-11
C12_91 V12 V91 2.640644565356635e-19

R12_92 V12 V92 1847.5890973461342
L12_92 V12 V92 3.571024117434769e-11
C12_92 V12 V92 1.8988067588957273e-19

R12_93 V12 V93 -1866.9837264209336
L12_93 V12 V93 1.0301195930883509e-11
C12_93 V12 V93 -1.4235433749718684e-20

R12_94 V12 V94 7064.221079841094
L12_94 V12 V94 8.361167812402327e-12
C12_94 V12 V94 1.1188748208976224e-19

R12_95 V12 V95 1811.7573744858887
L12_95 V12 V95 1.065211198419358e-11
C12_95 V12 V95 2.1530112399659985e-20

R12_96 V12 V96 426.18224536002344
L12_96 V12 V96 7.724093481307503e-12
C12_96 V12 V96 5.642605964676243e-20

R12_97 V12 V97 1727.8804069980838
L12_97 V12 V97 4.374247464811745e-12
C12_97 V12 V97 2.2748592566582135e-19

R12_98 V12 V98 40806.947168130224
L12_98 V12 V98 8.452784262040092e-12
C12_98 V12 V98 2.1910568864077383e-19

R12_99 V12 V99 6401.886312815834
L12_99 V12 V99 -2.616131989176589e-11
C12_99 V12 V99 -2.996147631654696e-19

R12_100 V12 V100 -393.1167709584979
L12_100 V12 V100 7.4371241699142e-12
C12_100 V12 V100 -2.647227082308095e-19

R12_101 V12 V101 -3479.322151728601
L12_101 V12 V101 -5.7327224354483215e-12
C12_101 V12 V101 -6.068700068512257e-20

R12_102 V12 V102 8708.398126869371
L12_102 V12 V102 -7.1378386640985975e-12
C12_102 V12 V102 -1.4536796232429977e-19

R12_103 V12 V103 -2070.1079783961063
L12_103 V12 V103 -3.43428149858132e-11
C12_103 V12 V103 1.104887623627293e-19

R12_104 V12 V104 10598.889528786533
L12_104 V12 V104 -8.896939663277551e-12
C12_104 V12 V104 9.340811164531266e-20

R12_105 V12 V105 -802.9735496107965
L12_105 V12 V105 -4.915271719472223e-12
C12_105 V12 V105 -1.1376353039919665e-19

R12_106 V12 V106 -1108.1891601995767
L12_106 V12 V106 2.8596872941973643e-11
C12_106 V12 V106 -1.9062990329372718e-19

R12_107 V12 V107 -11032.331583937575
L12_107 V12 V107 3.024571510303447e-11
C12_107 V12 V107 1.6668309282786466e-19

R12_108 V12 V108 762.8666233173742
L12_108 V12 V108 -4.507748289702776e-12
C12_108 V12 V108 2.7000768079466106e-20

R12_109 V12 V109 1232.252007203751
L12_109 V12 V109 1.1364923799022141e-09
C12_109 V12 V109 1.9805572400377458e-19

R12_110 V12 V110 1046.5734447549914
L12_110 V12 V110 1.589774047837392e-10
C12_110 V12 V110 1.4285125632955031e-19

R12_111 V12 V111 -2267.31319742668
L12_111 V12 V111 3.334775335078042e-11
C12_111 V12 V111 -3.530535620300605e-20

R12_112 V12 V112 -562.8405995804634
L12_112 V12 V112 3.170069729245797e-12
C12_112 V12 V112 1.545358991550645e-19

R12_113 V12 V113 -11021.332022999157
L12_113 V12 V113 4.563793694606701e-12
C12_113 V12 V113 5.823706449632389e-20

R12_114 V12 V114 1218.575166866566
L12_114 V12 V114 3.1300979633607697e-11
C12_114 V12 V114 1.566106860708747e-19

R12_115 V12 V115 657.7991219359039
L12_115 V12 V115 -1.0903427910668886e-11
C12_115 V12 V115 -1.30238109490657e-19

R12_116 V12 V116 666.3488313877322
L12_116 V12 V116 -5.295334535626604e-12
C12_116 V12 V116 -1.434755226778113e-19

R12_117 V12 V117 4449.78041864881
L12_117 V12 V117 1.1226362857788287e-11
C12_117 V12 V117 -1.796816187470039e-19

R12_118 V12 V118 -640.8023756697677
L12_118 V12 V118 -2.4987952084282857e-11
C12_118 V12 V118 -2.1399531326374714e-19

R12_119 V12 V119 -1396.2679178863125
L12_119 V12 V119 -1.676026027703855e-11
C12_119 V12 V119 -6.729650507794933e-20

R12_120 V12 V120 -540.2834632944011
L12_120 V12 V120 -4.783947347977133e-12
C12_120 V12 V120 -1.811211732509692e-19

R12_121 V12 V121 -8261.12114406875
L12_121 V12 V121 -2.237094237466939e-12
C12_121 V12 V121 9.48846102870864e-20

R12_122 V12 V122 4089.492169630031
L12_122 V12 V122 -5.912936414020551e-11
C12_122 V12 V122 2.527348443527765e-20

R12_123 V12 V123 -1229.0879741576318
L12_123 V12 V123 7.114995063401861e-12
C12_123 V12 V123 1.710698488753649e-19

R12_124 V12 V124 4532.2562532314705
L12_124 V12 V124 1.9248001434754616e-12
C12_124 V12 V124 4.263263432689288e-19

R12_125 V12 V125 -561.1120060599254
L12_125 V12 V125 -5.813393601980622e-12
C12_125 V12 V125 4.0804647998021914e-20

R12_126 V12 V126 2340.949037125724
L12_126 V12 V126 1.217328170143899e-11
C12_126 V12 V126 1.2567810270570483e-19

R12_127 V12 V127 734.7891700324966
L12_127 V12 V127 3.2885492985272584e-11
C12_127 V12 V127 1.2177114218315904e-20

R12_128 V12 V128 504.7771235905029
L12_128 V12 V128 -2.733183662735107e-11
C12_128 V12 V128 -4.39478936305363e-20

R12_129 V12 V129 556.8536714770208
L12_129 V12 V129 2.425943040239206e-12
C12_129 V12 V129 1.0718449238526044e-19

R12_130 V12 V130 2240.996145662986
L12_130 V12 V130 2.9533177248765e-10
C12_130 V12 V130 -1.3845160126904998e-19

R12_131 V12 V131 -772.4712112164542
L12_131 V12 V131 -8.482230826336343e-12
C12_131 V12 V131 -1.0843139366146944e-19

R12_132 V12 V132 -483.78098223416345
L12_132 V12 V132 -4.591777099221129e-12
C12_132 V12 V132 -2.553745087577654e-19

R12_133 V12 V133 1543.1164996076238
L12_133 V12 V133 3.038586263952842e-11
C12_133 V12 V133 -1.796303503320659e-19

R12_134 V12 V134 -1614.852281735145
L12_134 V12 V134 -2.977893068270176e-11
C12_134 V12 V134 1.92284143722703e-21

R12_135 V12 V135 -56923.27685025052
L12_135 V12 V135 1.8566228774231587e-11
C12_135 V12 V135 8.794241609838125e-20

R12_136 V12 V136 -1512.048955781769
L12_136 V12 V136 4.842724838262411e-12
C12_136 V12 V136 2.4904154385150155e-19

R12_137 V12 V137 -597.3718588085355
L12_137 V12 V137 -1.1118842703657494e-11
C12_137 V12 V137 -7.317691279893633e-20

R12_138 V12 V138 1813.7604373892084
L12_138 V12 V138 2.3928152714055015e-11
C12_138 V12 V138 6.970831116659188e-20

R12_139 V12 V139 595.1293262719341
L12_139 V12 V139 -9.329116771668784e-12
C12_139 V12 V139 -1.705899936141856e-19

R12_140 V12 V140 2763.0366404716815
L12_140 V12 V140 -2.152660434860205e-12
C12_140 V12 V140 -2.5536967225093123e-19

R12_141 V12 V141 -1953.559651949821
L12_141 V12 V141 -1.028978295660385e-11
C12_141 V12 V141 2.797573732144768e-19

R12_142 V12 V142 969.6458482714354
L12_142 V12 V142 1.4590340891480997e-11
C12_142 V12 V142 -1.0654512299130024e-20

R12_143 V12 V143 -839.2572590109424
L12_143 V12 V143 5.0300329349438384e-12
C12_143 V12 V143 1.0149088631145353e-19

R12_144 V12 V144 328.4171696170674
L12_144 V12 V144 4.028855440825725e-12
C12_144 V12 V144 6.958766161765106e-20

R12_145 V12 V145 651.9470006551372
L12_145 V12 V145 6.425673767149553e-11
C12_145 V12 V145 1.081443312312724e-19

R12_146 V12 V146 -2150.3298007504472
L12_146 V12 V146 1.642807598395906e-11
C12_146 V12 V146 -6.66803491222982e-20

R12_147 V12 V147 880.2808980038302
L12_147 V12 V147 1.7823713104522772e-11
C12_147 V12 V147 1.572679628294746e-19

R12_148 V12 V148 -184.70622855341347
L12_148 V12 V148 4.720915510870285e-12
C12_148 V12 V148 1.4885440686176033e-19

R12_149 V12 V149 2797.3132260568473
L12_149 V12 V149 -1.565141253816507e-11
C12_149 V12 V149 -3.7485267381414307e-19

R12_150 V12 V150 -474.8319388086282
L12_150 V12 V150 -5.019192673190721e-12
C12_150 V12 V150 2.344902175557474e-19

R12_151 V12 V151 -1092.732154974455
L12_151 V12 V151 -4.422403552485687e-12
C12_151 V12 V151 -7.321061138350204e-20

R12_152 V12 V152 773.2996217477449
L12_152 V12 V152 -3.695547185712781e-12
C12_152 V12 V152 -2.354217238353702e-20

R12_153 V12 V153 -1718.86134600121
L12_153 V12 V153 -1.001300553892785e-11
C12_153 V12 V153 -7.307938191587121e-20

R12_154 V12 V154 663.980294807331
L12_154 V12 V154 -9.458786158806437e-12
C12_154 V12 V154 -1.1869574359215884e-19

R12_155 V12 V155 354.89234515386124
L12_155 V12 V155 -7.330952144316092e-12
C12_155 V12 V155 -1.7126408437718778e-19

R12_156 V12 V156 -617.400296022463
L12_156 V12 V156 -4.579474788555645e-12
C12_156 V12 V156 -1.50553240580113e-19

R12_157 V12 V157 -631.7992933324979
L12_157 V12 V157 7.615808161271886e-12
C12_157 V12 V157 3.6523348586756204e-19

R12_158 V12 V158 -937.0731890556303
L12_158 V12 V158 4.361493291553192e-12
C12_158 V12 V158 -1.819370802301791e-20

R12_159 V12 V159 -346.15497219057323
L12_159 V12 V159 6.988105620735822e-12
C12_159 V12 V159 6.648729251255038e-20

R12_160 V12 V160 244.57892508953339
L12_160 V12 V160 1.655382253871404e-12
C12_160 V12 V160 9.599697444906978e-21

R12_161 V12 V161 1143.543484775953
L12_161 V12 V161 -1.527775044109829e-11
C12_161 V12 V161 4.076440238457331e-20

R12_162 V12 V162 -36088.5042584647
L12_162 V12 V162 2.0270260320035865e-11
C12_162 V12 V162 -7.487764402333652e-20

R12_163 V12 V163 -11004.417609561295
L12_163 V12 V163 5.641894708979727e-12
C12_163 V12 V163 1.216657089368192e-20

R12_164 V12 V164 -168.97121333358942
L12_164 V12 V164 7.198513736397416e-12
C12_164 V12 V164 -3.6427799080974266e-20

R12_165 V12 V165 -556.410658890846
L12_165 V12 V165 -4.627740363207858e-12
C12_165 V12 V165 -1.2137783816896646e-19

R12_166 V12 V166 -1413.5403918012858
L12_166 V12 V166 -3.1599589995971497e-12
C12_166 V12 V166 1.1647647846227182e-19

R12_167 V12 V167 -718.2123137069483
L12_167 V12 V167 -1.2410068858897129e-11
C12_167 V12 V167 2.6268433969865115e-20

R12_168 V12 V168 223.3027530367643
L12_168 V12 V168 -1.2887800205588884e-12
C12_168 V12 V168 5.868780444377641e-20

R12_169 V12 V169 -2150.412664440419
L12_169 V12 V169 6.590941606231604e-12
C12_169 V12 V169 9.180871888004644e-20

R12_170 V12 V170 -3171.669187441406
L12_170 V12 V170 1.518661995768618e-11
C12_170 V12 V170 -7.100367419537235e-20

R12_171 V12 V171 749.5194064245898
L12_171 V12 V171 -4.917036116579832e-12
C12_171 V12 V171 -4.791240853992527e-20

R12_172 V12 V172 1014.1193691998631
L12_172 V12 V172 5.871328098911924e-12
C12_172 V12 V172 -5.458204539461373e-20

R12_173 V12 V173 1866.589227021092
L12_173 V12 V173 1.0337523542449887e-11
C12_173 V12 V173 -7.80780421822035e-20

R12_174 V12 V174 543.0403687762565
L12_174 V12 V174 4.309196501863251e-12
C12_174 V12 V174 1.5267483038195998e-20

R12_175 V12 V175 -69651.25076956824
L12_175 V12 V175 5.848399092266901e-12
C12_175 V12 V175 -1.502871582073616e-19

R12_176 V12 V176 -438.11079471102596
L12_176 V12 V176 2.2900755872468344e-12
C12_176 V12 V176 -1.637966558037483e-19

R12_177 V12 V177 -877.6858137593383
L12_177 V12 V177 -3.1152383250074745e-11
C12_177 V12 V177 5.130558490909609e-20

R12_178 V12 V178 -857.1021465334458
L12_178 V12 V178 -3.198606043959364e-11
C12_178 V12 V178 6.764789294194006e-20

R12_179 V12 V179 1373682.0923077094
L12_179 V12 V179 9.545205940089252e-12
C12_179 V12 V179 1.868056139817504e-19

R12_180 V12 V180 2426.916589092923
L12_180 V12 V180 -4.743174236569745e-12
C12_180 V12 V180 2.0526917556196873e-19

R12_181 V12 V181 1093.5466155478282
L12_181 V12 V181 -4.771172288778553e-11
C12_181 V12 V181 8.316611876162115e-20

R12_182 V12 V182 965.0292387594774
L12_182 V12 V182 -6.727899667790833e-12
C12_182 V12 V182 -8.827417349738965e-20

R12_183 V12 V183 -1303.4365179993442
L12_183 V12 V183 2.7978491827828122e-11
C12_183 V12 V183 3.674389867882771e-20

R12_184 V12 V184 -1276.2669825648397
L12_184 V12 V184 -3.167390960591564e-11
C12_184 V12 V184 6.1133296677529776e-21

R12_185 V12 V185 -2780.9894231357293
L12_185 V12 V185 -5.5312657349131365e-12
C12_185 V12 V185 -8.397830174393013e-20

R12_186 V12 V186 29230.82858726173
L12_186 V12 V186 -7.693638447614624e-12
C12_186 V12 V186 6.995014891505631e-20

R12_187 V12 V187 2029.6552251004257
L12_187 V12 V187 -4.601338974006203e-12
C12_187 V12 V187 -1.6137784167917218e-19

R12_188 V12 V188 351.18371064138904
L12_188 V12 V188 -6.373697837379219e-12
C12_188 V12 V188 -1.525498689530782e-19

R12_189 V12 V189 -16275.572183476539
L12_189 V12 V189 6.564847048829609e-12
C12_189 V12 V189 -2.961501318601808e-20

R12_190 V12 V190 -992.0546921240851
L12_190 V12 V190 7.441316737181508e-12
C12_190 V12 V190 9.392547665052468e-20

R12_191 V12 V191 1630.756796624638
L12_191 V12 V191 -7.0775838773506e-12
C12_191 V12 V191 7.98959204363301e-21

R12_192 V12 V192 -5220.780866876636
L12_192 V12 V192 4.018517710737863e-12
C12_192 V12 V192 6.642283236141113e-20

R12_193 V12 V193 1290.9666024282344
L12_193 V12 V193 4.15279327226922e-12
C12_193 V12 V193 3.358972094269476e-20

R12_194 V12 V194 12858.705940711117
L12_194 V12 V194 3.5845521629741334e-12
C12_194 V12 V194 6.138455377807258e-20

R12_195 V12 V195 -829.0429165008829
L12_195 V12 V195 3.2933971231170797e-12
C12_195 V12 V195 1.055309208954255e-19

R12_196 V12 V196 -398.41123160207167
L12_196 V12 V196 1.434862676114468e-11
C12_196 V12 V196 -4.1260179892757523e-20

R12_197 V12 V197 11506.943733646294
L12_197 V12 V197 -6.755915922858174e-12
C12_197 V12 V197 7.490482243298513e-20

R12_198 V12 V198 -1152.8600972949023
L12_198 V12 V198 -6.500446505473268e-12
C12_198 V12 V198 2.9895806187149324e-20

R12_199 V12 V199 -385.45859838172055
L12_199 V12 V199 4.586029542258455e-11
C12_199 V12 V199 4.8386868279685496e-20

R12_200 V12 V200 326.4583256731352
L12_200 V12 V200 -9.420645402223638e-12
C12_200 V12 V200 -2.1569645539136135e-20

R13_13 V13 0 -126.00385989689562
L13_13 V13 0 3.0482400088464765e-13
C13_13 V13 0 3.9383492496306183e-19

R13_14 V13 V14 -6780.416052450479
L13_14 V13 V14 -3.134709541976162e-12
C13_14 V13 V14 -2.839326447330141e-19

R13_15 V13 V15 -12022.486694005944
L13_15 V13 V15 -3.042379028858527e-12
C13_15 V13 V15 -2.460075820905288e-19

R13_16 V13 V16 -7346.796401485821
L13_16 V13 V16 -2.3137089570990345e-12
C13_16 V13 V16 -2.895770296405162e-19

R13_17 V13 V17 -3011.2523130939935
L13_17 V13 V17 5.009110549693235e-12
C13_17 V13 V17 3.088568956995593e-19

R13_18 V13 V18 11716.37104195479
L13_18 V13 V18 -3.789965172908577e-11
C13_18 V13 V18 9.74092945339988e-20

R13_19 V13 V19 -29561.608342075517
L13_19 V13 V19 -1.433794421012195e-10
C13_19 V13 V19 8.112431690279547e-20

R13_20 V13 V20 -14958.262013415713
L13_20 V13 V20 -4.452993805033883e-11
C13_20 V13 V20 1.1064918394184378e-19

R13_21 V13 V21 -359.99750665982714
L13_21 V13 V21 1.0681544549446716e-12
C13_21 V13 V21 2.0394115482278144e-19

R13_22 V13 V22 -1657.1583025558589
L13_22 V13 V22 4.875832125013876e-12
C13_22 V13 V22 4.8030666715415087e-20

R13_23 V13 V23 -2780.1612393774717
L13_23 V13 V23 6.807490397726985e-12
C13_23 V13 V23 4.803733963648493e-20

R13_24 V13 V24 -2026.4124519853353
L13_24 V13 V24 5.4236351308178865e-12
C13_24 V13 V24 7.209454217200691e-20

R13_25 V13 V25 487.4146911153406
L13_25 V13 V25 -1.917467069899801e-12
C13_25 V13 V25 -3.3072029311280966e-19

R13_26 V13 V26 2950.337447577797
L13_26 V13 V26 -3.055630004043532e-11
C13_26 V13 V26 -1.5524562356090967e-20

R13_27 V13 V27 6601.930381848594
L13_27 V13 V27 -4.086709956587255e-11
C13_27 V13 V27 -5.869597193486824e-20

R13_28 V13 V28 4004.3351320115075
L13_28 V13 V28 -2.8625553798122453e-11
C13_28 V13 V28 -1.093320473171663e-19

R13_29 V13 V29 432.53163928872436
L13_29 V13 V29 -3.194096336439338e-12
C13_29 V13 V29 -1.327475601495674e-20

R13_30 V13 V30 5648.210376248685
L13_30 V13 V30 -2.4802687450278462e-11
C13_30 V13 V30 -4.232664007488101e-20

R13_31 V13 V31 6104.780620911593
L13_31 V13 V31 -3.9589115749817914e-11
C13_31 V13 V31 -3.260881995924e-20

R13_32 V13 V32 3966.532609328343
L13_32 V13 V32 -4.857206020719313e-11
C13_32 V13 V32 -7.591090495181866e-20

R13_33 V13 V33 1417.9136517271963
L13_33 V13 V33 -1.4509737246478524e-12
C13_33 V13 V33 -1.465491316943614e-19

R13_34 V13 V34 -14260.393803541076
L13_34 V13 V34 -4.876663420307575e-12
C13_34 V13 V34 -5.266776968960244e-20

R13_35 V13 V35 -4722.624787163759
L13_35 V13 V35 -8.337784361960327e-12
C13_35 V13 V35 -4.310756617014498e-20

R13_36 V13 V36 -2882.1492638017126
L13_36 V13 V36 -6.156086871859577e-12
C13_36 V13 V36 -1.2375223764101673e-19

R13_37 V13 V37 -1243.0772162289502
L13_37 V13 V37 2.344558220165781e-12
C13_37 V13 V37 4.186035137000437e-19

R13_38 V13 V38 -7936.759753724742
L13_38 V13 V38 8.244245743772312e-11
C13_38 V13 V38 8.542616947326816e-20

R13_39 V13 V39 -7121.070237091603
L13_39 V13 V39 1.2026745869961204e-11
C13_39 V13 V39 1.2876498605622395e-19

R13_40 V13 V40 -4502.3322991335035
L13_40 V13 V40 7.832250887306913e-12
C13_40 V13 V40 1.8044884239572273e-19

R13_41 V13 V41 -3102.8462225859585
L13_41 V13 V41 1.0898092659956589e-11
C13_41 V13 V41 2.6535822064161876e-21

R13_42 V13 V42 -5800.666433961604
L13_42 V13 V42 7.920206877795165e-12
C13_42 V13 V42 5.565539827839546e-20

R13_43 V13 V43 -3893.657020493182
L13_43 V13 V43 1.1043910951784982e-11
C13_43 V13 V43 1.2085435158776526e-20

R13_44 V13 V44 -3007.4581594178007
L13_44 V13 V44 7.314020403650692e-12
C13_44 V13 V44 -2.132465883389119e-20

R13_45 V13 V45 776.3586993387174
L13_45 V13 V45 -1.2607575522181094e-11
C13_45 V13 V45 -2.1288210342894827e-19

R13_46 V13 V46 25348.30722618353
L13_46 V13 V46 4.411614044365082e-12
C13_46 V13 V46 1.1447502770166302e-19

R13_47 V13 V47 -52742.57233893063
L13_47 V13 V47 1.4538280341306424e-11
C13_47 V13 V47 -4.945295540144957e-21

R13_48 V13 V48 10490.329431211187
L13_48 V13 V48 9.312447328862292e-12
C13_48 V13 V48 -1.532412837048176e-20

R13_49 V13 V49 794.871918547179
L13_49 V13 V49 -3.0771740176613184e-12
C13_49 V13 V49 -7.886967000081961e-20

R13_50 V13 V50 -8890.971218223478
L13_50 V13 V50 -4.468101192055956e-12
C13_50 V13 V50 -1.6686681249243924e-19

R13_51 V13 V51 -14797.635329101106
L13_51 V13 V51 -5.393631108532629e-12
C13_51 V13 V51 -1.4714317901848287e-19

R13_52 V13 V52 -5080.486530527386
L13_52 V13 V52 -4.210686360062411e-12
C13_52 V13 V52 -2.1261133107387481e-19

R13_53 V13 V53 1800.4987495252833
L13_53 V13 V53 -1.509723231607951e-11
C13_53 V13 V53 8.27998839051095e-20

R13_54 V13 V54 5758.877184835049
L13_54 V13 V54 -5.68890505373678e-12
C13_54 V13 V54 -7.031578858208533e-20

R13_55 V13 V55 4554.500376379942
L13_55 V13 V55 -1.3590715806305473e-11
C13_55 V13 V55 -1.5823362427983672e-20

R13_56 V13 V56 7500.395914160168
L13_56 V13 V56 -6.440001027342591e-12
C13_56 V13 V56 -6.326192475900285e-20

R13_57 V13 V57 -26580.735346266556
L13_57 V13 V57 6.120397462871687e-12
C13_57 V13 V57 4.506972804913158e-19

R13_58 V13 V58 -3987.4145809345428
L13_58 V13 V58 3.6109096737574845e-12
C13_58 V13 V58 2.1404441395110775e-19

R13_59 V13 V59 -2855.3938593935127
L13_59 V13 V59 3.397598648732434e-12
C13_59 V13 V59 2.3770040934756595e-19

R13_60 V13 V60 -1960.8061110816282
L13_60 V13 V60 2.3890244096500316e-12
C13_60 V13 V60 3.0012564654795557e-19

R13_61 V13 V61 -3389.7554321176885
L13_61 V13 V61 -5.056986077595889e-12
C13_61 V13 V61 -3.3949408876164495e-19

R13_62 V13 V62 43792.92934141948
L13_62 V13 V62 6.2354610595596306e-12
C13_62 V13 V62 1.2962551353299804e-19

R13_63 V13 V63 -150465.68877906335
L13_63 V13 V63 9.878819213807728e-12
C13_63 V13 V63 8.029238175396392e-20

R13_64 V13 V64 15994.93530563629
L13_64 V13 V64 7.074762515050474e-12
C13_64 V13 V64 6.252266050200351e-20

R13_65 V13 V65 1029.3957801336692
L13_65 V13 V65 -3.306459369589559e-12
C13_65 V13 V65 -2.1576922179638364e-19

R13_66 V13 V66 -8977.578231503363
L13_66 V13 V66 -3.676120657320538e-12
C13_66 V13 V66 -1.7537536916536724e-19

R13_67 V13 V67 -8714.805596941093
L13_67 V13 V67 -2.9327285373074064e-12
C13_67 V13 V67 -2.756079282667049e-19

R13_68 V13 V68 -12169.042031622854
L13_68 V13 V68 -2.523537117483182e-12
C13_68 V13 V68 -3.8719892838803893e-19

R13_69 V13 V69 1789.943757067364
L13_69 V13 V69 5.09550426371734e-11
C13_69 V13 V69 -7.249268196404887e-21

R13_70 V13 V70 -9854.5416997829
L13_70 V13 V70 1.1019905281996563e-10
C13_70 V13 V70 -6.496717132299532e-20

R13_71 V13 V71 -15371.839498092362
L13_71 V13 V71 6.67195370973076e-11
C13_71 V13 V71 -2.4389140626856882e-20

R13_72 V13 V72 -11849.23319554469
L13_72 V13 V72 -2.0183966454104708e-11
C13_72 V13 V72 -3.6614197019859167e-20

R13_73 V13 V73 4608.744260666085
L13_73 V13 V73 4.8654859617532375e-12
C13_73 V13 V73 3.7000582988698046e-19

R13_74 V13 V74 6759.090477692668
L13_74 V13 V74 3.003694267973736e-12
C13_74 V13 V74 2.775451358654618e-19

R13_75 V13 V75 6958.967964377572
L13_75 V13 V75 2.7950995712989135e-12
C13_75 V13 V75 2.6357328583649473e-19

R13_76 V13 V76 63466.46261113189
L13_76 V13 V76 2.799721563057745e-12
C13_76 V13 V76 2.7736210874300556e-19

R13_77 V13 V77 -4274.017774611052
L13_77 V13 V77 -6.799229338798971e-12
C13_77 V13 V77 1.0022743635296612e-19

R13_78 V13 V78 9654.519188231248
L13_78 V13 V78 -5.29804861995984e-12
C13_78 V13 V78 -1.3296072453996337e-19

R13_79 V13 V79 -32882.97119124974
L13_79 V13 V79 -4.7920460355062654e-12
C13_79 V13 V79 -6.749076264458506e-20

R13_80 V13 V80 -43549.3504117318
L13_80 V13 V80 -5.064167235110812e-12
C13_80 V13 V80 -7.743557645615062e-20

R13_81 V13 V81 539.3928017277613
L13_81 V13 V81 -3.2738100912439978e-12
C13_81 V13 V81 -3.18275291797857e-19

R13_82 V13 V82 -3738.2687622188246
L13_82 V13 V82 -6.115647093280522e-12
C13_82 V13 V82 -6.09966905688894e-20

R13_83 V13 V83 -2100.927912593019
L13_83 V13 V83 -8.427389093335237e-12
C13_83 V13 V83 -6.575666982665329e-20

R13_84 V13 V84 -2269.4774798298363
L13_84 V13 V84 -1.1042363538679654e-11
C13_84 V13 V84 -1.2875058094820816e-19

R13_85 V13 V85 -18978.792582616195
L13_85 V13 V85 4.708826557228907e-12
C13_85 V13 V85 4.013070708004874e-20

R13_86 V13 V86 -1418.1495182176184
L13_86 V13 V86 4.589512066027558e-12
C13_86 V13 V86 8.982672054946058e-20

R13_87 V13 V87 -4965.752956619174
L13_87 V13 V87 5.827176400596386e-12
C13_87 V13 V87 -8.677872628418044e-21

R13_88 V13 V88 -3777.7548785270687
L13_88 V13 V88 8.459765331889387e-12
C13_88 V13 V88 -6.01926815962754e-20

R13_89 V13 V89 13827.330156945689
L13_89 V13 V89 -3.330575927570578e-12
C13_89 V13 V89 -1.6187746429751732e-19

R13_90 V13 V90 1989.01595551951
L13_90 V13 V90 8.777801917099245e-12
C13_90 V13 V90 -8.617408857036354e-21

R13_91 V13 V91 2845.062626142881
L13_91 V13 V91 6.054831113073674e-12
C13_91 V13 V91 2.6809419509448768e-20

R13_92 V13 V92 5885.91883318582
L13_92 V13 V92 4.782068859111873e-12
C13_92 V13 V92 1.0570807015590003e-19

R13_93 V13 V93 908.7305626518315
L13_93 V13 V93 -1.881629622472122e-11
C13_93 V13 V93 1.6293793782577087e-19

R13_94 V13 V94 2824.690182538131
L13_94 V13 V94 -4.888780657791745e-12
C13_94 V13 V94 -1.7685401428581483e-20

R13_95 V13 V95 7819.876921101599
L13_95 V13 V95 -6.098529107837624e-12
C13_95 V13 V95 3.473022626838241e-20

R13_96 V13 V96 3950.58760646074
L13_96 V13 V96 -4.871509627005712e-12
C13_96 V13 V96 4.50396451454749e-20

R13_97 V13 V97 1426.7733873079137
L13_97 V13 V97 1.4705217173635907e-11
C13_97 V13 V97 4.146855173931642e-19

R13_98 V13 V98 -1005.3670203806406
L13_98 V13 V98 9.496591526374298e-12
C13_98 V13 V98 3.965430192450086e-20

R13_99 V13 V99 -962.1365771250443
L13_99 V13 V99 -9.329947547204844e-12
C13_99 V13 V99 -6.780097839845156e-20

R13_100 V13 V100 -912.4690417753735
L13_100 V13 V100 -6.000054068182254e-11
C13_100 V13 V100 -1.4823821574315187e-19

R13_101 V13 V101 -1971.9821444808374
L13_101 V13 V101 -6.260473200830085e-12
C13_101 V13 V101 -3.7654345808687724e-19

R13_102 V13 V102 -24726.918089665043
L13_102 V13 V102 9.914385552270134e-12
C13_102 V13 V102 5.960568033548422e-20

R13_103 V13 V103 19239.985088035708
L13_103 V13 V103 4.334206651362322e-12
C13_103 V13 V103 1.0470412969674761e-19

R13_104 V13 V104 -11254.75576150082
L13_104 V13 V104 3.5736226378009715e-12
C13_104 V13 V104 1.1415233465205013e-19

R13_105 V13 V105 421.49683105519676
L13_105 V13 V105 -3.828249663538614e-12
C13_105 V13 V105 -1.3915898904420096e-19

R13_106 V13 V106 -4696.180679888889
L13_106 V13 V106 -2.061067988452139e-11
C13_106 V13 V106 -1.2460524718806167e-19

R13_107 V13 V107 9160.945025039995
L13_107 V13 V107 3.213454888674687e-11
C13_107 V13 V107 -1.8992719427857287e-20

R13_108 V13 V108 4414.0363058560615
L13_108 V13 V108 -7.90755195355836e-12
C13_108 V13 V108 -7.681970183527815e-20

R13_109 V13 V109 -2042.0917249080555
L13_109 V13 V109 7.426971317249474e-12
C13_109 V13 V109 1.5622872889090993e-19

R13_110 V13 V110 9135.921064453425
L13_110 V13 V110 -6.570623691099224e-11
C13_110 V13 V110 3.541579183174214e-21

R13_111 V13 V111 -9302.313613850207
L13_111 V13 V111 -1.3570696672416318e-11
C13_111 V13 V111 -1.3448030344282628e-19

R13_112 V13 V112 -5326.591862977784
L13_112 V13 V112 8.706477688319555e-11
C13_112 V13 V112 5.624158139656193e-21

R13_113 V13 V113 5201.174120282204
L13_113 V13 V113 -7.137387474697716e-12
C13_113 V13 V113 1.1838390339739484e-19

R13_114 V13 V114 -10763.575264221021
L13_114 V13 V114 1.0525610815557008e-11
C13_114 V13 V114 1.5490010647469877e-19

R13_115 V13 V115 -6958.383907517659
L13_115 V13 V115 -3.685723336891857e-10
C13_115 V13 V115 1.2457532558916837e-19

R13_116 V13 V116 -14417.398684274878
L13_116 V13 V116 -5.5585716654680705e-11
C13_116 V13 V116 1.1553376655050264e-19

R13_117 V13 V117 846.6477218170145
L13_117 V13 V117 2.7854239495729878e-11
C13_117 V13 V117 2.277513116228876e-19

R13_118 V13 V118 -18819.892770419814
L13_118 V13 V118 -4.802995706123287e-11
C13_118 V13 V118 -1.5129768915556435e-19

R13_119 V13 V119 -3789.712028483909
L13_119 V13 V119 -7.650238149931904e-09
C13_119 V13 V119 -8.561603019295848e-20

R13_120 V13 V120 -2312.711937463982
L13_120 V13 V120 5.712817962100933e-11
C13_120 V13 V120 -1.182926102031245e-19

R13_121 V13 V121 -3388.6888700568093
L13_121 V13 V121 -2.610568862357003e-12
C13_121 V13 V121 -4.56671880532664e-19

R13_122 V13 V122 -3471.3759230437704
L13_122 V13 V122 -1.3427530601256124e-11
C13_122 V13 V122 -1.0922512283112495e-20

R13_123 V13 V123 6853.163517211708
L13_123 V13 V123 2.0543927258724272e-10
C13_123 V13 V123 6.074273637691785e-20

R13_124 V13 V124 3978.892931837478
L13_124 V13 V124 1.9417887509177127e-11
C13_124 V13 V124 7.652780825011327e-20

R13_125 V13 V125 746.1198188458682
L13_125 V13 V125 -1.2005248468718249e-11
C13_125 V13 V125 -1.7783201974809703e-19

R13_126 V13 V126 -98870.81707518714
L13_126 V13 V126 1.4409218021290645e-11
C13_126 V13 V126 -2.909963264226976e-20

R13_127 V13 V127 13415.656073521253
L13_127 V13 V127 3.0839073200694303e-11
C13_127 V13 V127 -5.693156344301303e-22

R13_128 V13 V128 3237.322608720086
L13_128 V13 V128 -2.4105225540896515e-11
C13_128 V13 V128 -3.804961164570408e-20

R13_129 V13 V129 230380.11046950248
L13_129 V13 V129 1.0440022516401297e-11
C13_129 V13 V129 3.3746665203178027e-19

R13_130 V13 V130 5640.36154654018
L13_130 V13 V130 2.444251106465312e-11
C13_130 V13 V130 4.808157283091902e-20

R13_131 V13 V131 -8174.174137762083
L13_131 V13 V131 -7.488757043818054e-10
C13_131 V13 V131 -3.020502947124316e-20

R13_132 V13 V132 -1672.2642793385664
L13_132 V13 V132 1.5972096542337487e-10
C13_132 V13 V132 -9.959037894762138e-21

R13_133 V13 V133 -1164.2398483602603
L13_133 V13 V133 3.665556433421377e-12
C13_133 V13 V133 1.9032211442239583e-19

R13_134 V13 V134 -1451.6194455971872
L13_134 V13 V134 8.959114124844567e-12
C13_134 V13 V134 5.2189488322660115e-20

R13_135 V13 V135 12554.843452796285
L13_135 V13 V135 9.291376136615683e-12
C13_135 V13 V135 6.722228458950332e-20

R13_136 V13 V136 3886.257630664953
L13_136 V13 V136 6.709077029466034e-12
C13_136 V13 V136 1.8452712081925715e-19

R13_137 V13 V137 766.6875083149381
L13_137 V13 V137 -3.2885602341632776e-11
C13_137 V13 V137 -5.856400061724121e-20

R13_138 V13 V138 1114.3317465913972
L13_138 V13 V138 -9.87901697739732e-12
C13_138 V13 V138 -7.565414550672578e-20

R13_139 V13 V139 -3419.795865637325
L13_139 V13 V139 -4.855393776685174e-12
C13_139 V13 V139 -1.428093930433876e-19

R13_140 V13 V140 -3832.73278655865
L13_140 V13 V140 -3.7398477797332995e-12
C13_140 V13 V140 -2.0275981445642244e-19

R13_141 V13 V141 -1129.4792615459269
L13_141 V13 V141 -7.7137041964197e-12
C13_141 V13 V141 -2.20326404336469e-19

R13_142 V13 V142 -1897.60277328407
L13_142 V13 V142 -2.1300029740239666e-11
C13_142 V13 V142 -2.7308660527203096e-20

R13_143 V13 V143 -5708.815148488161
L13_143 V13 V143 6.91574211666831e-12
C13_143 V13 V143 1.3723559055694921e-19

R13_144 V13 V144 -2485.549190191442
L13_144 V13 V144 1.1942780568965473e-11
C13_144 V13 V144 -3.901094558603696e-21

R13_145 V13 V145 629.7020239772484
L13_145 V13 V145 -6.852537024707354e-12
C13_145 V13 V145 -2.879319961867981e-20

R13_146 V13 V146 -1867.931740355695
L13_146 V13 V146 1.1883650906341211e-11
C13_146 V13 V146 7.094022423511038e-20

R13_147 V13 V147 3383.3080711717575
L13_147 V13 V147 9.830548013921401e-12
C13_147 V13 V147 -3.391802942687532e-20

R13_148 V13 V148 1465.425127440471
L13_148 V13 V148 5.345076527209096e-12
C13_148 V13 V148 2.825341962459575e-20

R13_149 V13 V149 -415.33310636630046
L13_149 V13 V149 -2.2908278508268036e-12
C13_149 V13 V149 -6.802681070927951e-20

R13_150 V13 V150 1365.6175680395954
L13_150 V13 V150 7.74590768692359e-12
C13_150 V13 V150 4.8301029754651127e-20

R13_151 V13 V151 2466.413602011815
L13_151 V13 V151 -1.1150192296189854e-11
C13_151 V13 V151 -9.243607410506707e-20

R13_152 V13 V152 -2522.6674799212396
L13_152 V13 V152 -1.598371373726784e-11
C13_152 V13 V152 2.3671149882019946e-20

R13_153 V13 V153 568.8795901004055
L13_153 V13 V153 3.286990244511646e-12
C13_153 V13 V153 1.9879895099585764e-19

R13_154 V13 V154 -5524.196261913944
L13_154 V13 V154 -1.675438269359721e-11
C13_154 V13 V154 4.919320856093019e-22

R13_155 V13 V155 -1076.6749261392372
L13_155 V13 V155 -9.593721389869967e-12
C13_155 V13 V155 -5.81963921223696e-20

R13_156 V13 V156 -26809.421212943904
L13_156 V13 V156 -2.106792779781095e-11
C13_156 V13 V156 -2.0320061121289253e-20

R13_157 V13 V157 659.2980673984508
L13_157 V13 V157 2.3112559726128606e-12
C13_157 V13 V157 4.1854436103107097e-19

R13_158 V13 V158 -3519.032474292358
L13_158 V13 V158 -4.014648654365631e-11
C13_158 V13 V158 -7.028550848191724e-20

R13_159 V13 V159 6805.089353303527
L13_159 V13 V159 1.1714671768719701e-11
C13_159 V13 V159 1.151772152029984e-19

R13_160 V13 V160 -4247.004997230091
L13_160 V13 V160 1.4408711072727384e-11
C13_160 V13 V160 2.430213918763968e-20

R13_161 V13 V161 1845.0613000760004
L13_161 V13 V161 -2.376528187052533e-12
C13_161 V13 V161 -4.286364205199313e-19

R13_162 V13 V162 -9723.017031728446
L13_162 V13 V162 2.2577679343305353e-10
C13_162 V13 V162 1.3111893947221617e-19

R13_163 V13 V163 -1524.6825158137708
L13_163 V13 V163 7.156794118324901e-12
C13_163 V13 V163 1.3540927871323623e-19

R13_164 V13 V164 -3779.1311575097197
L13_164 V13 V164 1.6656973311425207e-11
C13_164 V13 V164 -9.174665280593119e-21

R13_165 V13 V165 968.4928137195352
L13_165 V13 V165 -2.48112138684374e-12
C13_165 V13 V165 -2.0322257463087205e-19

R13_166 V13 V166 -1263.5868356561607
L13_166 V13 V166 3.349365211843901e-11
C13_166 V13 V166 -5.2857091526987586e-20

R13_167 V13 V167 -44733.88352726278
L13_167 V13 V167 -1.0821491223915511e-11
C13_167 V13 V167 -1.7712097755385995e-19

R13_168 V13 V168 -1308.6510971843968
L13_168 V13 V168 -8.06698297636588e-12
C13_168 V13 V168 -1.7939915389498101e-19

R13_169 V13 V169 -8618.466585895807
L13_169 V13 V169 -1.7364347046809937e-10
C13_169 V13 V169 1.4992946902843584e-19

R13_170 V13 V170 689.7228506282132
L13_170 V13 V170 -4.153952382713714e-12
C13_170 V13 V170 -1.4029990165171804e-19

R13_171 V13 V171 931.4168628407798
L13_171 V13 V171 -3.6110249739683597e-12
C13_171 V13 V171 -1.4347206001632436e-19

R13_172 V13 V172 1143.9235116837692
L13_172 V13 V172 -7.047300783883886e-12
C13_172 V13 V172 -1.3038460564201365e-20

R13_173 V13 V173 674.7573985028176
L13_173 V13 V173 3.536162507074634e-12
C13_173 V13 V173 3.613529047901385e-19

R13_174 V13 V174 -1200.7084219288304
L13_174 V13 V174 6.746730555907457e-12
C13_174 V13 V174 2.9661335349547525e-19

R13_175 V13 V175 -901.0052970704435
L13_175 V13 V175 3.0064586135410202e-12
C13_175 V13 V175 2.2571133361894355e-19

R13_176 V13 V176 -1149.6353775415648
L13_176 V13 V176 2.6447868300021456e-12
C13_176 V13 V176 2.590507791517425e-19

R13_177 V13 V177 -1347.5512830163973
L13_177 V13 V177 -4.3730512891290354e-12
C13_177 V13 V177 -1.8153130499308701e-19

R13_178 V13 V178 35643.011373033325
L13_178 V13 V178 3.842598410834813e-12
C13_178 V13 V178 2.2907197737218143e-20

R13_179 V13 V179 21066.68594148763
L13_179 V13 V179 8.796039869133547e-12
C13_179 V13 V179 7.865190548950261e-20

R13_180 V13 V180 3629.877194787324
L13_180 V13 V180 1.0932506054363966e-11
C13_180 V13 V180 -6.047376883462023e-21

R13_181 V13 V181 -1214.3021785643487
L13_181 V13 V181 -4.747316169114023e-12
C13_181 V13 V181 -3.78236554424513e-19

R13_182 V13 V182 1887.5694161785325
L13_182 V13 V182 -5.553794762058575e-12
C13_182 V13 V182 -1.072757904065128e-19

R13_183 V13 V183 2427.1078331371173
L13_183 V13 V183 -5.878180198299924e-12
C13_183 V13 V183 -4.178059048216989e-20

R13_184 V13 V184 2597.5166512422466
L13_184 V13 V184 -3.6075697497955475e-12
C13_184 V13 V184 -1.0934360328417415e-19

R13_185 V13 V185 370.0902967546091
L13_185 V13 V185 2.3685080726934073e-12
C13_185 V13 V185 3.201694127646232e-19

R13_186 V13 V186 -873.9067538244286
L13_186 V13 V186 -2.2611118305517415e-12
C13_186 V13 V186 -2.3134892157619726e-19

R13_187 V13 V187 -2828.5929913554323
L13_187 V13 V187 -5.872178516880992e-12
C13_187 V13 V187 -1.591232935400232e-19

R13_188 V13 V188 -3654.6640834618206
L13_188 V13 V188 -4.445521530232524e-12
C13_188 V13 V188 -1.4711875633704442e-19

R13_189 V13 V189 -345.6735734565041
L13_189 V13 V189 9.174091507462425e-12
C13_189 V13 V189 3.916273490230288e-20

R13_190 V13 V190 4669.6953306901
L13_190 V13 V190 4.064320007857161e-12
C13_190 V13 V190 1.390464083688648e-19

R13_191 V13 V191 1195.2931358709554
L13_191 V13 V191 3.722676744977321e-12
C13_191 V13 V191 5.0610442729714193e-20

R13_192 V13 V192 1625.1353265155992
L13_192 V13 V192 1.863627047086957e-12
C13_192 V13 V192 2.4590469901316876e-19

R13_193 V13 V193 37385.56799891134
L13_193 V13 V193 -2.504450846425713e-12
C13_193 V13 V193 1.43767588401534e-19

R13_194 V13 V194 969.9841224019669
L13_194 V13 V194 2.4583777747901265e-12
C13_194 V13 V194 2.284999316549016e-19

R13_195 V13 V195 -15834.230788936897
L13_195 V13 V195 2.0714103805585976e-11
C13_195 V13 V195 5.2203050233520107e-20

R13_196 V13 V196 -14555.709617831904
L13_196 V13 V196 1.6011359500285553e-11
C13_196 V13 V196 1.2905644371269706e-20

R13_197 V13 V197 619.0743783956336
L13_197 V13 V197 3.318728774091407e-11
C13_197 V13 V197 -2.712029304663626e-19

R13_198 V13 V198 -1231.6888040231272
L13_198 V13 V198 -3.277142979082369e-12
C13_198 V13 V198 -2.47557350673271e-20

R13_199 V13 V199 -828.7223519623586
L13_199 V13 V199 -2.993066523078131e-12
C13_199 V13 V199 1.2654958832315251e-19

R13_200 V13 V200 -1010.5640088436639
L13_200 V13 V200 -1.8617617726702783e-12
C13_200 V13 V200 -1.7739889573186443e-19

R14_14 V14 0 -196.141262028668
L14_14 V14 0 1.0855794415151526e-12
C14_14 V14 0 -1.1212805638438888e-18

R14_15 V14 V15 -4344.728492265129
L14_15 V14 V15 -1.4383273058084853e-12
C14_15 V14 V15 -4.490433740547944e-19

R14_16 V14 V16 -4449.44516652368
L14_16 V14 V16 -1.0757241000114447e-12
C14_16 V14 V16 -5.69096579129594e-19

R14_17 V14 V17 14924.996201235255
L14_17 V14 V17 1.11976155120817e-10
C14_17 V14 V17 9.226845246972861e-20

R14_18 V14 V18 -3082.3151976365143
L14_18 V14 V18 5.12299892965732e-11
C14_18 V14 V18 2.1196591940898842e-19

R14_19 V14 V19 -9739.444665028865
L14_19 V14 V19 -2.1300885031314583e-11
C14_19 V14 V19 7.160665503457923e-20

R14_20 V14 V20 -7093.594224531532
L14_20 V14 V20 -8.670853977761804e-12
C14_20 V14 V20 8.232328372751126e-20

R14_21 V14 V21 -4216.850708157822
L14_21 V14 V21 -2.0491277493753946e-11
C14_21 V14 V21 -4.631713669990203e-20

R14_22 V14 V22 -1091.6583175096293
L14_22 V14 V22 7.549685604069579e-13
C14_22 V14 V22 5.957418374379075e-19

R14_23 V14 V23 -4654.881094723086
L14_23 V14 V23 7.902779458584564e-12
C14_23 V14 V23 1.139785033359647e-19

R14_24 V14 V24 -4267.224363696228
L14_24 V14 V24 8.11478048130724e-12
C14_24 V14 V24 1.298538683451395e-19

R14_25 V14 V25 4624.280115060827
L14_25 V14 V25 1.9609939559464956e-11
C14_25 V14 V25 8.674055781393473e-21

R14_26 V14 V26 1656.812634100172
L14_26 V14 V26 -1.2992130831360684e-12
C14_26 V14 V26 -4.424807722691862e-19

R14_27 V14 V27 5526.948919698097
L14_27 V14 V27 2.4503219186970454e-11
C14_27 V14 V27 -4.203431001699051e-20

R14_28 V14 V28 4402.293782938281
L14_28 V14 V28 4.960966540966531e-12
C14_28 V14 V28 2.0399736756174395e-20

R14_29 V14 V29 7879.561145752887
L14_29 V14 V29 2.92345238749887e-12
C14_29 V14 V29 2.3110217789916056e-19

R14_30 V14 V30 889.9828822849587
L14_30 V14 V30 -1.5210982172250671e-12
C14_30 V14 V30 -1.9045831872358205e-19

R14_31 V14 V31 3180.5234885965724
L14_31 V14 V31 6.293322415954013e-11
C14_31 V14 V31 -1.9693584856479073e-20

R14_32 V14 V32 3037.99344408105
L14_32 V14 V32 1.3264098324652723e-11
C14_32 V14 V32 -4.878063545942954e-20

R14_33 V14 V33 -24042.108714151225
L14_33 V14 V33 -1.3027226973532006e-12
C14_33 V14 V33 -3.452194595372391e-19

R14_34 V14 V34 -2181.158812928357
L14_34 V14 V34 8.284695716110865e-12
C14_34 V14 V34 3.633086495610207e-19

R14_35 V14 V35 -4424.295832476534
L14_35 V14 V35 -4.5356044993238884e-12
C14_35 V14 V35 -1.0030220782863473e-19

R14_36 V14 V36 -2617.0223830933423
L14_36 V14 V36 -3.4579296600117145e-12
C14_36 V14 V36 -1.9814345793368738e-19

R14_37 V14 V37 -30256.82875060155
L14_37 V14 V37 -5.028609640390374e-12
C14_37 V14 V37 -3.6563608516640785e-20

R14_38 V14 V38 -2670.0098777143016
L14_38 V14 V38 4.264479305684053e-12
C14_38 V14 V38 3.7832199328388074e-20

R14_39 V14 V39 -3988.0734195182445
L14_39 V14 V39 -6.469042350964752e-11
C14_39 V14 V39 2.0818658318794473e-20

R14_40 V14 V40 -2927.1524277609988
L14_40 V14 V40 8.703550629151959e-11
C14_40 V14 V40 5.531042500840376e-20

R14_41 V14 V41 7274.282761522254
L14_41 V14 V41 2.5409215216744925e-12
C14_41 V14 V41 2.887254902335151e-19

R14_42 V14 V42 -2206.541576257557
L14_42 V14 V42 -3.071647224085304e-12
C14_42 V14 V42 -1.3832782595522564e-19

R14_43 V14 V43 -34088.21491420261
L14_43 V14 V43 8.584425971517593e-12
C14_43 V14 V43 7.040668091181265e-20

R14_44 V14 V44 -399242.1396372106
L14_44 V14 V44 4.838524605469443e-12
C14_44 V14 V44 8.061164445438942e-20

R14_45 V14 V45 6076.328355922947
L14_45 V14 V45 4.025473514644346e-12
C14_45 V14 V45 9.250339636964721e-20

R14_46 V14 V46 1233.8136503522107
L14_46 V14 V46 1.0034199282988514e-11
C14_46 V14 V46 5.291980729261529e-20

R14_47 V14 V47 5470.8849630961395
L14_47 V14 V47 4.4885866761644405e-12
C14_47 V14 V47 1.1291630307680777e-19

R14_48 V14 V48 3262.7411487322674
L14_48 V14 V48 2.9329931779442963e-12
C14_48 V14 V48 1.6683129685839674e-19

R14_49 V14 V49 -30800.41673705945
L14_49 V14 V49 -3.0107784214030634e-12
C14_49 V14 V49 -1.525958710531492e-19

R14_50 V14 V50 2125.6122362086
L14_50 V14 V50 -4.439609092162392e-12
C14_50 V14 V50 -8.733742144116015e-20

R14_51 V14 V51 22356.25990019196
L14_51 V14 V51 -3.429290835165667e-12
C14_51 V14 V51 -2.31702042611596e-19

R14_52 V14 V52 -11403.015347494504
L14_52 V14 V52 -2.8869014411509605e-12
C14_52 V14 V52 -3.152250700858164e-19

R14_53 V14 V53 11124.082132711706
L14_53 V14 V53 -2.420635703356565e-12
C14_53 V14 V53 -1.973181217135386e-19

R14_54 V14 V54 -2201.226544244983
L14_54 V14 V54 2.9911429364762967e-12
C14_54 V14 V54 2.360113369141511e-19

R14_55 V14 V55 -9752.017333232841
L14_55 V14 V55 -1.1413486296372941e-11
C14_55 V14 V55 -3.969270695240839e-20

R14_56 V14 V56 -3047.803395890529
L14_56 V14 V56 -4.506073954613361e-12
C14_56 V14 V56 -1.4855641470760697e-19

R14_57 V14 V57 87458.56790103884
L14_57 V14 V57 4.135790487445106e-12
C14_57 V14 V57 3.076197101091832e-19

R14_58 V14 V58 4296.869078056024
L14_58 V14 V58 -2.2196351949184733e-12
C14_58 V14 V58 -1.843154740796595e-19

R14_59 V14 V59 -19763.65204003686
L14_59 V14 V59 2.6317248689854005e-12
C14_59 V14 V59 2.621369343239834e-19

R14_60 V14 V60 -10784.682597454888
L14_60 V14 V60 2.0309992026649947e-12
C14_60 V14 V60 3.1541985338708666e-19

R14_61 V14 V61 17381.66448521804
L14_61 V14 V61 4.672864600016989e-12
C14_61 V14 V61 2.701051011322814e-20

R14_62 V14 V62 -2366.9756660029416
L14_62 V14 V62 -3.764468562518669e-12
C14_62 V14 V62 -8.433052853672006e-20

R14_63 V14 V63 26585.6624260071
L14_63 V14 V63 -1.2130059864792794e-11
C14_63 V14 V63 -5.986188034797166e-20

R14_64 V14 V64 5941.057941879974
L14_64 V14 V64 1.906782937199666e-09
C14_64 V14 V64 -5.1223708422981875e-20

R14_65 V14 V65 10563.183265867237
L14_65 V14 V65 -4.038625773514789e-12
C14_65 V14 V65 -9.932641385744342e-20

R14_66 V14 V66 1865.8262061704904
L14_66 V14 V66 1.8368338916389187e-12
C14_66 V14 V66 3.9526911376201627e-19

R14_67 V14 V67 -227627.39641042557
L14_67 V14 V67 -4.188632278496158e-12
C14_67 V14 V67 -1.541705694842226e-19

R14_68 V14 V68 10770.06357561867
L14_68 V14 V68 -6.7171854889682446e-12
C14_68 V14 V68 -1.3178548224965944e-19

R14_69 V14 V69 -6646.019553736471
L14_69 V14 V69 -8.927150837293827e-12
C14_69 V14 V69 -1.238284289199688e-19

R14_70 V14 V70 2353.570864231869
L14_70 V14 V70 -2.875573982417293e-12
C14_70 V14 V70 -4.004123199169466e-19

R14_71 V14 V71 8787.834773604938
L14_71 V14 V71 3.926283968906882e-12
C14_71 V14 V71 1.306562961089742e-19

R14_72 V14 V72 11611.955822425905
L14_72 V14 V72 5.431797805202678e-12
C14_72 V14 V72 9.640765688931593e-20

R14_73 V14 V73 2852.9100850671393
L14_73 V14 V73 1.1124797455896465e-11
C14_73 V14 V73 1.5480385078426724e-19

R14_74 V14 V74 -1529.372627970845
L14_74 V14 V74 -2.0317140827784114e-12
C14_74 V14 V74 -9.920666701930177e-20

R14_75 V14 V75 20002.592487977094
L14_75 V14 V75 1.1372021751594004e-11
C14_75 V14 V75 5.916082787858332e-20

R14_76 V14 V76 -3702.3834525039288
L14_76 V14 V76 -7.834730051893005e-12
C14_76 V14 V76 -1.0220681359789782e-19

R14_77 V14 V77 -12351.986385618537
L14_77 V14 V77 -1.2109311163602684e-10
C14_77 V14 V77 1.2634472420807168e-19

R14_78 V14 V78 6187.478588362647
L14_78 V14 V78 1.8859219145590965e-12
C14_78 V14 V78 2.577202723980056e-19

R14_79 V14 V79 -3960.6414866896494
L14_79 V14 V79 -6.591784725074625e-12
C14_79 V14 V79 -6.8730822427373e-20

R14_80 V14 V80 -11738.990857641907
L14_80 V14 V80 2.0947121038004724e-11
C14_80 V14 V80 5.535516703092321e-20

R14_81 V14 V81 5036.7660205471475
L14_81 V14 V81 -1.5241460523610772e-11
C14_81 V14 V81 -6.339746986879841e-20

R14_82 V14 V82 4201.606708484987
L14_82 V14 V82 1.3889113977293657e-11
C14_82 V14 V82 1.4413352169410634e-19

R14_83 V14 V83 20631.403468312295
L14_83 V14 V83 -8.153837585096511e-11
C14_83 V14 V83 1.7967578442837923e-20

R14_84 V14 V84 6004.202007724739
L14_84 V14 V84 4.642594023027778e-12
C14_84 V14 V84 1.0629383395537143e-19

R14_85 V14 V85 -9192.733189650906
L14_85 V14 V85 9.362837362833625e-12
C14_85 V14 V85 3.205204075922479e-21

R14_86 V14 V86 1286.7967907989653
L14_86 V14 V86 -8.015895839167032e-12
C14_86 V14 V86 -1.1788525288128847e-19

R14_87 V14 V87 26675.74024705264
L14_87 V14 V87 2.5437952128281924e-11
C14_87 V14 V87 -6.265477746925608e-20

R14_88 V14 V88 -26245.33971435619
L14_88 V14 V88 -8.409048325072623e-12
C14_88 V14 V88 -1.7576794685544103e-19

R14_89 V14 V89 -127074.50632460625
L14_89 V14 V89 -5.143399868075868e-12
C14_89 V14 V89 -1.247557292534543e-19

R14_90 V14 V90 -1035.423786124328
L14_90 V14 V90 -2.47209947657149e-12
C14_90 V14 V90 -2.9867047068199876e-19

R14_91 V14 V91 15040.905062826647
L14_91 V14 V91 3.2022145121976583e-12
C14_91 V14 V91 1.3012973291831517e-19

R14_92 V14 V92 -17131.819293120767
L14_92 V14 V92 3.7442764004190944e-12
C14_92 V14 V92 7.80749537764633e-20

R14_93 V14 V93 5337.265313207377
L14_93 V14 V93 -1.1340970019389466e-11
C14_93 V14 V93 5.896640454338125e-20

R14_94 V14 V94 -3260.171416240934
L14_94 V14 V94 3.129083004437783e-12
C14_94 V14 V94 2.66770960023692e-19

R14_95 V14 V95 -30469.839495780718
L14_95 V14 V95 -1.4477822417679406e-10
C14_95 V14 V95 9.457370906056423e-20

R14_96 V14 V96 -12052.385271691894
L14_96 V14 V96 -3.2977116892148937e-11
C14_96 V14 V96 1.442948812037368e-19

R14_97 V14 V97 -3987.3064048223005
L14_97 V14 V97 5.380054117810751e-12
C14_97 V14 V97 3.1943351212900155e-19

R14_98 V14 V98 1034.9983420986014
L14_98 V14 V98 -8.179609087971657e-12
C14_98 V14 V98 2.5398466841727934e-20

R14_99 V14 V99 -1994.1008849789225
L14_99 V14 V99 -3.0572604422805664e-12
C14_99 V14 V99 -2.5248428228013276e-19

R14_100 V14 V100 -2835.880611155097
L14_100 V14 V100 -3.621184648488756e-11
C14_100 V14 V100 -2.0094373943460401e-19

R14_101 V14 V101 4488.217153585745
L14_101 V14 V101 -4.887814249988068e-12
C14_101 V14 V101 -1.953758498462208e-19

R14_102 V14 V102 -1422.9658019628005
L14_102 V14 V102 1.145100985495847e-11
C14_102 V14 V102 2.7167080096216565e-20

R14_103 V14 V103 2983.531553621835
L14_103 V14 V103 -4.7205867348240113e-11
C14_103 V14 V103 -5.61568616881648e-20

R14_104 V14 V104 2444.189140657277
L14_104 V14 V104 5.485713713828055e-11
C14_104 V14 V104 -2.9696572229657935e-20

R14_105 V14 V105 4351.364741482113
L14_105 V14 V105 -3.0730600481577665e-12
C14_105 V14 V105 -1.9621980745975637e-19

R14_106 V14 V106 663.6670251503458
L14_106 V14 V106 -1.5546308112114172e-11
C14_106 V14 V106 -1.4955651036536438e-19

R14_107 V14 V107 4419.067199133647
L14_107 V14 V107 2.720229327226342e-12
C14_107 V14 V107 2.8372947223580324e-19

R14_108 V14 V108 26202.817058254823
L14_108 V14 V108 -1.1791379113643365e-10
C14_108 V14 V108 9.202717315584485e-20

R14_109 V14 V109 -2142.253777659074
L14_109 V14 V109 3.620270256239962e-12
C14_109 V14 V109 2.3082050690836667e-19

R14_110 V14 V110 -843.1890063184474
L14_110 V14 V110 -1.7467609347275883e-12
C14_110 V14 V110 -2.054000784482998e-19

R14_111 V14 V111 13266.399605202621
L14_111 V14 V111 8.006856683479366e-12
C14_111 V14 V111 8.116055424635545e-22

R14_112 V14 V112 -20634.478985510024
L14_112 V14 V112 6.009493640286589e-12
C14_112 V14 V112 6.775265237647533e-20

R14_113 V14 V113 2965.972185478238
L14_113 V14 V113 7.05812970980787e-12
C14_113 V14 V113 2.0060075134536454e-19

R14_114 V14 V114 -932.3110410331496
L14_114 V14 V114 2.6122331045351904e-12
C14_114 V14 V114 4.370989741559781e-19

R14_115 V14 V115 -1696.4801182918497
L14_115 V14 V115 -2.1163253908783788e-12
C14_115 V14 V115 -2.0486053285549348e-19

R14_116 V14 V116 -2912.686050973034
L14_116 V14 V116 -3.827486902416068e-12
C14_116 V14 V116 -5.65295769075985e-20

R14_117 V14 V117 -36649.19938879565
L14_117 V14 V117 -2.337563264268074e-12
C14_117 V14 V117 -1.239267269589716e-19

R14_118 V14 V118 473.8745516230454
L14_118 V14 V118 4.362805714895148e-12
C14_118 V14 V118 -1.4439033543665957e-19

R14_119 V14 V119 2392.990141684653
L14_119 V14 V119 1.049618963713158e-11
C14_119 V14 V119 -3.1580332507798926e-20

R14_120 V14 V120 3538.5169066084054
L14_120 V14 V120 -3.037406990235591e-11
C14_120 V14 V120 -1.47060078889044e-19

R14_121 V14 V121 -9893.552991942275
L14_121 V14 V121 -4.321867910267188e-12
C14_121 V14 V121 -2.1031163574222168e-19

R14_122 V14 V122 -92495.24761942994
L14_122 V14 V122 -8.446709958437119e-12
C14_122 V14 V122 -6.191129556580154e-20

R14_123 V14 V123 2126.932949225721
L14_123 V14 V123 4.885321202559318e-12
C14_123 V14 V123 1.3044459758440741e-19

R14_124 V14 V124 2080.4514096713633
L14_124 V14 V124 3.4995602386685754e-12
C14_124 V14 V124 2.2181677757029633e-19

R14_125 V14 V125 1907.4123810062592
L14_125 V14 V125 2.6748536901397843e-12
C14_125 V14 V125 4.739212278750542e-20

R14_126 V14 V126 -846.1324980960774
L14_126 V14 V126 -3.573136772326497e-12
C14_126 V14 V126 3.103830816116328e-20

R14_127 V14 V127 -1148.6952454105872
L14_127 V14 V127 -8.581728010306312e-12
C14_127 V14 V127 8.827270713675866e-20

R14_128 V14 V128 -1287.2042556549175
L14_128 V14 V128 -5.56178442208522e-12
C14_128 V14 V128 6.911833835351703e-20

R14_129 V14 V129 -2418.377052021783
L14_129 V14 V129 6.77524227739442e-12
C14_129 V14 V129 3.878493078951952e-19

R14_130 V14 V130 -85128.80298930242
L14_130 V14 V130 -6.245088433105778e-12
C14_130 V14 V130 -1.2110283829493804e-19

R14_131 V14 V131 1445.5977215738997
L14_131 V14 V131 2.2843463784388738e-11
C14_131 V14 V131 -1.3528548626870572e-19

R14_132 V14 V132 1366.165960464924
L14_132 V14 V132 -1.4971840650486766e-11
C14_132 V14 V132 -2.699485562909832e-19

R14_133 V14 V133 -2672.5374406589
L14_133 V14 V133 -1.7430570810877397e-12
C14_133 V14 V133 -2.9178095185561966e-19

R14_134 V14 V134 721.1630141706431
L14_134 V14 V134 1.1963417804228632e-12
C14_134 V14 V134 3.272997903482548e-19

R14_135 V14 V135 2131.746024694151
L14_135 V14 V135 3.171451976823514e-11
C14_135 V14 V135 -5.135281027179932e-20

R14_136 V14 V136 1200.262393480391
L14_136 V14 V136 3.5565662757105356e-12
C14_136 V14 V136 1.5753904234882741e-19

R14_137 V14 V137 931.4887399024584
L14_137 V14 V137 1.3571038930130301e-11
C14_137 V14 V137 -1.988629595273439e-19

R14_138 V14 V138 -1204.4236470330188
L14_138 V14 V138 -1.8583232032058285e-12
C14_138 V14 V138 -2.176809300845197e-19

R14_139 V14 V139 -887.900575980008
L14_139 V14 V139 -3.3552363715668984e-12
C14_139 V14 V139 -2.3478914527121427e-20

R14_140 V14 V140 -789.9521121245839
L14_140 V14 V140 -2.1768240523042383e-12
C14_140 V14 V140 -1.0813585980695375e-19

R14_141 V14 V141 6661.014836137286
L14_141 V14 V141 1.3764251640753908e-12
C14_141 V14 V141 4.61111153105103e-19

R14_142 V14 V142 -466.69417476447455
L14_142 V14 V142 -8.641417427145292e-13
C14_142 V14 V142 -1.2213872964497073e-19

R14_143 V14 V143 1571.4957763674213
L14_143 V14 V143 3.947977577403018e-12
C14_143 V14 V143 1.9066003359801306e-19

R14_144 V14 V144 -5846.540163454101
L14_144 V14 V144 2.4997376274224427e-11
C14_144 V14 V144 5.623237275414849e-20

R14_145 V14 V145 -1021.1985084053114
L14_145 V14 V145 -2.3147114434209386e-12
C14_145 V14 V145 1.2960984082430056e-19

R14_146 V14 V146 307.82651695607154
L14_146 V14 V146 8.880116602209555e-13
C14_146 V14 V146 1.3588167278611793e-19

R14_147 V14 V147 -3061.3317061055436
L14_147 V14 V147 9.405524232411286e-12
C14_147 V14 V147 -1.6930104115578153e-20

R14_148 V14 V148 666.1883560356418
L14_148 V14 V148 3.195201290872939e-12
C14_148 V14 V148 7.201926059021951e-20

R14_149 V14 V149 9147.713817424055
L14_149 V14 V149 -9.97391236714176e-13
C14_149 V14 V149 -7.771037689509118e-19

R14_150 V14 V150 991.0743831947788
L14_150 V14 V150 1.037992590992713e-12
C14_150 V14 V150 4.43163519918921e-19

R14_151 V14 V151 19822.31909791141
L14_151 V14 V151 -3.3319517684919275e-12
C14_151 V14 V151 -1.191630722824123e-19

R14_152 V14 V152 -472.3756929435962
L14_152 V14 V152 -3.709914634969576e-12
C14_152 V14 V152 1.4141863849991347e-20

R14_153 V14 V153 1132.4223574744387
L14_153 V14 V153 2.581330616589322e-12
C14_153 V14 V153 3.991322238131445e-20

R14_154 V14 V154 -596.7691526223426
L14_154 V14 V154 -1.9132538688121873e-12
C14_154 V14 V154 -3.860797377967552e-19

R14_155 V14 V155 -639.0829904466483
L14_155 V14 V155 -4.9475118807449354e-12
C14_155 V14 V155 -1.4140789842623158e-19

R14_156 V14 V156 425.7352366733596
L14_156 V14 V156 1.3762097210517994e-11
C14_156 V14 V156 -1.3029460740357805e-19

R14_157 V14 V157 -7756.745891958435
L14_157 V14 V157 1.1344770215472414e-12
C14_157 V14 V157 8.102931565426078e-19

R14_158 V14 V158 -5593.40077386748
L14_158 V14 V158 -8.255370878091543e-13
C14_158 V14 V158 -2.2511886253212643e-21

R14_159 V14 V159 417.2687515499585
L14_159 V14 V159 2.5842824646300117e-12
C14_159 V14 V159 2.5487202372713706e-20

R14_160 V14 V160 2073.915324441487
L14_160 V14 V160 3.6166444428220437e-12
C14_160 V14 V160 -4.5785707863625096e-20

R14_161 V14 V161 -1109.4390971763376
L14_161 V14 V161 -3.283992392438341e-12
C14_161 V14 V161 -6.903663886105892e-20

R14_162 V14 V162 1035.8353911171635
L14_162 V14 V162 6.3377082188844294e-12
C14_162 V14 V162 4.872505109336026e-20

R14_163 V14 V163 -1063.7419041156725
L14_163 V14 V163 2.3437335829026248e-11
C14_163 V14 V163 1.8163792937385648e-19

R14_164 V14 V164 -1365.7465220790834
L14_164 V14 V164 -5.2131343037530974e-12
C14_164 V14 V164 6.614037024055252e-21

R14_165 V14 V165 861.9370853012421
L14_165 V14 V165 -1.7012631507276396e-12
C14_165 V14 V165 -4.628875033093877e-19

R14_166 V14 V166 823.7565488171313
L14_166 V14 V166 7.497112884472689e-13
C14_166 V14 V166 5.734869707444284e-20

R14_167 V14 V167 5049.226891334893
L14_167 V14 V167 -4.869585186969094e-12
C14_167 V14 V167 -7.904377282800268e-21

R14_168 V14 V168 -1056.5118554816088
L14_168 V14 V168 -7.078805548575834e-12
C14_168 V14 V168 9.113062225547792e-20

R14_169 V14 V169 1228.4271064433137
L14_169 V14 V169 4.415264923216863e-12
C14_169 V14 V169 1.120767770143293e-19

R14_170 V14 V170 -678.0386985292207
L14_170 V14 V170 -8.5575141412335e-13
C14_170 V14 V170 -2.8690900996576617e-19

R14_171 V14 V171 11635.306881164339
L14_171 V14 V171 -2.7421350242095443e-12
C14_171 V14 V171 -3.384706839159057e-19

R14_172 V14 V172 1092.9470271406467
L14_172 V14 V172 -1.8428914013009714e-11
C14_172 V14 V172 -2.0838290195397615e-19

R14_173 V14 V173 -1465.2677466402026
L14_173 V14 V173 1.3016136545437149e-11
C14_173 V14 V173 2.3798814511459754e-19

R14_174 V14 V174 -947.4953184859049
L14_174 V14 V174 -1.4984204606324163e-12
C14_174 V14 V174 3.303366042613411e-19

R14_175 V14 V175 162749.79983322427
L14_175 V14 V175 8.269548361316072e-12
C14_175 V14 V175 3.6175845643310175e-20

R14_176 V14 V176 -12087.237200452148
L14_176 V14 V176 1.2169402080618128e-11
C14_176 V14 V176 8.845780201773863e-21

R14_177 V14 V177 1819.0888135419987
L14_177 V14 V177 -4.871314158699049e-12
C14_177 V14 V177 -1.3842185301571675e-19

R14_178 V14 V178 556.5253609627855
L14_178 V14 V178 8.537937462014161e-13
C14_178 V14 V178 6.604626882833554e-20

R14_179 V14 V179 -3284.852813096248
L14_179 V14 V179 2.4987755460384126e-12
C14_179 V14 V179 3.2094636326580117e-19

R14_180 V14 V180 9452.586942562635
L14_180 V14 V180 2.9089702650278074e-12
C14_180 V14 V180 2.4840014790793626e-19

R14_181 V14 V181 -14275.71839416186
L14_181 V14 V181 6.122862681100342e-12
C14_181 V14 V181 -1.2975081451085615e-20

R14_182 V14 V182 -2981.228383484411
L14_182 V14 V182 -1.744834870478211e-12
C14_182 V14 V182 -1.828301009847337e-19

R14_183 V14 V183 1138.2782670170996
L14_183 V14 V183 5.637428513864828e-12
C14_183 V14 V183 3.369194640931519e-20

R14_184 V14 V184 2314.0292013627613
L14_184 V14 V184 1.7038097318943425e-11
C14_184 V14 V184 -8.597569287122263e-20

R14_185 V14 V185 -3950.086126578146
L14_185 V14 V185 7.401510526492677e-12
C14_185 V14 V185 6.6659715985474e-20

R14_186 V14 V186 -1148.5191831776897
L14_186 V14 V186 -2.7554751276270678e-12
C14_186 V14 V186 1.5098292729153718e-20

R14_187 V14 V187 -1704.9894508231046
L14_187 V14 V187 -2.32975084304186e-12
C14_187 V14 V187 -2.891014389431819e-19

R14_188 V14 V188 -667.6167380862616
L14_188 V14 V188 -1.6948185196773147e-12
C14_188 V14 V188 -2.24387271210091e-19

R14_189 V14 V189 1759.0681987985508
L14_189 V14 V189 -6.7656650000268e-12
C14_189 V14 V189 -1.7479803713747472e-19

R14_190 V14 V190 871.07448454492
L14_190 V14 V190 3.944036281703814e-12
C14_190 V14 V190 1.933271304568279e-19

R14_191 V14 V191 -2547.512257709415
L14_191 V14 V191 -3.3388724365109017e-12
C14_191 V14 V191 -1.6691109358545967e-19

R14_192 V14 V192 2720.5076364678403
L14_192 V14 V192 9.746059130252373e-12
C14_192 V14 V192 -1.7468104768488665e-20

R14_193 V14 V193 -3292.220550365204
L14_193 V14 V193 1.522295704089366e-11
C14_193 V14 V193 1.4926655792524098e-19

R14_194 V14 V194 -2162.3866192144083
L14_194 V14 V194 -9.409634939444367e-12
C14_194 V14 V194 1.1853987637462082e-19

R14_195 V14 V195 1252.3220827691912
L14_195 V14 V195 1.3797378779669698e-12
C14_195 V14 V195 4.073829988911563e-19

R14_196 V14 V196 966.4910294993916
L14_196 V14 V196 1.4821792481470979e-12
C14_196 V14 V196 2.8454603053139126e-19

R14_197 V14 V197 -2213.706427432508
L14_197 V14 V197 8.126360284450875e-12
C14_197 V14 V197 6.57987719375987e-20

R14_198 V14 V198 -1607.0678396450785
L14_198 V14 V198 -5.7120113509582144e-12
C14_198 V14 V198 -6.880895877505021e-20

R14_199 V14 V199 4632.485460207744
L14_199 V14 V199 1.9340460347544033e-11
C14_199 V14 V199 1.6312380341564942e-19

R14_200 V14 V200 -1235.4993977899637
L14_200 V14 V200 -5.042744053427586e-12
C14_200 V14 V200 -4.7083400518542467e-20

R15_15 V15 0 -363.04169092890163
L15_15 V15 0 -3.68265484821125e-12
C15_15 V15 0 -5.75619600900809e-19

R15_16 V15 V16 -3050.702134279139
L15_16 V15 V16 -9.779039999152105e-13
C15_16 V15 V16 -5.664484541273758e-19

R15_17 V15 V17 36442.70547946566
L15_17 V15 V17 -5.1758244946825204e-11
C15_17 V15 V17 6.993710461125659e-20

R15_18 V15 V18 28396.68651003468
L15_18 V15 V18 -4.854014583857682e-12
C15_18 V15 V18 -8.996132352038301e-21

R15_19 V15 V19 -1457.477433966877
L15_19 V15 V19 6.376424917651686e-12
C15_19 V15 V19 3.2791187288166478e-19

R15_20 V15 V20 -3264.5626016737865
L15_20 V15 V20 -1.1488460923121427e-11
C15_20 V15 V20 1.407296232970152e-19

R15_21 V15 V21 -6533.005339187655
L15_21 V15 V21 -6.472655781729472e-12
C15_21 V15 V21 -3.7772584223581685e-20

R15_22 V15 V22 -3247.3886590103434
L15_22 V15 V22 3.267255058881294e-12
C15_22 V15 V22 1.6527134796613261e-19

R15_23 V15 V23 -1728.9274067029974
L15_23 V15 V23 1.2976613384005898e-12
C15_23 V15 V23 3.119573915587655e-19

R15_24 V15 V24 -3326.3958052578437
L15_24 V15 V24 1.1156612411575659e-11
C15_24 V15 V24 1.0095920979085354e-19

R15_25 V15 V25 6095.718913407179
L15_25 V15 V25 7.730583845599614e-12
C15_25 V15 V25 2.9121984821565625e-20

R15_26 V15 V26 3130.3971893253324
L15_26 V15 V26 -1.0562864533919996e-11
C15_26 V15 V26 -2.248033137852029e-20

R15_27 V15 V27 2833.4336592307523
L15_27 V15 V27 -3.1029370950800626e-12
C15_27 V15 V27 -2.821302603691475e-19

R15_28 V15 V28 3339.8493130333495
L15_28 V15 V28 4.328769537776355e-12
C15_28 V15 V28 2.8145497338639793e-20

R15_29 V15 V29 15817.900946350439
L15_29 V15 V29 2.5806922555822062e-12
C15_29 V15 V29 1.7624968563013584e-19

R15_30 V15 V30 5977.607579603452
L15_30 V15 V30 4.207686516692752e-11
C15_30 V15 V30 1.9738075636164295e-20

R15_31 V15 V31 777.5454202669462
L15_31 V15 V31 -4.083994252525558e-12
C15_31 V15 V31 -2.168827573875939e-19

R15_32 V15 V32 2042.832142043016
L15_32 V15 V32 6.22239598584136e-12
C15_32 V15 V32 -9.178164827131137e-20

R15_33 V15 V33 -9053.105160237568
L15_33 V15 V33 -1.3933151280916291e-12
C15_33 V15 V33 -2.6882941894019604e-19

R15_34 V15 V34 -7550.475553204466
L15_34 V15 V34 -3.55414952092668e-12
C15_34 V15 V34 9.848879931247408e-21

R15_35 V15 V35 -1914.7432358139893
L15_35 V15 V35 -8.422602577198952e-11
C15_35 V15 V35 2.172486240751123e-19

R15_36 V15 V36 -2645.92438486831
L15_36 V15 V36 -2.549757554318639e-12
C15_36 V15 V36 -1.8726343853390294e-19

R15_37 V15 V37 -15494.96993584837
L15_37 V15 V37 -4.42156802385083e-12
C15_37 V15 V37 -2.9201822354230824e-20

R15_38 V15 V38 -10127.42898616844
L15_38 V15 V38 -4.040639134388644e-12
C15_38 V15 V38 -1.1125050826158672e-19

R15_39 V15 V39 -1056.2812627644032
L15_39 V15 V39 2.0682997667682478e-12
C15_39 V15 V39 3.096664314690038e-19

R15_40 V15 V40 -1591.5899206650993
L15_40 V15 V40 2.145620557886002e-11
C15_40 V15 V40 1.48720611325279e-19

R15_41 V15 V41 6401.80897393564
L15_41 V15 V41 2.4961019585574057e-12
C15_41 V15 V41 2.319558499628892e-19

R15_42 V15 V42 8882.19491068675
L15_42 V15 V42 9.51090911796794e-12
C15_42 V15 V42 1.3310093588667664e-19

R15_43 V15 V43 -4230.02132088362
L15_43 V15 V43 -1.7196245819819665e-12
C15_43 V15 V43 -3.27641362665119e-19

R15_44 V15 V44 10035.554297672863
L15_44 V15 V44 9.225765784006986e-12
C15_44 V15 V44 -5.560479505216972e-20

R15_45 V15 V45 8704.583891064882
L15_45 V15 V45 3.179896009200769e-12
C15_45 V15 V45 9.008477681979766e-20

R15_46 V15 V46 4481.773983469251
L15_46 V15 V46 2.0613117555376745e-12
C15_46 V15 V46 2.030816760022065e-19

R15_47 V15 V47 1067.1516063831655
L15_47 V15 V47 -9.749257270681719e-11
C15_47 V15 V47 -1.2867826148655435e-19

R15_48 V15 V48 2284.8168396436095
L15_48 V15 V48 2.330149584129111e-12
C15_48 V15 V48 1.244027998463729e-19

R15_49 V15 V49 -12127.838100002944
L15_49 V15 V49 -3.6004416145562216e-12
C15_49 V15 V49 -8.299601857128228e-20

R15_50 V15 V50 35796.97744729958
L15_50 V15 V50 -2.312392814242551e-12
C15_50 V15 V50 -1.4951087838301638e-19

R15_51 V15 V51 2399.3534920481698
L15_51 V15 V51 2.7264193399189185e-12
C15_51 V15 V51 1.6131640355918818e-19

R15_52 V15 V52 -18009.1734275853
L15_52 V15 V52 -4.432745162286172e-12
C15_52 V15 V52 -1.3105569334713904e-19

R15_53 V15 V53 9095.09858398265
L15_53 V15 V53 -2.173955873833927e-12
C15_53 V15 V53 -2.0447852871475458e-19

R15_54 V15 V54 -26411.365142208026
L15_54 V15 V54 -2.47829019563018e-12
C15_54 V15 V54 -1.4824420236428057e-19

R15_55 V15 V55 -3215.524762890221
L15_55 V15 V55 1.2370443394402305e-11
C15_55 V15 V55 1.8448629997423146e-19

R15_56 V15 V56 -3475.8576655860784
L15_56 V15 V56 -2.1269938346284952e-12
C15_56 V15 V56 -2.0427077789615089e-19

R15_57 V15 V57 -12637.849892837345
L15_57 V15 V57 5.164002695095057e-12
C15_57 V15 V57 2.4832340591085057e-19

R15_58 V15 V58 4129.318562680848
L15_58 V15 V58 4.3521632257764945e-12
C15_58 V15 V58 1.3471070575645068e-19

R15_59 V15 V59 -2082.7056570938103
L15_59 V15 V59 -2.827318687644149e-12
C15_59 V15 V59 -9.604652402235813e-20

R15_60 V15 V60 -3892.9053192032984
L15_60 V15 V60 2.3457900995762306e-12
C15_60 V15 V60 2.0269424930624421e-19

R15_61 V15 V61 12236.923696222184
L15_61 V15 V61 3.0135059449895023e-12
C15_61 V15 V61 9.60756238172682e-20

R15_62 V15 V62 -5443.600397821989
L15_62 V15 V62 4.026258134271542e-12
C15_62 V15 V62 1.7113279690757128e-19

R15_63 V15 V63 91047.49327559912
L15_63 V15 V63 -3.840895118631353e-12
C15_63 V15 V63 -1.8309940566615153e-19

R15_64 V15 V64 5719.848163495112
L15_64 V15 V64 5.5069983620034494e-12
C15_64 V15 V64 4.26081129435889e-20

R15_65 V15 V65 27323.691144640477
L15_65 V15 V65 -5.250048135968318e-12
C15_65 V15 V65 -9.06546676301824e-20

R15_66 V15 V66 11307.279565615272
L15_66 V15 V66 -3.826646037065715e-12
C15_66 V15 V66 -6.966812180056779e-20

R15_67 V15 V67 2226.239883470271
L15_67 V15 V67 1.8747403409928856e-12
C15_67 V15 V67 2.44705779696796e-19

R15_68 V15 V68 4137.60736918334
L15_68 V15 V68 -6.60102522651901e-12
C15_68 V15 V68 -8.745316598460793e-20

R15_69 V15 V69 -39318.516702051915
L15_69 V15 V69 -4.349366915544413e-12
C15_69 V15 V69 -1.2510827063474404e-19

R15_70 V15 V70 10622.59762343009
L15_70 V15 V70 -8.677216793387389e-12
C15_70 V15 V70 -1.2550987602581962e-19

R15_71 V15 V71 2343.0998181629643
L15_71 V15 V71 -8.904956001778362e-12
C15_71 V15 V71 -1.6032468677473165e-19

R15_72 V15 V72 5112.252615578186
L15_72 V15 V72 8.151628228566953e-12
C15_72 V15 V72 1.882430408687027e-20

R15_73 V15 V73 4468.558004816736
L15_73 V15 V73 7.590223243817416e-12
C15_73 V15 V73 1.4749030951932055e-19

R15_74 V15 V74 -7035.003434426585
L15_74 V15 V74 1.3691455650559997e-11
C15_74 V15 V74 9.351702613360172e-20

R15_75 V15 V75 -1794.283776597152
L15_75 V15 V75 -1.87769461346131e-12
C15_75 V15 V75 -7.461013527022066e-20

R15_76 V15 V76 -2227.6449553989423
L15_76 V15 V76 -6.508671085228255e-12
C15_76 V15 V76 -9.678633911634654e-20

R15_77 V15 V77 -4922.89173571815
L15_77 V15 V77 -3.579004401044839e-11
C15_77 V15 V77 5.866948750631224e-20

R15_78 V15 V78 9591.664358954085
L15_78 V15 V78 -1.4664166034745856e-11
C15_78 V15 V78 -1.0131454830527804e-19

R15_79 V15 V79 -2028.458709364106
L15_79 V15 V79 2.336845511500401e-12
C15_79 V15 V79 1.8805193402222884e-19

R15_80 V15 V80 -4646.284961747446
L15_80 V15 V80 3.4955742460866236e-11
C15_80 V15 V80 6.010903865516613e-20

R15_81 V15 V81 19884.29795911146
L15_81 V15 V81 -1.909360781037075e-11
C15_81 V15 V81 -6.324084774106272e-20

R15_82 V15 V82 -37357.99291844696
L15_82 V15 V82 9.208185185814071e-12
C15_82 V15 V82 1.107363023560258e-19

R15_83 V15 V83 2866.5935795443024
L15_83 V15 V83 9.104589031265124e-12
C15_83 V15 V83 -2.2954781884710308e-20

R15_84 V15 V84 3839.374874231251
L15_84 V15 V84 3.6242546241017427e-12
C15_84 V15 V84 6.904467990413868e-20

R15_85 V15 V85 -358602.1058945014
L15_85 V15 V85 4.779926470375019e-12
C15_85 V15 V85 5.753510830270223e-20

R15_86 V15 V86 2882.773289556706
L15_86 V15 V86 5.589899272095837e-12
C15_86 V15 V86 8.706011849070341e-20

R15_87 V15 V87 1527.5945083135634
L15_87 V15 V87 -2.145504281251013e-12
C15_87 V15 V87 -2.892294875600447e-19

R15_88 V15 V88 8672.99114379041
L15_88 V15 V88 -6.8174192113973664e-12
C15_88 V15 V88 -1.9552298634655668e-19

R15_89 V15 V89 7306.631300287105
L15_89 V15 V89 -4.289132118929984e-12
C15_89 V15 V89 -9.315321048338666e-20

R15_90 V15 V90 -8734.243952851275
L15_90 V15 V90 -1.6914408469130676e-12
C15_90 V15 V90 -2.706832729701238e-19

R15_91 V15 V91 -6432.083006545446
L15_91 V15 V91 9.333367748946693e-13
C15_91 V15 V91 4.610023142706373e-19

R15_92 V15 V92 78529.56289227252
L15_92 V15 V92 3.6209704122660108e-12
C15_92 V15 V92 1.5801447724600688e-19

R15_93 V15 V93 15515.768678375276
L15_93 V15 V93 -5.2233673415280794e-12
C15_93 V15 V93 -6.06484673362821e-20

R15_94 V15 V94 -5334.055276619125
L15_94 V15 V94 1.7625163495936338e-11
C15_94 V15 V94 8.863584092603026e-20

R15_95 V15 V95 -824.9803109507917
L15_95 V15 V95 -3.1367608745938904e-12
C15_95 V15 V95 2.387013508559276e-20

R15_96 V15 V96 -1962.4881706372098
L15_96 V15 V96 -9.923733119409875e-12
C15_96 V15 V96 8.052552513932581e-20

R15_97 V15 V97 -2411.574502468296
L15_97 V15 V97 2.683369175342752e-12
C15_97 V15 V97 3.723430102051284e-19

R15_98 V15 V98 3335.436245851317
L15_98 V15 V98 2.300535461878721e-12
C15_98 V15 V98 2.121847143754306e-19

R15_99 V15 V99 799.2453644555708
L15_99 V15 V99 -1.0096663148424072e-12
C15_99 V15 V99 -4.877361798200942e-19

R15_100 V15 V100 5598.269437375442
L15_100 V15 V100 -2.2014993835482672e-11
C15_100 V15 V100 -2.3990237520367833e-19

R15_101 V15 V101 4497.689963755267
L15_101 V15 V101 -3.6289773226871842e-12
C15_101 V15 V101 -1.320414848167901e-19

R15_102 V15 V102 -5880.351200119776
L15_102 V15 V102 -3.99554761477966e-12
C15_102 V15 V102 -1.2032242502360397e-19

R15_103 V15 V103 -11779.760287417768
L15_103 V15 V103 9.088914820991343e-13
C15_103 V15 V103 4.422505137811545e-19

R15_104 V15 V104 3984.6444706505326
L15_104 V15 V104 4.615453973051693e-12
C15_104 V15 V104 1.0723135466934448e-19

R15_105 V15 V105 2680.6997231427413
L15_105 V15 V105 -3.682518823132169e-12
C15_105 V15 V105 -1.837230988709672e-19

R15_106 V15 V106 1626.1164985077817
L15_106 V15 V106 -2.8554113683152976e-12
C15_106 V15 V106 -2.178726554625593e-19

R15_107 V15 V107 -2365.0034297610437
L15_107 V15 V107 -4.485184961159364e-12
C15_107 V15 V107 -6.771650533515686e-20

R15_108 V15 V108 -35161.48441084053
L15_108 V15 V108 -8.458526141390096e-12
C15_108 V15 V108 3.891429200069723e-20

R15_109 V15 V109 -4542.5894470724115
L15_109 V15 V109 2.741348825112449e-12
C15_109 V15 V109 2.0895720819726081e-19

R15_110 V15 V110 -2149.2610723430616
L15_110 V15 V110 5.916608461912095e-12
C15_110 V15 V110 9.701407910224196e-20

R15_111 V15 V111 652.8848607437856
L15_111 V15 V111 -8.019099270760428e-12
C15_111 V15 V111 -1.448470920406154e-19

R15_112 V15 V112 2324.7230412424115
L15_112 V15 V112 5.5139884148079334e-11
C15_112 V15 V112 2.2930468126454607e-20

R15_113 V15 V113 -6650.122365265165
L15_113 V15 V113 -2.24523965299208e-11
C15_113 V15 V113 9.262804877954507e-20

R15_114 V15 V114 -1650.8965862187206
L15_114 V15 V114 2.8227529888834284e-12
C15_114 V15 V114 2.6522997381304025e-19

R15_115 V15 V115 -660.3171218742835
L15_115 V15 V115 -1.7784869285224403e-12
C15_115 V15 V115 6.968395407371975e-20

R15_116 V15 V116 -1341.78249180783
L15_116 V15 V116 -7.336018558675785e-12
C15_116 V15 V116 -9.645058037755554e-21

R15_117 V15 V117 -3885.914262003541
L15_117 V15 V117 -1.858400162049141e-12
C15_117 V15 V117 -8.851851954329717e-20

R15_118 V15 V118 1062.1079096818603
L15_118 V15 V118 -2.820822170439788e-12
C15_118 V15 V118 -3.382264887232612e-19

R15_119 V15 V119 1340.9078960052655
L15_119 V15 V119 4.4100442232467896e-12
C15_119 V15 V119 -5.719152223705097e-20

R15_120 V15 V120 2226.228378166757
L15_120 V15 V120 -1.1984358799072192e-11
C15_120 V15 V120 -1.8738780579021057e-19

R15_121 V15 V121 8046.081227009662
L15_121 V15 V121 8.78841175697351e-12
C15_121 V15 V121 -3.644779209313554e-20

R15_122 V15 V122 74675.7533444701
L15_122 V15 V122 2.3217083858447853e-11
C15_122 V15 V122 2.6154934865688663e-20

R15_123 V15 V123 1069.4048259092774
L15_123 V15 V123 1.3587469763324203e-12
C15_123 V15 V123 1.490304811665369e-19

R15_124 V15 V124 1713.8883740545173
L15_124 V15 V124 3.2335015678721213e-12
C15_124 V15 V124 2.655678664274935e-19

R15_125 V15 V125 1208.785497467888
L15_125 V15 V125 2.322720368717693e-12
C15_125 V15 V125 -2.9492103931124414e-20

R15_126 V15 V126 -3818.134656659761
L15_126 V15 V126 1.9558377564546246e-12
C15_126 V15 V126 2.1623169507688999e-19

R15_127 V15 V127 -792.520453526888
L15_127 V15 V127 -1.028486009897956e-12
C15_127 V15 V127 -1.3281698185526964e-19

R15_128 V15 V128 -1329.4118455663315
L15_128 V15 V128 -1.6857208086693964e-11
C15_128 V15 V128 7.856155415819016e-20

R15_129 V15 V129 -1174.274006925098
L15_129 V15 V129 -4.442375763569044e-12
C15_129 V15 V129 1.947130635310563e-19

R15_130 V15 V130 -2360.4044940865306
L15_130 V15 V130 -2.435935991800596e-12
C15_130 V15 V130 -1.684468997715786e-19

R15_131 V15 V131 1789.899602580352
L15_131 V15 V131 2.704307957842841e-12
C15_131 V15 V131 -1.4543878245482682e-20

R15_132 V15 V132 2138.346822902746
L15_132 V15 V132 -3.98805012045566e-12
C15_132 V15 V132 -3.3670357711186544e-19

R15_133 V15 V133 -1755.9148113816889
L15_133 V15 V133 -2.3258902297596324e-12
C15_133 V15 V133 -1.0198234690152757e-19

R15_134 V15 V134 4262.6401000157675
L15_134 V15 V134 2.979067471093756e-12
C15_134 V15 V134 -1.0287464243287899e-20

R15_135 V15 V135 1795.526955857982
L15_135 V15 V135 9.520996005957731e-13
C15_135 V15 V135 3.2475751877411584e-19

R15_136 V15 V136 1941.7584636670156
L15_136 V15 V136 3.8394740553631135e-12
C15_136 V15 V136 2.0817361085126077e-19

R15_137 V15 V137 1069.444670862823
L15_137 V15 V137 2.6793667601418743e-12
C15_137 V15 V137 -8.424388857477251e-20

R15_138 V15 V138 -5071.137053142428
L15_138 V15 V138 6.615331918347263e-12
C15_138 V15 V138 1.129678390085945e-19

R15_139 V15 V139 -1028.2162197873647
L15_139 V15 V139 -5.727727367933321e-13
C15_139 V15 V139 -5.364545903031022e-19

R15_140 V15 V140 -1022.1269008545947
L15_140 V15 V140 -2.819139733292647e-12
C15_140 V15 V140 -1.762626469066019e-19

R15_141 V15 V141 1326.7310297765844
L15_141 V15 V141 1.4844619742839274e-12
C15_141 V15 V141 2.321659805728685e-19

R15_142 V15 V142 -3496.2172100928387
L15_142 V15 V142 -1.5386655265413127e-12
C15_142 V15 V142 -1.7290232869263884e-20

R15_143 V15 V143 1259.971074586634
L15_143 V15 V143 -2.0277192111114155e-11
C15_143 V15 V143 1.86702463753303e-19

R15_144 V15 V144 2458.2147274743766
L15_144 V15 V144 -9.227463870088945e-11
C15_144 V15 V144 2.5518173497141354e-20

R15_145 V15 V145 -823.9642778979974
L15_145 V15 V145 -1.720450918615186e-12
C15_145 V15 V145 6.030433100922351e-20

R15_146 V15 V146 2150.3392566980283
L15_146 V15 V146 3.9366336834920576e-12
C15_146 V15 V146 -5.82352084171897e-20

R15_147 V15 V147 -528.5530981019552
L15_147 V15 V147 7.255205871743591e-13
C15_147 V15 V147 3.705322647032325e-19

R15_148 V15 V148 -6893.616165984601
L15_148 V15 V148 6.366340390375283e-12
C15_148 V15 V148 1.4727605149322846e-19

R15_149 V15 V149 -47336.57825494568
L15_149 V15 V149 -9.593464905089888e-13
C15_149 V15 V149 -4.0202401452954146e-19

R15_150 V15 V150 979.830603877302
L15_150 V15 V150 1.4860547429252791e-12
C15_150 V15 V150 1.6389288577059577e-19

R15_151 V15 V151 245.68262610729977
L15_151 V15 V151 2.419870615120325e-12
C15_151 V15 V151 -2.0000178082190274e-19

R15_152 V15 V152 4449.358525314393
L15_152 V15 V152 -2.027342537240272e-11
C15_152 V15 V152 -1.0647728176838771e-20

R15_153 V15 V153 4384.602501560767
L15_153 V15 V153 1.8308055013901148e-12
C15_153 V15 V153 4.0737678213917104e-20

R15_154 V15 V154 -3832.50262563645
L15_154 V15 V154 -6.354800773026825e-12
C15_154 V15 V154 -5.562891919609413e-20

R15_155 V15 V155 -127.74017235312303
L15_155 V15 V155 -6.137050196469265e-13
C15_155 V15 V155 -3.467311118764911e-19

R15_156 V15 V156 2344.8313590252883
L15_156 V15 V156 2.9884661427666064e-11
C15_156 V15 V156 -1.167578835085363e-19

R15_157 V15 V157 3668.641661837064
L15_157 V15 V157 1.1120140303393102e-12
C15_157 V15 V157 4.2756542292775996e-19

R15_158 V15 V158 4523.8279980873585
L15_158 V15 V158 -2.6211593296456997e-12
C15_158 V15 V158 -6.654318820963248e-20

R15_159 V15 V159 383.71090008697865
L15_159 V15 V159 -1.0922753715914119e-11
C15_159 V15 V159 3.0932302795976905e-19

R15_160 V15 V160 -3620.820173160584
L15_160 V15 V160 9.663710899503925e-12
C15_160 V15 V160 1.1771404586616163e-20

R15_161 V15 V161 -5411.145089599862
L15_161 V15 V161 -2.839493803055434e-12
C15_161 V15 V161 -1.5547353078834408e-19

R15_162 V15 V162 6561.725796163748
L15_162 V15 V162 -4.597712217255551e-12
C15_162 V15 V162 -3.144709785164511e-20

R15_163 V15 V163 560.9381031951258
L15_163 V15 V163 1.0017916330127298e-12
C15_163 V15 V163 -4.2039048058270843e-20

R15_164 V15 V164 993.2481358861706
L15_164 V15 V164 9.919264634477085e-12
C15_164 V15 V164 -4.85186524308254e-20

R15_165 V15 V165 2883.878638499196
L15_165 V15 V165 -3.538683986171261e-12
C15_165 V15 V165 -1.116423180075884e-19

R15_166 V15 V166 4712.645786939695
L15_166 V15 V166 2.0849048123547786e-12
C15_166 V15 V166 7.997628425843186e-20

R15_167 V15 V167 3305.345726265702
L15_167 V15 V167 -1.6862203438286836e-11
C15_167 V15 V167 -6.190152828386046e-20

R15_168 V15 V168 -895.8358225496919
L15_168 V15 V168 -6.991881159840781e-12
C15_168 V15 V168 -1.8110977417860814e-20

R15_169 V15 V169 1937.8447586977377
L15_169 V15 V169 3.598239790112593e-12
C15_169 V15 V169 1.731530438949319e-19

R15_170 V15 V170 3034.3017174759652
L15_170 V15 V170 -2.970173098986709e-12
C15_170 V15 V170 -1.111940782447214e-19

R15_171 V15 V171 -331.74667674330794
L15_171 V15 V171 -1.1051655354006227e-12
C15_171 V15 V171 -6.83129140963389e-20

R15_172 V15 V172 -3561.3994248171794
L15_172 V15 V172 -5.70601400781402e-12
C15_172 V15 V172 -3.3302430518629775e-20

R15_173 V15 V173 -1994.8331553027335
L15_173 V15 V173 -4.839156960809972e-12
C15_173 V15 V173 3.013574748140454e-20

R15_174 V15 V174 -988.3798915012806
L15_174 V15 V174 -3.308400846899771e-12
C15_174 V15 V174 1.3526231618340132e-19

R15_175 V15 V175 506.58994536238123
L15_175 V15 V175 -1.1127946023160949e-11
C15_175 V15 V175 -1.103125520133046e-19

R15_176 V15 V176 39034.609684984316
L15_176 V15 V176 1.099942755152479e-10
C15_176 V15 V176 -1.9610388473197336e-20

R15_177 V15 V177 1391.8191267166878
L15_177 V15 V177 8.467286067943164e-12
C15_177 V15 V177 -3.996881931142994e-20

R15_178 V15 V178 1502.154188509652
L15_178 V15 V178 1.9252966111780106e-12
C15_178 V15 V178 4.206187715929711e-20

R15_179 V15 V179 -645.4332950051236
L15_179 V15 V179 1.1321477805830821e-12
C15_179 V15 V179 2.168591156570685e-19

R15_180 V15 V180 2046.1157998298572
L15_180 V15 V180 2.172286561425036e-12
C15_180 V15 V180 1.450801073473564e-19

R15_181 V15 V181 -3254.4666070697626
L15_181 V15 V181 -1.3208570683775425e-11
C15_181 V15 V181 -4.27503083063394e-20

R15_182 V15 V182 -1570.5359535554003
L15_182 V15 V182 -2.2284684021216278e-12
C15_182 V15 V182 -1.1733944582880702e-19

R15_183 V15 V183 629.6726449032298
L15_183 V15 V183 5.8954414909211595e-12
C15_183 V15 V183 5.484405494997768e-20

R15_184 V15 V184 5433.342177963162
L15_184 V15 V184 1.0726190789881241e-11
C15_184 V15 V184 -4.117176410709059e-20

R15_185 V15 V185 -3168.1132137264017
L15_185 V15 V185 -4.0696860666731616e-11
C15_185 V15 V185 2.931793931480886e-20

R15_186 V15 V186 -4238.155865826055
L15_186 V15 V186 -9.141200304402746e-12
C15_186 V15 V186 -7.409290974663839e-22

R15_187 V15 V187 -7124.89701207373
L15_187 V15 V187 -1.2524762869213749e-12
C15_187 V15 V187 -2.542351752699042e-19

R15_188 V15 V188 -704.3010401376756
L15_188 V15 V188 -1.5921152270628434e-12
C15_188 V15 V188 -1.416915283057673e-19

R15_189 V15 V189 1639.4310481989835
L15_189 V15 V189 7.03155761830888e-12
C15_189 V15 V189 1.6305190590943475e-20

R15_190 V15 V190 1616.518711003153
L15_190 V15 V190 4.833007405446021e-12
C15_190 V15 V190 1.0318981392559245e-19

R15_191 V15 V191 -1136.4359697842697
L15_191 V15 V191 -2.218759138956251e-11
C15_191 V15 V191 5.1447092677534894e-20

R15_192 V15 V192 6109.332440236892
L15_192 V15 V192 9.248667546360035e-11
C15_192 V15 V192 9.354420305250977e-20

R15_193 V15 V193 -13480.148232409147
L15_193 V15 V193 4.659870949081879e-11
C15_193 V15 V193 6.714523964709025e-20

R15_194 V15 V194 -2852.0210273179205
L15_194 V15 V194 6.328876016780293e-12
C15_194 V15 V194 1.3856279190238718e-19

R15_195 V15 V195 1336.411623209165
L15_195 V15 V195 9.361279508094089e-12
C15_195 V15 V195 -2.8953257762912416e-20

R15_196 V15 V196 554.4481907967687
L15_196 V15 V196 1.298126971774987e-12
C15_196 V15 V196 7.312705405316411e-20

R15_197 V15 V197 -32953.379921149564
L15_197 V15 V197 -9.623511536268294e-12
C15_197 V15 V197 -8.26712712500604e-20

R15_198 V15 V198 2533.08076590676
L15_198 V15 V198 -5.039318836703379e-12
C15_198 V15 V198 -2.8696785305854936e-21

R15_199 V15 V199 5529.263349515481
L15_199 V15 V199 -4.3002510575561526e-11
C15_199 V15 V199 5.516127820917462e-20

R15_200 V15 V200 -1515.0771381824304
L15_200 V15 V200 -2.66163167224248e-12
C15_200 V15 V200 -1.2276051703116914e-19

R16_16 V16 0 -172.5935068636525
L16_16 V16 0 -4.5062105672473887e-13
C16_16 V16 0 -9.338260015016283e-19

R16_17 V16 V17 -120800.50638179117
L16_17 V16 V17 -2.9685262698375804e-11
C16_17 V16 V17 7.545829338067049e-20

R16_18 V16 V18 -71835.85311092332
L16_18 V16 V18 -3.6565228960957006e-12
C16_18 V16 V18 -6.3799425067686675e-21

R16_19 V16 V19 -5716.006993963141
L16_19 V16 V19 -1.2841857767650654e-10
C16_19 V16 V19 1.2141646331856542e-19

R16_20 V16 V20 -1171.6090265947948
L16_20 V16 V20 1.6793527202047054e-11
C16_20 V16 V20 3.2950815059095855e-19

R16_21 V16 V21 -3130.4189069477097
L16_21 V16 V21 -3.4273624564986837e-12
C16_21 V16 V21 -5.3973019792244156e-20

R16_22 V16 V22 -2853.6266778662225
L16_22 V16 V22 3.0905021629340726e-12
C16_22 V16 V22 1.876351984305703e-19

R16_23 V16 V23 -4077.248904706127
L16_23 V16 V23 8.257226316533345e-11
C16_23 V16 V23 4.55583328856904e-20

R16_24 V16 V24 -1672.5019394766234
L16_24 V16 V24 1.4942012179659626e-12
C16_24 V16 V24 3.870274419693453e-19

R16_25 V16 V25 3638.5120109757963
L16_25 V16 V25 4.6222154362994676e-12
C16_25 V16 V25 6.399469876243665e-20

R16_26 V16 V26 3028.531720199151
L16_26 V16 V26 -2.0537270848157734e-11
C16_26 V16 V26 2.0495349090985953e-20

R16_27 V16 V27 3968.1329091518733
L16_27 V16 V27 5.830220746307187e-12
C16_27 V16 V27 6.924741168562043e-20

R16_28 V16 V28 2345.3616286645984
L16_28 V16 V28 1.4822162979519242e-11
C16_28 V16 V28 -3.001162101031104e-19

R16_29 V16 V29 5472.69881563478
L16_29 V16 V29 1.7350265933462666e-12
C16_29 V16 V29 2.1768229978912e-19

R16_30 V16 V30 5185.790271559923
L16_30 V16 V30 1.1780223014776284e-11
C16_30 V16 V30 1.0266283590005147e-20

R16_31 V16 V31 2573.2809932348423
L16_31 V16 V31 7.545388827203329e-12
C16_31 V16 V31 4.24785016841407e-21

R16_32 V16 V32 709.9495818890072
L16_32 V16 V32 2.0868768374211434e-09
C16_32 V16 V32 -2.373275672455189e-19

R16_33 V16 V33 -7654.572692456552
L16_33 V16 V33 -1.0671223504579109e-12
C16_33 V16 V33 -3.2365822267019486e-19

R16_34 V16 V34 -4527.917529264442
L16_34 V16 V34 -2.874079316981834e-12
C16_34 V16 V34 2.2785432058318122e-20

R16_35 V16 V35 -5029.2213359086645
L16_35 V16 V35 -2.0171086859814266e-12
C16_35 V16 V35 -7.029740640055602e-20

R16_36 V16 V36 -1205.1238775595139
L16_36 V16 V36 -4.115983838258583e-12
C16_36 V16 V36 -3.639100509448885e-21

R16_37 V16 V37 -6805.82422061943
L16_37 V16 V37 -2.7841745261452728e-12
C16_37 V16 V37 -6.384068752745479e-20

R16_38 V16 V38 -6216.898985613768
L16_38 V16 V38 -2.608240249044271e-12
C16_38 V16 V38 -1.4661193059381898e-19

R16_39 V16 V39 -2509.3113144404756
L16_39 V16 V39 -1.6226409048940803e-11
C16_39 V16 V39 5.845284807134928e-20

R16_40 V16 V40 -838.0258771671175
L16_40 V16 V40 2.2160043318919868e-12
C16_40 V16 V40 2.84162111867963e-19

R16_41 V16 V41 5830.319155117949
L16_41 V16 V41 1.7436092956838288e-12
C16_41 V16 V41 3.021897135173732e-19

R16_42 V16 V42 10201.91217291977
L16_42 V16 V42 5.290380430592675e-12
C16_42 V16 V42 1.6218767395276036e-19

R16_43 V16 V43 6473.479669994769
L16_43 V16 V43 5.587954317224114e-11
C16_43 V16 V43 5.112595349767858e-20

R16_44 V16 V44 -6758.641753541043
L16_44 V16 V44 -2.286535005845644e-12
C16_44 V16 V44 -3.164362078112987e-19

R16_45 V16 V45 4989.7550506226335
L16_45 V16 V45 2.1363659326856386e-12
C16_45 V16 V45 1.101417492308187e-19

R16_46 V16 V46 3554.776950377216
L16_46 V16 V46 1.4094483619208672e-12
C16_46 V16 V46 2.5896695320804534e-19

R16_47 V16 V47 2965.7931509754067
L16_47 V16 V47 2.5424380488846127e-12
C16_47 V16 V47 9.476798940148406e-20

R16_48 V16 V48 793.3139300313393
L16_48 V16 V48 2.686408626921759e-12
C16_48 V16 V48 -5.3975147564343354e-20

R16_49 V16 V49 -13148.262857028512
L16_49 V16 V49 -2.848043326131665e-12
C16_49 V16 V49 -9.541065238874982e-20

R16_50 V16 V50 -24559.949920894825
L16_50 V16 V50 -1.7567708268607138e-12
C16_50 V16 V50 -1.7426813903646822e-19

R16_51 V16 V51 14280.97637008561
L16_51 V16 V51 -2.85185258497595e-12
C16_51 V16 V51 -1.141777421996443e-19

R16_52 V16 V52 9010.216913560924
L16_52 V16 V52 3.0879376053395374e-12
C16_52 V16 V52 9.192610934994818e-20

R16_53 V16 V53 9886.907445965939
L16_53 V16 V53 -1.6825240159577542e-12
C16_53 V16 V53 -2.378116169667254e-19

R16_54 V16 V54 -8008.140759566976
L16_54 V16 V54 -1.7945255863698078e-12
C16_54 V16 V54 -1.8426337213203134e-19

R16_55 V16 V55 -43645.22045042748
L16_55 V16 V55 -2.5896485209605345e-12
C16_55 V16 V55 -1.0685826904399534e-19

R16_56 V16 V56 -1300.135764288366
L16_56 V16 V56 -2.976178227774622e-12
C16_56 V16 V56 -3.485147638095268e-20

R16_57 V16 V57 -8986.35555536624
L16_57 V16 V57 4.182578758801154e-12
C16_57 V16 V57 2.7453043223707984e-19

R16_58 V16 V58 3643.682143554625
L16_58 V16 V58 2.812475728992856e-12
C16_58 V16 V58 1.6643348774756484e-19

R16_59 V16 V59 -7373.7414692906605
L16_59 V16 V59 2.4518447575359636e-12
C16_59 V16 V59 2.5835537258275313e-19

R16_60 V16 V60 -1723.4660747378812
L16_60 V16 V60 -8.564723950378843e-12
C16_60 V16 V60 1.5245135213841423e-21

R16_61 V16 V61 8506.168520813217
L16_61 V16 V61 2.1699859746861474e-12
C16_61 V16 V61 1.2446534535810717e-19

R16_62 V16 V62 -5911.560014959706
L16_62 V16 V62 2.9757099627774513e-12
C16_62 V16 V62 1.7762718784793534e-19

R16_63 V16 V63 11329.322316769745
L16_63 V16 V63 -8.2479080799435e-11
C16_63 V16 V63 -4.111615677084291e-21

R16_64 V16 V64 4283.533355239415
L16_64 V16 V64 2.3278527416483957e-11
C16_64 V16 V64 -2.264385221366602e-19

R16_65 V16 V65 11643.22773350044
L16_65 V16 V65 -4.9226040731154176e-12
C16_65 V16 V65 -1.0421932250197953e-19

R16_66 V16 V66 28984.587721732954
L16_66 V16 V66 -3.0420280482726564e-12
C16_66 V16 V66 -5.422533363245634e-20

R16_67 V16 V67 -43796.81383199425
L16_67 V16 V67 -2.0062386767925224e-12
C16_67 V16 V67 -1.8460452506404698e-19

R16_68 V16 V68 1669.2724187454426
L16_68 V16 V68 1.4565864599401738e-12
C16_68 V16 V68 2.226207748925432e-19

R16_69 V16 V69 -13510.633988528034
L16_69 V16 V69 -3.0953728697191376e-12
C16_69 V16 V69 -1.330245442116044e-19

R16_70 V16 V70 10007.985280671217
L16_70 V16 V70 -7.029360598240399e-12
C16_70 V16 V70 -1.2491936693070608e-19

R16_71 V16 V71 7493.226698072833
L16_71 V16 V71 2.148165737844155e-12
C16_71 V16 V71 1.109905063436381e-19

R16_72 V16 V72 2059.6834269546002
L16_72 V16 V72 -5.129218824004921e-12
C16_72 V16 V72 -1.6498628499285292e-19

R16_73 V16 V73 4732.43904787204
L16_73 V16 V73 4.730394040875985e-12
C16_73 V16 V73 1.814074178495078e-19

R16_74 V16 V74 -5642.140163005811
L16_74 V16 V74 1.1335542980808056e-11
C16_74 V16 V74 6.30999231219721e-20

R16_75 V16 V75 12754.267708743073
L16_75 V16 V75 3.0070682237773234e-11
C16_75 V16 V75 7.059534731190095e-20

R16_76 V16 V76 -828.6625662402762
L16_76 V16 V76 -9.460811306521368e-13
C16_76 V16 V76 -2.373533218569201e-19

R16_77 V16 V77 -5516.754706717355
L16_77 V16 V77 -2.3002120180905318e-11
C16_77 V16 V77 4.257596524281636e-20

R16_78 V16 V78 4884.70301039368
L16_78 V16 V78 -1.0865171184739792e-11
C16_78 V16 V78 -7.649738693949159e-20

R16_79 V16 V79 -2945.170164165716
L16_79 V16 V79 -2.9415925056405846e-12
C16_79 V16 V79 -8.255590811881486e-20

R16_80 V16 V80 -24554.836418030747
L16_80 V16 V80 1.0072833568023257e-12
C16_80 V16 V80 3.811360322141224e-19

R16_81 V16 V81 4488.912567545307
L16_81 V16 V81 -3.992390358056699e-11
C16_81 V16 V81 -3.316811564661146e-20

R16_82 V16 V82 -30477.819254033107
L16_82 V16 V82 6.4515165530681656e-12
C16_82 V16 V82 1.3698358795509596e-19

R16_83 V16 V83 5383.98635332204
L16_83 V16 V83 -1.1641879677855051e-11
C16_83 V16 V83 2.850925898426905e-20

R16_84 V16 V84 2264.3075862346295
L16_84 V16 V84 2.5126966473071095e-12
C16_84 V16 V84 -8.694931086232931e-20

R16_85 V16 V85 -51896.81648302331
L16_85 V16 V85 3.640056463563902e-12
C16_85 V16 V85 5.957979185804172e-20

R16_86 V16 V86 4282.932814092398
L16_86 V16 V86 5.624383603686733e-12
C16_86 V16 V86 4.807856709822295e-20

R16_87 V16 V87 9863.561037670846
L16_87 V16 V87 -1.0106501278299895e-11
C16_87 V16 V87 -1.2283911323056656e-19

R16_88 V16 V88 1744.1407210012667
L16_88 V16 V88 -1.1645089947103586e-12
C16_88 V16 V88 -3.1908908769811006e-19

R16_89 V16 V89 19681.37766383126
L16_89 V16 V89 -2.2056501380539195e-12
C16_89 V16 V89 -1.1316935634809825e-19

R16_90 V16 V90 -6636.824201499539
L16_90 V16 V90 -1.1360947414655854e-12
C16_90 V16 V90 -2.706822270375219e-19

R16_91 V16 V91 3048.4259613692957
L16_91 V16 V91 1.5726565499660124e-12
C16_91 V16 V91 2.5256571233677764e-19

R16_92 V16 V92 -2174.964525167858
L16_92 V16 V92 7.200238078358471e-13
C16_92 V16 V92 4.10851176993551e-19

R16_93 V16 V93 5375.066517401207
L16_93 V16 V93 -4.42745091901054e-12
C16_93 V16 V93 -4.7980482266077754e-20

R16_94 V16 V94 -13135.173190442847
L16_94 V16 V94 7.162579783253434e-12
C16_94 V16 V94 1.2977476844723055e-19

R16_95 V16 V95 -2983.4411169959444
L16_95 V16 V95 -1.1588849261494454e-11
C16_95 V16 V95 5.750716835364675e-20

R16_96 V16 V96 -673.7420363805775
L16_96 V16 V96 -1.4378555929258874e-12
C16_96 V16 V96 -1.1301013459879041e-20

R16_97 V16 V97 -2442.158844999512
L16_97 V16 V97 1.6734101442182467e-12
C16_97 V16 V97 3.937257062053275e-19

R16_98 V16 V98 3971.9460520828757
L16_98 V16 V98 1.5680697043856977e-12
C16_98 V16 V98 1.994032606756538e-19

R16_99 V16 V99 -10733.811846383165
L16_99 V16 V99 -1.1371527905714836e-12
C16_99 V16 V99 -2.844177063990959e-19

R16_100 V16 V100 524.4428619396538
L16_100 V16 V100 -2.7776034268023524e-12
C16_100 V16 V100 -4.3357827667591076e-19

R16_101 V16 V101 4368.255944170581
L16_101 V16 V101 -2.2533698726057985e-12
C16_101 V16 V101 -1.3601413138362557e-19

R16_102 V16 V102 -4401.3678846367575
L16_102 V16 V102 -2.5352047181668724e-12
C16_102 V16 V102 -1.3590916953608434e-19

R16_103 V16 V103 3416.166992242909
L16_103 V16 V103 4.054515294476169e-12
C16_103 V16 V103 6.720327559614049e-20

R16_104 V16 V104 -7692.369785101834
L16_104 V16 V104 7.917561675224083e-13
C16_104 V16 V104 4.2603465199816285e-19

R16_105 V16 V105 2248.6906332031986
L16_105 V16 V105 -2.7378939172888895e-12
C16_105 V16 V105 -2.0200078022333597e-19

R16_106 V16 V106 1390.5469773356785
L16_106 V16 V106 -2.9887167391958595e-12
C16_106 V16 V106 -1.72878324719802e-19

R16_107 V16 V107 6429.57091671247
L16_107 V16 V107 2.4122755629268734e-12
C16_107 V16 V107 1.7992762034999367e-19

R16_108 V16 V108 -1007.364956700831
L16_108 V16 V108 -9.104902508575305e-13
C16_108 V16 V108 -1.9357329921116442e-19

R16_109 V16 V109 -1996.916014796325
L16_109 V16 V109 2.302959047549765e-12
C16_109 V16 V109 2.2547047958097385e-19

R16_110 V16 V110 -1569.1053208784654
L16_110 V16 V110 1.4701445390945806e-11
C16_110 V16 V110 5.839905435855526e-20

R16_111 V16 V111 2699.8217130352987
L16_111 V16 V111 1.906342467373936e-11
C16_111 V16 V111 -5.1009435545001284e-20

R16_112 V16 V112 712.1558313012167
L16_112 V16 V112 2.915921245487204e-12
C16_112 V16 V112 -2.5860846729367552e-20

R16_113 V16 V113 15773.289680035956
L16_113 V16 V113 9.950730814525156e-12
C16_113 V16 V113 1.323877401680683e-19

R16_114 V16 V114 -1767.2346560589085
L16_114 V16 V114 1.8203515001227908e-12
C16_114 V16 V114 2.605803025439666e-19

R16_115 V16 V115 -909.8660587730142
L16_115 V16 V115 -1.8967433426992657e-12
C16_115 V16 V115 -1.2763555412839865e-19

R16_116 V16 V116 -942.2656007204583
L16_116 V16 V116 -3.4622352481976527e-12
C16_116 V16 V116 1.588331707452306e-19

R16_117 V16 V117 -5158.693467509823
L16_117 V16 V117 -1.4065636731114906e-12
C16_117 V16 V117 -1.3347694501480468e-19

R16_118 V16 V118 910.9880732372612
L16_118 V16 V118 -3.392484514159778e-12
C16_118 V16 V118 -3.146486417041215e-19

R16_119 V16 V119 2144.518369683554
L16_119 V16 V119 -6.10044412900391e-10
C16_119 V16 V119 -1.1595591019564074e-19

R16_120 V16 V120 982.3376741937703
L16_120 V16 V120 -3.937517312431287e-12
C16_120 V16 V120 -2.8995333017633768e-19

R16_121 V16 V121 -8339.468859970739
L16_121 V16 V121 1.918725167669736e-11
C16_121 V16 V121 -5.2331496265742313e-20

R16_122 V16 V122 -7154.188726442807
L16_122 V16 V122 -2.3043576965489368e-11
C16_122 V16 V122 2.594891033099106e-20

R16_123 V16 V123 1556.844132068852
L16_123 V16 V123 2.111199910430598e-12
C16_123 V16 V123 1.833320634105062e-19

R16_124 V16 V124 4351.064359259777
L16_124 V16 V124 7.277047417247679e-13
C16_124 V16 V124 3.5590950259060015e-19

R16_125 V16 V125 1106.6177076014283
L16_125 V16 V125 1.567090027746459e-12
C16_125 V16 V125 -5.995387473058093e-21

R16_126 V16 V126 -3870.5133686856516
L16_126 V16 V126 1.4120985439506448e-12
C16_126 V16 V126 1.883694586234151e-19

R16_127 V16 V127 -1128.20891552274
L16_127 V16 V127 4.52113064293121e-12
C16_127 V16 V127 1.3650134415578472e-19

R16_128 V16 V128 -764.9228058634063
L16_128 V16 V128 -9.39140942685835e-13
C16_128 V16 V128 -2.734556517434149e-20

R16_129 V16 V129 -1140.4543299545687
L16_129 V16 V129 -4.095165615010317e-12
C16_129 V16 V129 2.4505129359787595e-19

R16_130 V16 V130 -2976.6780065871394
L16_130 V16 V130 -1.8386111307286052e-12
C16_130 V16 V130 -1.8644386042218574e-19

R16_131 V16 V131 1286.356164592335
L16_131 V16 V131 -2.6669642562035515e-12
C16_131 V16 V131 -2.4599417660109535e-19

R16_132 V16 V132 824.0908904340548
L16_132 V16 V132 1.709818740603531e-11
C16_132 V16 V132 -2.857469249683312e-19

R16_133 V16 V133 -2519.768444519337
L16_133 V16 V133 -1.7025340657942558e-12
C16_133 V16 V133 -1.7053976556982085e-19

R16_134 V16 V134 2006.6598026424986
L16_134 V16 V134 2.2882924153274244e-12
C16_134 V16 V134 2.78557319228292e-20

R16_135 V16 V135 15997.02747508695
L16_135 V16 V135 5.526817081962106e-12
C16_135 V16 V135 9.744469054058347e-21

R16_136 V16 V136 1714.9945888501193
L16_136 V16 V136 6.954264818308986e-13
C16_136 V16 V136 4.415311760159831e-19

R16_137 V16 V137 1320.2072355334758
L16_137 V16 V137 2.0434292453296824e-12
C16_137 V16 V137 -1.276814031913412e-19

R16_138 V16 V138 -2212.3637323165567
L16_138 V16 V138 4.45795959151742e-12
C16_138 V16 V138 8.669948502528505e-20

R16_139 V16 V139 -850.4150132647147
L16_139 V16 V139 -3.6614674908280105e-12
C16_139 V16 V139 -2.9665576608916355e-20

R16_140 V16 V140 -1716.7766832671116
L16_140 V16 V140 -5.79945973097486e-13
C16_140 V16 V140 -5.113664308146166e-19

R16_141 V16 V141 1681.6456215006008
L16_141 V16 V141 9.98914320041717e-13
C16_141 V16 V141 3.2821729978370423e-19

R16_142 V16 V142 -1868.5754037180336
L16_142 V16 V142 -1.2492489949537445e-12
C16_142 V16 V142 -4.05374714611199e-20

R16_143 V16 V143 1034.5460057619543
L16_143 V16 V143 2.856183766073592e-12
C16_143 V16 V143 1.2312331674126638e-19

R16_144 V16 V144 -600.0321057122989
L16_144 V16 V144 -3.0832104538023647e-12
C16_144 V16 V144 8.29102049257635e-20

R16_145 V16 V145 -970.7189043318502
L16_145 V16 V145 -1.3302017608561303e-12
C16_145 V16 V145 1.0692949243406431e-19

R16_146 V16 V146 2188.1979512777098
L16_146 V16 V146 4.775832761524581e-12
C16_146 V16 V146 -4.255213563271701e-20

R16_147 V16 V147 -1549.9332317530818
L16_147 V16 V147 2.538364200879918e-12
C16_147 V16 V147 1.3104544430550857e-19

R16_148 V16 V148 275.77604284200737
L16_148 V16 V148 4.881469261042217e-13
C16_148 V16 V148 4.421157854714705e-19

R16_149 V16 V149 -9401.492065530056
L16_149 V16 V149 -7.175825905803382e-13
C16_149 V16 V149 -5.505408030382445e-19

R16_150 V16 V150 796.7395032088149
L16_150 V16 V150 1.0260095713160224e-12
C16_150 V16 V150 2.600252815773586e-19

R16_151 V16 V151 3010.942802119762
L16_151 V16 V151 -2.5268196070392288e-12
C16_151 V16 V151 -1.0762410995978064e-19

R16_152 V16 V152 -999.7988597044242
L16_152 V16 V152 3.1028181126208637e-10
C16_152 V16 V152 -1.5841105056248084e-19

R16_153 V16 V153 -8439.84435620102
L16_153 V16 V153 2.6477707279856904e-12
C16_153 V16 V153 -3.561516439900029e-21

R16_154 V16 V154 -803.7180682229695
L16_154 V16 V154 -2.096856333009218e-12
C16_154 V16 V154 -1.424805279676112e-19

R16_155 V16 V155 -552.5211082512777
L16_155 V16 V155 -1.641319523702872e-12
C16_155 V16 V155 -1.540994405896606e-19

R16_156 V16 V156 1399.8882864548482
L16_156 V16 V156 -1.0199830452666728e-12
C16_156 V16 V156 -2.971717725445516e-19

R16_157 V16 V157 1151.475450984404
L16_157 V16 V157 7.023650467725885e-13
C16_157 V16 V157 5.751015816415581e-19

R16_158 V16 V158 1067.6672664833202
L16_158 V16 V158 -2.5595113919914016e-12
C16_158 V16 V158 -5.1596491987916946e-20

R16_159 V16 V159 515.1575130305562
L16_159 V16 V159 3.445671000194996e-12
C16_159 V16 V159 4.242417036147035e-20

R16_160 V16 V160 -463.76052258024754
L16_160 V16 V160 -1.5381310524628259e-12
C16_160 V16 V160 1.764983163774021e-19

R16_161 V16 V161 -1980.1585078318963
L16_161 V16 V161 -1.5236872478736831e-12
C16_161 V16 V161 -1.0415287861516522e-19

R16_162 V16 V162 9678.533954371205
L16_162 V16 V162 -2.618050243678485e-12
C16_162 V16 V162 -3.4287484021703285e-20

R16_163 V16 V163 6205.600800466384
L16_163 V16 V163 4.5469306037497844e-12
C16_163 V16 V163 9.04609007759164e-20

R16_164 V16 V164 250.7198842971996
L16_164 V16 V164 8.597783706904139e-13
C16_164 V16 V164 -9.169449141545898e-20

R16_165 V16 V165 987.3894216065711
L16_165 V16 V165 -3.83522609777719e-12
C16_165 V16 V165 -1.9455852989230195e-19

R16_166 V16 V166 2421.6049587312586
L16_166 V16 V166 1.4256311432791823e-12
C16_166 V16 V166 1.205852187210208e-19

R16_167 V16 V167 1046.9208069993956
L16_167 V16 V167 -7.396332144338919e-12
C16_167 V16 V167 -2.133952486200711e-20

R16_168 V16 V168 -305.4271660667277
L16_168 V16 V168 -2.6999444123481886e-12
C16_168 V16 V168 -1.3982093602344348e-20

R16_169 V16 V169 4052.0395651654408
L16_169 V16 V169 4.04600195503603e-12
C16_169 V16 V169 1.357989389254068e-19

R16_170 V16 V170 28507.37644978699
L16_170 V16 V170 -1.680383547619462e-12
C16_170 V16 V170 -1.6557092053993744e-19

R16_171 V16 V171 -935.7110146618412
L16_171 V16 V171 -1.3800695183797855e-12
C16_171 V16 V171 -1.6502395485447396e-19

R16_172 V16 V172 -1598.4412319670164
L16_172 V16 V172 -3.647964721904215e-12
C16_172 V16 V172 -3.603022992026502e-20

R16_173 V16 V173 -1901.0145418266295
L16_173 V16 V173 -3.2369204381328196e-12
C16_173 V16 V173 8.154710081978478e-20

R16_174 V16 V174 -967.1087850041486
L16_174 V16 V174 -2.8422811625287358e-12
C16_174 V16 V174 1.4628904336644203e-19

R16_175 V16 V175 15071.388483196082
L16_175 V16 V175 7.820521235746724e-12
C16_175 V16 V175 -2.284884839489055e-21

R16_176 V16 V176 571.8510945708884
L16_176 V16 V176 -2.6012039358187567e-12
C16_176 V16 V176 -2.325869973036779e-19

R16_177 V16 V177 1207.0570003297828
L16_177 V16 V177 6.474593553816228e-12
C16_177 V16 V177 -3.6254003238512287e-20

R16_178 V16 V178 1270.9148722657317
L16_178 V16 V178 1.3542780214750965e-12
C16_178 V16 V178 8.045333433021524e-20

R16_179 V16 V179 7052.877576924955
L16_179 V16 V179 1.5437374858509003e-12
C16_179 V16 V179 2.215987034069329e-19

R16_180 V16 V180 -2686.7837241020343
L16_180 V16 V180 8.904256906417557e-13
C16_180 V16 V180 3.302310119053969e-19

R16_181 V16 V181 -2800.2688435725727
L16_181 V16 V181 -1.803094403936794e-11
C16_181 V16 V181 -1.8926212411057252e-20

R16_182 V16 V182 -1321.9873322844776
L16_182 V16 V182 -1.7554780065022212e-12
C16_182 V16 V182 -1.3764676427044745e-19

R16_183 V16 V183 2105.2585010524276
L16_183 V16 V183 2.938284784008785e-12
C16_183 V16 V183 4.666382322810002e-20

R16_184 V16 V184 2337.192722163181
L16_184 V16 V184 6.467105402113443e-12
C16_184 V16 V184 -6.490294387117322e-20

R16_185 V16 V185 -4211.460921974944
L16_185 V16 V185 4.494039679884584e-10
C16_185 V16 V185 8.276139852400402e-21

R16_186 V16 V186 22288.897751153578
L16_186 V16 V186 2.7040824718239733e-10
C16_186 V16 V186 -2.8559968426316465e-20

R16_187 V16 V187 -2256.0211515277388
L16_187 V16 V187 -2.241404825181054e-12
C16_187 V16 V187 -2.251795813395955e-19

R16_188 V16 V188 -549.4568699293053
L16_188 V16 V188 -6.275511193297391e-13
C16_188 V16 V188 -1.812998970379488e-19

R16_189 V16 V189 2865.283488052405
L16_189 V16 V189 7.457992153026745e-12
C16_189 V16 V189 -3.605069657406428e-20

R16_190 V16 V190 1349.3956036215648
L16_190 V16 V190 4.997433242777082e-12
C16_190 V16 V190 1.372719691049836e-19

R16_191 V16 V191 -1818.081000902357
L16_191 V16 V191 -1.3771773174449989e-12
C16_191 V16 V191 -5.957569543965874e-20

R16_192 V16 V192 11308.796114733806
L16_192 V16 V192 1.1047288900188363e-12
C16_192 V16 V192 1.031349628329208e-19

R16_193 V16 V193 -2869.0334662533946
L16_193 V16 V193 1.162665592716487e-11
C16_193 V16 V193 1.1203647835548443e-19

R16_194 V16 V194 -8449.210282903969
L16_194 V16 V194 3.0823227876864268e-12
C16_194 V16 V194 1.5151351207077693e-19

R16_195 V16 V195 1059.2864931874299
L16_195 V16 V195 8.006600028600526e-13
C16_195 V16 V195 2.9390806316129505e-19

R16_196 V16 V196 632.0770957576534
L16_196 V16 V196 -2.6247539556514078e-12
C16_196 V16 V196 -1.4459328605849796e-19

R16_197 V16 V197 -3757.3301392566823
L16_197 V16 V197 -1.6623290549416894e-11
C16_197 V16 V197 -5.428011958023533e-20

R16_198 V16 V198 1796.788031524878
L16_198 V16 V198 -5.107752824184885e-12
C16_198 V16 V198 3.616860557520782e-21

R16_199 V16 V199 555.546655173683
L16_199 V16 V199 -6.509317254631615e-12
C16_199 V16 V199 1.2014616057893846e-20

R16_200 V16 V200 -561.6387424890428
L16_200 V16 V200 -1.3390075237919618e-11
C16_200 V16 V200 6.814266414121885e-20

R17_17 V17 0 -1382.3620918090242
L17_17 V17 0 -3.664882883708413e-13
C17_17 V17 0 -2.3072246727174757e-19

R17_18 V17 V18 -17315.8541097646
L17_18 V17 V18 -3.241075881586558e-12
C17_18 V17 V18 -2.0377510119340493e-19

R17_19 V17 V19 -11912.493086046738
L17_19 V17 V19 -3.3394939783219244e-12
C17_19 V17 V19 -2.1006292606755258e-19

R17_20 V17 V20 -7843.971591422908
L17_20 V17 V20 -2.328413193900024e-12
C17_20 V17 V20 -3.0074470021221588e-19

R17_21 V17 V21 -1749.2002575885374
L17_21 V17 V21 -2.2345496317897042e-12
C17_21 V17 V21 3.506814897879805e-19

R17_22 V17 V22 -15346.732991873085
L17_22 V17 V22 -4.503560763321473e-12
C17_22 V17 V22 3.606702873905449e-20

R17_23 V17 V23 -28988.24340403885
L17_23 V17 V23 -1.1897236140783584e-11
C17_23 V17 V23 1.0105014549558642e-19

R17_24 V17 V24 -14805.747765716273
L17_24 V17 V24 -9.72221059551701e-12
C17_24 V17 V24 1.2978273141652167e-19

R17_25 V17 V25 2034.6675191265304
L17_25 V17 V25 8.222978306529275e-13
C17_25 V17 V25 3.129092331047621e-19

R17_26 V17 V26 20067.970352343196
L17_26 V17 V26 2.5594086546811095e-12
C17_26 V17 V26 1.2464152461664236e-19

R17_27 V17 V27 31607.29279296491
L17_27 V17 V27 3.108440759198629e-12
C17_27 V17 V27 6.748760253592174e-20

R17_28 V17 V28 13647.472088899207
L17_28 V17 V28 2.038960109596194e-12
C17_28 V17 V28 1.2137140672676254e-19

R17_29 V17 V29 1217.9144422936406
L17_29 V17 V29 3.862693880602457e-12
C17_29 V17 V29 -1.4996462294609743e-19

R17_30 V17 V30 49196.85577753401
L17_30 V17 V30 1.1485018129070943e-11
C17_30 V17 V30 -1.1469551194385203e-20

R17_31 V17 V31 20192.285034815202
L17_31 V17 V31 2.146668577389437e-11
C17_31 V17 V31 -1.3361309924172646e-20

R17_32 V17 V32 8371.162795970999
L17_32 V17 V32 1.59812383235502e-11
C17_32 V17 V32 1.7871281187031304e-20

R17_33 V17 V33 29342.030163929383
L17_33 V17 V33 2.3778783218155196e-12
C17_33 V17 V33 2.097340483681374e-19

R17_34 V17 V34 -13658.158240710352
L17_34 V17 V34 -2.896490789570067e-11
C17_34 V17 V34 -8.643622763147182e-20

R17_35 V17 V35 -12217.090006076865
L17_35 V17 V35 -9.697808786980815e-11
C17_35 V17 V35 2.4012845515548096e-21

R17_36 V17 V36 -11454.03612621011
L17_36 V17 V36 -1.3650895763868366e-11
C17_36 V17 V36 4.064295580974453e-20

R17_37 V17 V37 -2135.322922239506
L17_37 V17 V37 -1.127144024569723e-12
C17_37 V17 V37 -4.150634966168723e-19

R17_38 V17 V38 -19786.622300091658
L17_38 V17 V38 -5.935399929060846e-12
C17_38 V17 V38 -1.4283478727978382e-20

R17_39 V17 V39 -12179.4580609642
L17_39 V17 V39 -4.184986358769281e-12
C17_39 V17 V39 -1.303991423931396e-19

R17_40 V17 V40 -7484.373533237382
L17_40 V17 V40 -2.819283671569171e-12
C17_40 V17 V40 -1.852946881225367e-19

R17_41 V17 V41 -18022.50035925305
L17_41 V17 V41 1.603283237997439e-11
C17_41 V17 V41 1.4334077570540392e-19

R17_42 V17 V42 -99217.3160167345
L17_42 V17 V42 1.6361971595385576e-11
C17_42 V17 V42 3.545893432056233e-20

R17_43 V17 V43 -79891.04441706097
L17_43 V17 V43 2.988227812126643e-11
C17_43 V17 V43 8.312065639869578e-20

R17_44 V17 V44 84913.41958430233
L17_44 V17 V44 1.2306791003406094e-11
C17_44 V17 V44 1.4992788918207576e-19

R17_45 V17 V45 1809.9115634764962
L17_45 V17 V45 1.9017661249817023e-12
C17_45 V17 V45 2.265758828489186e-19

R17_46 V17 V46 -83550.06483013454
L17_46 V17 V46 -1.1072559916733705e-11
C17_46 V17 V46 -8.15663020880265e-20

R17_47 V17 V47 -853539.6041219577
L17_47 V17 V47 2.042236901622458e-11
C17_47 V17 V47 1.8557113987032645e-20

R17_48 V17 V48 15619.090866859984
L17_48 V17 V48 6.1334428750329025e-12
C17_48 V17 V48 6.035272220608108e-20

R17_49 V17 V49 3162.2563418246623
L17_49 V17 V49 -6.251104699997084e-12
C17_49 V17 V49 -2.24993262436563e-19

R17_50 V17 V50 -15977.831938421383
L17_50 V17 V50 9.826912420476828e-12
C17_50 V17 V50 7.183043503130039e-20

R17_51 V17 V51 -58696.82217634558
L17_51 V17 V51 1.6659811822586462e-11
C17_51 V17 V51 -4.108847045074422e-21

R17_52 V17 V52 -42106.95613455819
L17_52 V17 V52 -3.094468598916784e-11
C17_52 V17 V52 -1.2794723849410278e-20

R17_53 V17 V53 27704.820849265212
L17_53 V17 V53 1.93645265245334e-12
C17_53 V17 V53 1.1051776418735685e-19

R17_54 V17 V54 44406.0170960909
L17_54 V17 V54 4.1278483991497936e-11
C17_54 V17 V54 -4.4964763434092966e-20

R17_55 V17 V55 39869.29846896676
L17_55 V17 V55 8.516361782163626e-12
C17_55 V17 V55 5.8242814228818985e-21

R17_56 V17 V56 -92677.95965896448
L17_56 V17 V56 4.376009383399253e-11
C17_56 V17 V56 -2.1894486273961895e-21

R17_57 V17 V57 -6273.052330054423
L17_57 V17 V57 -1.968145997078169e-12
C17_57 V17 V57 -1.7213058623046552e-19

R17_58 V17 V58 -15832.466979148077
L17_58 V17 V58 5.614916896743407e-11
C17_58 V17 V58 1.9951150339924814e-20

R17_59 V17 V59 -8902.150510735559
L17_59 V17 V59 -8.503703479760437e-12
C17_59 V17 V59 -4.8578968043397326e-20

R17_60 V17 V60 -6910.778812877557
L17_60 V17 V60 -5.799925909702521e-12
C17_60 V17 V60 -3.196991695435316e-20

R17_61 V17 V61 179766.35987838183
L17_61 V17 V61 6.34588498300835e-12
C17_61 V17 V61 9.185983850446602e-20

R17_62 V17 V62 559330.8731583292
L17_62 V17 V62 -1.59258767137778e-10
C17_62 V17 V62 -2.084195384222745e-20

R17_63 V17 V63 340742.4613620807
L17_63 V17 V63 -1.010558208481961e-11
C17_63 V17 V63 -1.0665410391076223e-20

R17_64 V17 V64 20165.50265662789
L17_64 V17 V64 -2.5681929897754025e-11
C17_64 V17 V64 1.4071748523716193e-20

R17_65 V17 V65 2507.555189392573
L17_65 V17 V65 2.4305184152904304e-11
C17_65 V17 V65 4.099827192728863e-20

R17_66 V17 V66 -15398.33580258399
L17_66 V17 V66 -4.936144322715843e-12
C17_66 V17 V66 -8.347489405439089e-20

R17_67 V17 V67 -54613.66841343519
L17_67 V17 V67 -7.032145932726376e-12
C17_67 V17 V67 -4.1108222873086136e-20

R17_68 V17 V68 24230.134648768202
L17_68 V17 V68 -1.429456715872776e-11
C17_68 V17 V68 -1.0069285707834115e-20

R17_69 V17 V69 8066.017184400607
L17_69 V17 V69 3.948082687264529e-12
C17_69 V17 V69 1.2979820911814916e-20

R17_70 V17 V70 -20936.954744272414
L17_70 V17 V70 6.407817362240509e-12
C17_70 V17 V70 8.927426196815469e-20

R17_71 V17 V71 -38923.2038177692
L17_71 V17 V71 4.543816890246599e-12
C17_71 V17 V71 6.060552376452755e-20

R17_72 V17 V72 -16239.097078801356
L17_72 V17 V72 4.700215088287097e-12
C17_72 V17 V72 4.0864620941915595e-20

R17_73 V17 V73 -6125.791182033996
L17_73 V17 V73 2.2889031673038642e-12
C17_73 V17 V73 1.5568059736037002e-19

R17_74 V17 V74 28902.414419589495
L17_74 V17 V74 4.222215300129269e-12
C17_74 V17 V74 5.0229764649404866e-20

R17_75 V17 V75 13254.700111580843
L17_75 V17 V75 5.791998875450603e-12
C17_75 V17 V75 8.505588585265104e-20

R17_76 V17 V76 48862.65866413223
L17_76 V17 V76 1.1822447751599918e-11
C17_76 V17 V76 9.356317398291618e-20

R17_77 V17 V77 -6421.0012368954485
L17_77 V17 V77 -1.5827740209062844e-12
C17_77 V17 V77 -3.2047113258775793e-19

R17_78 V17 V78 8950.683052219307
L17_78 V17 V78 -9.41553276801304e-12
C17_78 V17 V78 2.7048333035344774e-20

R17_79 V17 V79 -166636.42979462454
L17_79 V17 V79 -3.757790059291637e-12
C17_79 V17 V79 -1.1723105040087292e-19

R17_80 V17 V80 33645.848075199625
L17_80 V17 V80 -3.1994496936805977e-12
C17_80 V17 V80 -1.434586652504875e-19

R17_81 V17 V81 1275.4871457650859
L17_81 V17 V81 4.987774406718821e-12
C17_81 V17 V81 7.750268831743293e-20

R17_82 V17 V82 -5876.354299533418
L17_82 V17 V82 -3.4603970783792856e-12
C17_82 V17 V82 -1.915784398056562e-19

R17_83 V17 V83 -4047.1933580136774
L17_83 V17 V83 -4.22184016945587e-12
C17_83 V17 V83 -1.1580560337381765e-19

R17_84 V17 V84 -5833.784055447238
L17_84 V17 V84 -3.0475371606338613e-12
C17_84 V17 V84 -1.1645399438780792e-19

R17_85 V17 V85 15866.20794011015
L17_85 V17 V85 2.238591878759256e-12
C17_85 V17 V85 2.984253446201149e-19

R17_86 V17 V86 -2775.5152525404374
L17_86 V17 V86 6.444952389634608e-12
C17_86 V17 V86 3.9810338094524205e-20

R17_87 V17 V87 -62472.48092165932
L17_87 V17 V87 4.8878636308889934e-12
C17_87 V17 V87 1.3127293192356575e-19

R17_88 V17 V88 -28761.680133169215
L17_88 V17 V88 2.8123966672581704e-12
C17_88 V17 V88 2.0100354238633444e-19

R17_89 V17 V89 -4564.294569202963
L17_89 V17 V89 2.899543496717217e-12
C17_89 V17 V89 -1.8649945009088072e-20

R17_90 V17 V90 3002.2712515148296
L17_90 V17 V90 4.82631561457994e-12
C17_90 V17 V90 1.8959543117309812e-19

R17_91 V17 V91 4438.348072008937
L17_91 V17 V91 7.359476776810747e-12
C17_91 V17 V91 3.403879513643509e-20

R17_92 V17 V92 9446.419415601797
L17_92 V17 V92 2.1121277066795162e-11
C17_92 V17 V92 -2.149144719905904e-20

R17_93 V17 V93 2600.050480349194
L17_93 V17 V93 -1.6352728399236493e-12
C17_93 V17 V93 -2.7604727442463095e-19

R17_94 V17 V94 7721.258272145161
L17_94 V17 V94 -6.785796827026896e-12
C17_94 V17 V94 -1.35600868860596e-19

R17_95 V17 V95 71047.33563235994
L17_95 V17 V95 -5.153366571719093e-12
C17_95 V17 V95 -1.076638430380453e-19

R17_96 V17 V96 22873.41654181438
L17_96 V17 V96 -3.5530875910802404e-12
C17_96 V17 V96 -1.4332277553431622e-19

R17_97 V17 V97 11164.670740748572
L17_97 V17 V97 9.371952169294348e-12
C17_97 V17 V97 -3.960119523965059e-20

R17_98 V17 V98 -2145.9506240214723
L17_98 V17 V98 -1.7816417239600425e-11
C17_98 V17 V98 -6.922473821455319e-20

R17_99 V17 V99 -2269.6822012377356
L17_99 V17 V99 -2.499642527045739e-11
C17_99 V17 V99 -9.450681460828085e-21

R17_100 V17 V100 -3077.070027660351
L17_100 V17 V100 -1.1140951832116321e-11
C17_100 V17 V100 4.294762734469269e-20

R17_101 V17 V101 -6937.83819035965
L17_101 V17 V101 1.929329967977553e-12
C17_101 V17 V101 2.258368826004789e-19

R17_102 V17 V102 25720.148698152912
L17_102 V17 V102 1.5768092769259182e-11
C17_102 V17 V102 5.969408155605115e-20

R17_103 V17 V103 19619.671980129835
L17_103 V17 V103 2.0868823472679388e-11
C17_103 V17 V103 2.159820705509313e-20

R17_104 V17 V104 194898.06115487497
L17_104 V17 V104 3.494541430060518e-11
C17_104 V17 V104 1.5983885248579823e-20

R17_105 V17 V105 1083.439227741107
L17_105 V17 V105 -5.009748295355262e-10
C17_105 V17 V105 1.0664982135100035e-19

R17_106 V17 V106 -10104.380305704768
L17_106 V17 V106 8.597343524739706e-11
C17_106 V17 V106 7.183541897412588e-20

R17_107 V17 V107 15297.775823493868
L17_107 V17 V107 8.979432207342932e-11
C17_107 V17 V107 1.6519787120132935e-20

R17_108 V17 V108 29749.82462910896
L17_108 V17 V108 4.871237924141293e-12
C17_108 V17 V108 7.757863423459221e-20

R17_109 V17 V109 -3053.4314910246126
L17_109 V17 V109 8.234855404817476e-12
C17_109 V17 V109 -1.377407931220798e-19

R17_110 V17 V110 15614.497987234723
L17_110 V17 V110 -1.977380526480865e-11
C17_110 V17 V110 -3.457190698306669e-20

R17_111 V17 V111 -33670.91582500962
L17_111 V17 V111 1.7456757248653703e-11
C17_111 V17 V111 1.9556759380802687e-20

R17_112 V17 V112 -15128.012344832088
L17_112 V17 V112 -8.898795883819291e-12
C17_112 V17 V112 -8.218925025241148e-20

R17_113 V17 V113 -12395.937450486756
L17_113 V17 V113 -3.938439940782535e-12
C17_113 V17 V113 -2.3964314954093606e-19

R17_114 V17 V114 -59964.77172402639
L17_114 V17 V114 -9.404703705669873e-12
C17_114 V17 V114 -1.1933815813763992e-19

R17_115 V17 V115 -11685.948765369576
L17_115 V17 V115 -1.1690409002853181e-11
C17_115 V17 V115 -5.149901878531182e-20

R17_116 V17 V116 -35270.57847215709
L17_116 V17 V116 -6.697537932784395e-12
C17_116 V17 V116 -7.984822137991317e-20

R17_117 V17 V117 2560.4827104801316
L17_117 V17 V117 -3.5598886794509673e-12
C17_117 V17 V117 1.2205309802324714e-19

R17_118 V17 V118 781693.9334050546
L17_118 V17 V118 2.7765367471730288e-11
C17_118 V17 V118 1.2433931677788662e-19

R17_119 V17 V119 -18303.14184033137
L17_119 V17 V119 1.0909085113977746e-11
C17_119 V17 V119 9.922569356886389e-20

R17_120 V17 V120 -7428.7186697259685
L17_120 V17 V120 6.251196275384456e-12
C17_120 V17 V120 1.5614457404082472e-19

R17_121 V17 V121 17238.701954543005
L17_121 V17 V121 1.5159295616589146e-12
C17_121 V17 V121 1.9576765865355412e-19

R17_122 V17 V122 -6567.565538471691
L17_122 V17 V122 9.915355108397822e-12
C17_122 V17 V122 2.4835858186751013e-20

R17_123 V17 V123 79178.54414636012
L17_123 V17 V123 -9.673549747636064e-12
C17_123 V17 V123 -6.62796852520085e-20

R17_124 V17 V124 13206.714478853537
L17_124 V17 V124 -9.291831647914755e-12
C17_124 V17 V124 -1.0247274674840351e-19

R17_125 V17 V125 1801.474752226117
L17_125 V17 V125 4.043010354994837e-12
C17_125 V17 V125 -8.826529745761517e-21

R17_126 V17 V126 11459.570143434037
L17_126 V17 V126 7.511048004288986e-10
C17_126 V17 V126 -4.52856728571526e-21

R17_127 V17 V127 16115.76353377773
L17_127 V17 V127 -3.4590407590812934e-11
C17_127 V17 V127 -1.105294705796062e-20

R17_128 V17 V128 7923.456436034123
L17_128 V17 V128 2.8651468180937888e-11
C17_128 V17 V128 -8.161140519932958e-21

R17_129 V17 V129 -3663.3210466069486
L17_129 V17 V129 -5.969764051944717e-12
C17_129 V17 V129 4.882274067261565e-21

R17_130 V17 V130 20437.562485997358
L17_130 V17 V130 -7.27036588175587e-12
C17_130 V17 V130 -4.0371261585012485e-20

R17_131 V17 V131 -15083.090715109976
L17_131 V17 V131 1.6243540403466842e-11
C17_131 V17 V131 1.0232172861217944e-20

R17_132 V17 V132 -4023.9016498713795
L17_132 V17 V132 2.14046931495875e-11
C17_132 V17 V132 3.4695683042825025e-20

R17_133 V17 V133 -2119.37442759602
L17_133 V17 V133 -2.749637051768549e-12
C17_133 V17 V133 -2.9159849118312296e-19

R17_134 V17 V134 -3147.916646559147
L17_134 V17 V134 -1.3065273746932726e-11
C17_134 V17 V134 -1.552636815469445e-20

R17_135 V17 V135 114282.22755460948
L17_135 V17 V135 -7.751516462727659e-12
C17_135 V17 V135 -3.645969622938916e-20

R17_136 V17 V136 34991.31392647364
L17_136 V17 V136 -5.360895769153034e-12
C17_136 V17 V136 -1.2275757595133163e-19

R17_137 V17 V137 1395.2164089670944
L17_137 V17 V137 -2.6910020706895494e-12
C17_137 V17 V137 -5.6255609466817285e-21

R17_138 V17 V138 2265.939160904687
L17_138 V17 V138 2.018115425265885e-11
C17_138 V17 V138 4.477623060312034e-20

R17_139 V17 V139 -13675.588590407571
L17_139 V17 V139 3.369595452199294e-12
C17_139 V17 V139 1.1822981917180498e-19

R17_140 V17 V140 197127.3580996365
L17_140 V17 V140 4.200662335419468e-12
C17_140 V17 V140 1.5924304810722487e-19

R17_141 V17 V141 -5189.79569946041
L17_141 V17 V141 1.233210370597958e-12
C17_141 V17 V141 3.207215963660457e-19

R17_142 V17 V142 -5934.438953454837
L17_142 V17 V142 5.850361117216575e-12
C17_142 V17 V142 2.7708918273073776e-20

R17_143 V17 V143 -9003.446441134725
L17_143 V17 V143 -3.765372169747372e-12
C17_143 V17 V143 -1.083073268098068e-19

R17_144 V17 V144 -5452.686481977983
L17_144 V17 V144 -1.696441966675597e-11
C17_144 V17 V144 -1.015470734163044e-20

R17_145 V17 V145 2035.1041482403832
L17_145 V17 V145 2.8348214826224514e-12
C17_145 V17 V145 -5.616193043154686e-20

R17_146 V17 V146 -2591.3548143706057
L17_146 V17 V146 -9.40324051857525e-12
C17_146 V17 V146 -6.454350369278177e-20

R17_147 V17 V147 4556.258622420687
L17_147 V17 V147 -3.1261381847504025e-10
C17_147 V17 V147 -8.034114871756296e-21

R17_148 V17 V148 2956.300286505959
L17_148 V17 V148 3.284223631206153e-11
C17_148 V17 V148 -2.8030487601359285e-20

R17_149 V17 V149 -706.8061152453951
L17_149 V17 V149 -2.483637520317437e-12
C17_149 V17 V149 6.279907198356393e-20

R17_150 V17 V150 3305.819797097402
L17_150 V17 V150 -1.0061942334345579e-10
C17_150 V17 V150 -2.7436086055779977e-20

R17_151 V17 V151 7449.612459717541
L17_151 V17 V151 2.3772206373714007e-12
C17_151 V17 V151 8.819772164201636e-20

R17_152 V17 V152 -6610.167507145001
L17_152 V17 V152 9.809190201240709e-12
C17_152 V17 V152 -1.9046174077158867e-20

R17_153 V17 V153 1016.368880400691
L17_153 V17 V153 -3.4845376098036443e-12
C17_153 V17 V153 -1.169684446454503e-19

R17_154 V17 V154 -77793.03752871597
L17_154 V17 V154 -6.120992103490616e-10
C17_154 V17 V154 1.536675542547901e-20

R17_155 V17 V155 -3214.0762777455016
L17_155 V17 V155 2.5814939051919707e-11
C17_155 V17 V155 3.388096316589447e-20

R17_156 V17 V156 -9653.160055368986
L17_156 V17 V156 -3.787897944338023e-10
C17_156 V17 V156 4.766478157570358e-20

R17_157 V17 V157 2129.11141679908
L17_157 V17 V157 -1.3679598608296462e-11
C17_157 V17 V157 -3.3781885377236474e-19

R17_158 V17 V158 -37963.06687487754
L17_158 V17 V158 4.1125465010308264e-11
C17_158 V17 V158 4.010385419747549e-20

R17_159 V17 V159 35096.8024652239
L17_159 V17 V159 -2.2597091728788345e-12
C17_159 V17 V159 -7.024207557469059e-20

R17_160 V17 V160 -42285.60908345705
L17_160 V17 V160 -3.236478143796666e-12
C17_160 V17 V160 -2.0783620233639968e-20

R17_161 V17 V161 2181.977991773713
L17_161 V17 V161 5.454940919414346e-12
C17_161 V17 V161 3.189474366021738e-19

R17_162 V17 V162 -4078.2332422372324
L17_162 V17 V162 -1.250212688575538e-11
C17_162 V17 V162 -8.191711848905921e-20

R17_163 V17 V163 -3520.0587751433177
L17_163 V17 V163 -3.817231437721138e-12
C17_163 V17 V163 -9.915014481632063e-20

R17_164 V17 V164 -17285.22099945731
L17_164 V17 V164 -1.0545878196997577e-10
C17_164 V17 V164 7.639235193588524e-21

R17_165 V17 V165 19962.13218186812
L17_165 V17 V165 1.2244372259273504e-12
C17_165 V17 V165 2.338231573256159e-19

R17_166 V17 V166 -2531.971762629989
L17_166 V17 V166 2.5447629253877743e-12
C17_166 V17 V166 5.1367786494045306e-20

R17_167 V17 V167 13721.55993257711
L17_167 V17 V167 2.025831421870117e-12
C17_167 V17 V167 1.2298069674769333e-19

R17_168 V17 V168 -3392.7454536559558
L17_168 V17 V168 2.5964007994177604e-12
C17_168 V17 V168 1.0816931405277835e-19

R17_169 V17 V169 11262.460890525328
L17_169 V17 V169 -4.303691566857531e-12
C17_169 V17 V169 -1.9395501375401991e-19

R17_170 V17 V170 1543.1017090546466
L17_170 V17 V170 -6.427748280720369e-12
C17_170 V17 V170 6.226294867057298e-20

R17_171 V17 V171 3107.5374568361544
L17_171 V17 V171 5.487574580731664e-12
C17_171 V17 V171 8.269412846319234e-20

R17_172 V17 V172 4890.480066651188
L17_172 V17 V172 -9.529653753992265e-12
C17_172 V17 V172 -8.261860838790966e-25

R17_173 V17 V173 1768.1003930076074
L17_173 V17 V173 -1.4890359691380666e-12
C17_173 V17 V173 -2.191883434306611e-19

R17_174 V17 V174 -2905.49708192284
L17_174 V17 V174 -1.7474927746468608e-12
C17_174 V17 V174 -1.845165742160099e-19

R17_175 V17 V175 -2660.688308671681
L17_175 V17 V175 -2.1842482109474037e-12
C17_175 V17 V175 -1.4167508318496483e-19

R17_176 V17 V176 -4358.377953398823
L17_176 V17 V176 -1.7364859792520827e-12
C17_176 V17 V176 -1.6638572114010383e-19

R17_177 V17 V177 -1790.6346148127018
L17_177 V17 V177 4.6784766130538e-12
C17_177 V17 V177 1.5996369383277536e-19

R17_178 V17 V178 10405.925495845777
L17_178 V17 V178 6.625333062903838e-12
C17_178 V17 V178 -2.3424849128152995e-20

R17_179 V17 V179 16520.920637043742
L17_179 V17 V179 -2.3285282224593105e-11
C17_179 V17 V179 -7.225689136229367e-20

R17_180 V17 V180 4356.23266579262
L17_180 V17 V180 4.1244310404988175e-12
C17_180 V17 V180 -1.0635122845307154e-21

R17_181 V17 V181 -6438.5154284460605
L17_181 V17 V181 -6.255521900069484e-12
C17_181 V17 V181 2.000509063395287e-19

R17_182 V17 V182 8424.738864554654
L17_182 V17 V182 3.807096172844582e-12
C17_182 V17 V182 8.772041753058711e-20

R17_183 V17 V183 51929.2447734931
L17_183 V17 V183 -1.3081691686096429e-11
C17_183 V17 V183 3.6960008606605947e-20

R17_184 V17 V184 -12915.635126153977
L17_184 V17 V184 7.679566446853222e-12
C17_184 V17 V184 7.89909818795358e-20

R17_185 V17 V185 769.4087578865257
L17_185 V17 V185 1.7022005203163134e-12
C17_185 V17 V185 -1.9098315105196231e-19

R17_186 V17 V186 -1467.559067479634
L17_186 V17 V186 2.3958237534805134e-12
C17_186 V17 V186 1.7727009134422783e-19

R17_187 V17 V187 -7185.473782862091
L17_187 V17 V187 1.947624399915017e-12
C17_187 V17 V187 1.2841609155101707e-19

R17_188 V17 V188 -9847.454549159025
L17_188 V17 V188 1.8646612549017295e-12
C17_188 V17 V188 1.1647822781502018e-19

R17_189 V17 V189 -889.4142787708513
L17_189 V17 V189 1.842510291865178e-11
C17_189 V17 V189 2.088442075075713e-20

R17_190 V17 V190 6040.067897668857
L17_190 V17 V190 -3.1769741858442376e-12
C17_190 V17 V190 -1.0869974921340673e-19

R17_191 V17 V191 1720.0593026961346
L17_191 V17 V191 6.043613509601856e-12
C17_191 V17 V191 -4.9424280052847297e-20

R17_192 V17 V192 2116.4733067659226
L17_192 V17 V192 -3.4514936241392664e-12
C17_192 V17 V192 -1.9696148601505994e-19

R17_193 V17 V193 -1603.6582882031228
L17_193 V17 V193 -1.1212074976436605e-12
C17_193 V17 V193 -1.7151988887247858e-19

R17_194 V17 V194 1179.9841378486894
L17_194 V17 V194 -2.2849539658216776e-12
C17_194 V17 V194 -1.6327514208885034e-19

R17_195 V17 V195 -23145.666352847948
L17_195 V17 V195 -3.4717914332121943e-12
C17_195 V17 V195 -2.878070771913063e-20

R17_196 V17 V196 19756.860602522327
L17_196 V17 V196 -2.836057625803504e-12
C17_196 V17 V196 2.1669467933182484e-20

R17_197 V17 V197 969.811880617678
L17_197 V17 V197 4.807986059897501e-12
C17_197 V17 V197 1.924046701100097e-19

R17_198 V17 V198 -1418.7717422662545
L17_198 V17 V198 6.057928555926078e-12
C17_198 V17 V198 1.5613480441929936e-20

R17_199 V17 V199 -954.617543024966
L17_199 V17 V199 -4.8331233152973574e-12
C17_199 V17 V199 -9.008429759086692e-20

R17_200 V17 V200 -1192.3081354153655
L17_200 V17 V200 5.389772015239951e-12
C17_200 V17 V200 1.1400113765942765e-19

R18_18 V18 0 -1048.9709848926263
L18_18 V18 0 -7.933387871540071e-13
C18_18 V18 0 1.0984228326119438e-19

R18_19 V18 V19 -61171.0380310442
L18_19 V18 V19 -3.198922256019652e-12
C18_19 V18 V19 -2.528851975296677e-19

R18_20 V18 V20 -21826.56944790925
L18_20 V18 V20 -2.439946867429371e-12
C18_20 V18 V20 -3.461023907874015e-19

R18_21 V18 V21 9872.525396261113
L18_21 V18 V21 -4.442089400276349e-12
C18_21 V18 V21 5.804153393781182e-20

R18_22 V18 V22 -3884.098903669047
L18_22 V18 V22 2.3504251513252566e-12
C18_22 V18 V22 5.029695736157842e-19

R18_23 V18 V23 30349.991561866875
L18_23 V18 V23 8.923024112143204e-12
C18_23 V18 V23 1.2605668655702537e-19

R18_24 V18 V24 41989.42544816114
L18_24 V18 V24 6.552384185488055e-12
C18_24 V18 V24 1.7078885464946155e-19

R18_25 V18 V25 -31841.487236871075
L18_25 V18 V25 1.916929047858581e-12
C18_25 V18 V25 2.46545619337109e-19

R18_26 V18 V26 5270.962711529448
L18_26 V18 V26 9.010352976530927e-13
C18_26 V18 V26 6.370461548247894e-19

R18_27 V18 V27 112349.1822276584
L18_27 V18 V27 2.649355307465582e-12
C18_27 V18 V27 2.1789477876423694e-19

R18_28 V18 V28 53214.96578069055
L18_28 V18 V28 1.956229767184933e-12
C18_28 V18 V28 2.67341289269941e-19

R18_29 V18 V29 -32505.914369873746
L18_29 V18 V29 1.0593482336305075e-11
C18_29 V18 V29 -7.392687913330174e-20

R18_30 V18 V30 1810.2320985323142
L18_30 V18 V30 -1.4390654521847507e-12
C18_30 V18 V30 -5.282285229608787e-19

R18_31 V18 V31 -69201.94094209686
L18_31 V18 V31 -5.3333955297828614e-12
C18_31 V18 V31 -1.4206214718222968e-19

R18_32 V18 V32 22735.864494159832
L18_32 V18 V32 -4.4350170912473125e-12
C18_32 V18 V32 -1.3657850354723975e-19

R18_33 V18 V33 -12561.201704686831
L18_33 V18 V33 -1.0330206282873105e-11
C18_33 V18 V33 -4.487627980785918e-20

R18_34 V18 V34 -4335.202592502223
L18_34 V18 V34 -9.910421932377718e-12
C18_34 V18 V34 -7.516048572385523e-20

R18_35 V18 V35 -17405.713991065044
L18_35 V18 V35 -4.656283016708269e-12
C18_35 V18 V35 -1.04597562195999e-19

R18_36 V18 V36 -16082.721670731227
L18_36 V18 V36 -3.2226286947433727e-12
C18_36 V18 V36 -1.1686974842541839e-19

R18_37 V18 V37 -47199.73879825412
L18_37 V18 V37 -5.113420315174907e-12
C18_37 V18 V37 -9.38611931028406e-20

R18_38 V18 V38 -3841.34228448286
L18_38 V18 V38 3.381548940566769e-12
C18_38 V18 V38 2.972563799014696e-19

R18_39 V18 V39 77964.71479109405
L18_39 V18 V39 4.730115075524531e-12
C18_39 V18 V39 1.2542341229778885e-19

R18_40 V18 V40 -95195.53609931323
L18_40 V18 V40 3.976344219011452e-12
C18_40 V18 V40 1.3109495833458058e-19

R18_41 V18 V41 17848.1349558519
L18_41 V18 V41 -7.78059518676901e-11
C18_41 V18 V41 -2.8392880188111038e-21

R18_42 V18 V42 -5637.088858406703
L18_42 V18 V42 -1.8693440723773634e-11
C18_42 V18 V42 -7.669353400884282e-20

R18_43 V18 V43 54348.56367358448
L18_43 V18 V43 -5.8715973029873606e-12
C18_43 V18 V43 -8.445261206808525e-20

R18_44 V18 V44 20841.211440017465
L18_44 V18 V44 -5.882288820230969e-12
C18_44 V18 V44 -6.036047607603634e-20

R18_45 V18 V45 25800.045878332585
L18_45 V18 V45 2.809145182602048e-12
C18_45 V18 V45 1.8718771021128706e-19

R18_46 V18 V46 2889.3541458358345
L18_46 V18 V46 -1.9900798696684307e-12
C18_46 V18 V46 -3.296920519618302e-19

R18_47 V18 V47 -28420.032741341958
L18_47 V18 V47 -1.1294755428458608e-10
C18_47 V18 V47 -2.4488769485619246e-20

R18_48 V18 V48 68903.55546880928
L18_48 V18 V48 2.1558024084509386e-11
C18_48 V18 V48 -3.691989971608111e-21

R18_49 V18 V49 -13523.212429295707
L18_49 V18 V49 -7.362009782794085e-11
C18_49 V18 V49 -5.3329523593742795e-21

R18_50 V18 V50 4369.808785887581
L18_50 V18 V50 2.7657256895845894e-12
C18_50 V18 V50 3.4812249600633403e-19

R18_51 V18 V51 -63339.18099263648
L18_51 V18 V51 3.124863332602353e-12
C18_51 V18 V51 2.5251975075213312e-19

R18_52 V18 V52 152519.20818912395
L18_52 V18 V52 2.746362617241213e-12
C18_52 V18 V52 3.0877939111763893e-19

R18_53 V18 V53 -24785.802482598727
L18_53 V18 V53 -3.740629314326225e-12
C18_53 V18 V53 -2.29342351616222e-19

R18_54 V18 V54 -4151.179049452194
L18_54 V18 V54 5.068668826312651e-12
C18_54 V18 V54 3.8208471628219804e-20

R18_55 V18 V55 -17994.284394494996
L18_55 V18 V55 -3.3393482264747145e-12
C18_55 V18 V55 -2.2341812318596477e-19

R18_56 V18 V56 -9577.640971239554
L18_56 V18 V56 -2.475173676648315e-12
C18_56 V18 V56 -2.471512536754579e-19

R18_57 V18 V57 -34834.83880401522
L18_57 V18 V57 1.146893565027885e-11
C18_57 V18 V57 1.263972562897362e-20

R18_58 V18 V58 24238.809783517714
L18_58 V18 V58 -1.7416166647153101e-12
C18_58 V18 V58 -4.010596959127929e-19

R18_59 V18 V59 24474.72855006868
L18_59 V18 V59 -6.388843008037271e-12
C18_59 V18 V59 -1.6199281262975703e-19

R18_60 V18 V60 20791.299332371258
L18_60 V18 V60 -4.078912402259621e-12
C18_60 V18 V60 -2.154866732692152e-19

R18_61 V18 V61 15308.021589843029
L18_61 V18 V61 4.039830769312549e-12
C18_61 V18 V61 2.101699692700337e-19

R18_62 V18 V62 -6082.6982862736
L18_62 V18 V62 3.9446118051207685e-12
C18_62 V18 V62 1.7659632803883635e-19

R18_63 V18 V63 96268.11000695574
L18_63 V18 V63 3.164490139378936e-12
C18_63 V18 V63 2.5904140238647744e-19

R18_64 V18 V64 15702.059524330567
L18_64 V18 V64 1.9417877083085808e-12
C18_64 V18 V64 3.877731497688271e-19

R18_65 V18 V65 87137.1033626568
L18_65 V18 V65 -3.9911816088289535e-12
C18_65 V18 V65 -1.5847069614468278e-19

R18_66 V18 V66 3827.8983162547115
L18_66 V18 V66 5.140609116715543e-12
C18_66 V18 V66 8.486056157515132e-20

R18_67 V18 V67 -27035.84635102022
L18_67 V18 V67 -6.302500490163594e-12
C18_67 V18 V67 -7.636406999714226e-20

R18_68 V18 V68 196369.4286348464
L18_68 V18 V68 -9.914230236160605e-12
C18_68 V18 V68 -7.106876291354049e-20

R18_69 V18 V69 -9074.817557816097
L18_69 V18 V69 1.6711424363794458e-11
C18_69 V18 V69 5.199719783099652e-21

R18_70 V18 V70 4853.749744912518
L18_70 V18 V70 -4.784919088211924e-12
C18_70 V18 V70 -7.15809353116608e-20

R18_71 V18 V71 -207447.97844248128
L18_71 V18 V71 -1.2112275232284091e-11
C18_71 V18 V71 -1.0442819931031204e-19

R18_72 V18 V72 -29515.77191876217
L18_72 V18 V72 -3.1967775208216892e-12
C18_72 V18 V72 -2.5271284056371974e-19

R18_73 V18 V73 12995.489394801676
L18_73 V18 V73 3.9072917887643175e-12
C18_73 V18 V73 1.125235080746524e-19

R18_74 V18 V74 -2958.350096888496
L18_74 V18 V74 2.4172722897717864e-11
C18_74 V18 V74 -1.9794438205512558e-20

R18_75 V18 V75 11358.29165077204
L18_75 V18 V75 4.865140716484933e-12
C18_75 V18 V75 1.4073605610012887e-19

R18_76 V18 V76 36324.5251700623
L18_76 V18 V76 3.914599549960506e-12
C18_76 V18 V76 2.5004642855993024e-19

R18_77 V18 V77 -37288.54169058745
L18_77 V18 V77 -3.722631114692954e-12
C18_77 V18 V77 -2.0607956344976137e-19

R18_78 V18 V78 13732.67452197766
L18_78 V18 V78 -1.2560863711757863e-10
C18_78 V18 V78 -1.334770594267725e-19

R18_79 V18 V79 -26200.483003043744
L18_79 V18 V79 8.015814265183816e-11
C18_79 V18 V79 -2.5550305168795636e-20

R18_80 V18 V80 91226.25802927832
L18_80 V18 V80 1.090661687089373e-11
C18_80 V18 V80 -3.42621896069739e-20

R18_81 V18 V81 20688.905501443696
L18_81 V18 V81 5.804812520055818e-12
C18_81 V18 V81 8.972603014285531e-20

R18_82 V18 V82 13083.335114746
L18_82 V18 V82 1.0004313699416514e-11
C18_82 V18 V82 1.0006979346830453e-19

R18_83 V18 V83 -15133.616609062403
L18_83 V18 V83 -3.400693800451935e-12
C18_83 V18 V83 -1.5976756820417408e-19

R18_84 V18 V84 212177.9726524916
L18_84 V18 V84 -3.002512651588092e-12
C18_84 V18 V84 -1.9089665001450625e-19

R18_85 V18 V85 -22366.18165382968
L18_85 V18 V85 8.260120065578999e-12
C18_85 V18 V85 1.0576396139077212e-19

R18_86 V18 V86 2380.078173930862
L18_86 V18 V86 5.6195592359335445e-11
C18_86 V18 V86 1.5312763448531324e-19

R18_87 V18 V87 -26068.57673775101
L18_87 V18 V87 1.4654259063308677e-11
C18_87 V18 V87 9.59766583903763e-20

R18_88 V18 V88 -22698.9861801282
L18_88 V18 V88 9.131028981623702e-12
C18_88 V18 V88 1.6828599425069183e-19

R18_89 V18 V89 -12920.170257738195
L18_89 V18 V89 -2.4832299619853752e-11
C18_89 V18 V89 -1.3420711197116248e-20

R18_90 V18 V90 -2136.2968330447084
L18_90 V18 V90 -6.833251830154954e-12
C18_90 V18 V90 -2.50216556570853e-19

R18_91 V18 V91 20862.44472117794
L18_91 V18 V91 5.046430917990098e-12
C18_91 V18 V91 2.07744989583792e-20

R18_92 V18 V92 29165.361337063256
L18_92 V18 V92 9.913504302272304e-12
C18_92 V18 V92 -5.078698529470634e-20

R18_93 V18 V93 29955.55430319279
L18_93 V18 V93 -1.5634474395573304e-11
C18_93 V18 V93 -9.827138514397361e-20

R18_94 V18 V94 -4174.422207510895
L18_94 V18 V94 -2.1879988820959642e-11
C18_94 V18 V94 1.9586255059337986e-20

R18_95 V18 V95 7843.108414839269
L18_95 V18 V95 -8.412967240178528e-12
C18_95 V18 V95 -4.6734720493737004e-20

R18_96 V18 V96 14342.15454533007
L18_96 V18 V96 -6.384018991656204e-12
C18_96 V18 V96 -7.138050703554643e-20

R18_97 V18 V97 -6989.355174958898
L18_97 V18 V97 7.288311179237367e-12
C18_97 V18 V97 -5.63437903720833e-20

R18_98 V18 V98 2086.5408461711
L18_98 V18 V98 3.841955406810592e-12
C18_98 V18 V98 1.3035072857495272e-19

R18_99 V18 V99 -2534.7069664561186
L18_99 V18 V99 -6.247389210128627e-12
C18_99 V18 V99 -3.877543853844195e-20

R18_100 V18 V100 -4017.4672035499298
L18_100 V18 V100 2.8200518807386405e-10
C18_100 V18 V100 7.532058928362357e-20

R18_101 V18 V101 10198.346004049381
L18_101 V18 V101 -3.9602836838261026e-11
C18_101 V18 V101 9.096581056056638e-20

R18_102 V18 V102 -3026.4317466973057
L18_102 V18 V102 1.461708799901092e-11
C18_102 V18 V102 -1.3072142682744105e-19

R18_103 V18 V103 4950.63334178803
L18_103 V18 V103 1.526700319746757e-11
C18_103 V18 V103 1.8437527817168235e-20

R18_104 V18 V104 4151.623055017663
L18_104 V18 V104 4.3150890581729847e-11
C18_104 V18 V104 -1.4322096701745544e-20

R18_105 V18 V105 -43280.175924836214
L18_105 V18 V105 2.7563307622278465e-11
C18_105 V18 V105 8.500889428843351e-20

R18_106 V18 V106 1218.0818022589738
L18_106 V18 V106 -1.7569961302350933e-12
C18_106 V18 V106 7.509441056723255e-20

R18_107 V18 V107 9450.398815892508
L18_107 V18 V107 1.6777915767275815e-11
C18_107 V18 V107 2.4100129757077295e-20

R18_108 V18 V108 -269552.87033237214
L18_108 V18 V108 -1.1555885680906267e-11
C18_108 V18 V108 2.0241371915623795e-21

R18_109 V18 V109 -4985.657499323025
L18_109 V18 V109 4.336284246647172e-12
C18_109 V18 V109 -6.24446027669262e-20

R18_110 V18 V110 -1563.5157356547188
L18_110 V18 V110 4.086622609951509e-12
C18_110 V18 V110 -1.7857340805568644e-20

R18_111 V18 V111 -8203.69977336461
L18_111 V18 V111 -6.472256679744005e-11
C18_111 V18 V111 2.5274086436350905e-20

R18_112 V18 V112 -7267.1704457418855
L18_112 V18 V112 1.6510424150666308e-11
C18_112 V18 V112 -1.1502339712908826e-20

R18_113 V18 V113 7816.466290557087
L18_113 V18 V113 -5.3817312945148194e-12
C18_113 V18 V113 -1.6136545849885463e-19

R18_114 V18 V114 -1809.0375133703499
L18_114 V18 V114 1.83136424743104e-12
C18_114 V18 V114 3.485652593069228e-20

R18_115 V18 V115 -11144.58137900467
L18_115 V18 V115 -1.3385446386340254e-11
C18_115 V18 V115 -4.940069358871575e-20

R18_116 V18 V116 -23217.99381917632
L18_116 V18 V116 -4.386369182953919e-11
C18_116 V18 V116 -2.7656707282048085e-20

R18_117 V18 V117 -11890.282071418744
L18_117 V18 V117 -3.43832468405729e-12
C18_117 V18 V117 4.551633322421735e-20

R18_118 V18 V118 884.2616395431778
L18_118 V18 V118 -1.2220184094926685e-12
C18_118 V18 V118 -4.47596706528157e-20

R18_119 V18 V119 6313.937638652953
L18_119 V18 V119 -1.3045991092526456e-11
C18_119 V18 V119 5.207908132267322e-20

R18_120 V18 V120 11767.123196969233
L18_120 V18 V120 -8.41323198460358e-12
C18_120 V18 V120 7.189145475732291e-20

R18_121 V18 V121 17730.43279551943
L18_121 V18 V121 2.3391379765375572e-12
C18_121 V18 V121 1.646413822898206e-19

R18_122 V18 V122 -67789.35178385528
L18_122 V18 V122 4.015184110417084e-11
C18_122 V18 V122 -5.1984361037135106e-20

R18_123 V18 V123 7665.90430566925
L18_123 V18 V123 1.4552380281333e-11
C18_123 V18 V123 6.4345927913244514e-21

R18_124 V18 V124 5226.819568274718
L18_124 V18 V124 8.561493309258954e-12
C18_124 V18 V124 -5.47285654623928e-20

R18_125 V18 V125 4629.698535784659
L18_125 V18 V125 7.259507491085711e-12
C18_125 V18 V125 -3.0257578580932866e-20

R18_126 V18 V126 -1343.575046370849
L18_126 V18 V126 1.1805816307617358e-12
C18_126 V18 V126 2.175271909074995e-19

R18_127 V18 V127 -2627.0346737628875
L18_127 V18 V127 5.443890280961206e-12
C18_127 V18 V127 -2.6379971408986984e-20

R18_128 V18 V128 -2636.7227925487546
L18_128 V18 V128 7.783730647079209e-12
C18_128 V18 V128 -1.2409611170812829e-21

R18_129 V18 V129 -3069.903636460019
L18_129 V18 V129 -5.632654253364421e-12
C18_129 V18 V129 -5.166851245078859e-20

R18_130 V18 V130 6500.610026361373
L18_130 V18 V130 -1.7586874501471384e-12
C18_130 V18 V130 -1.1066795782412579e-19

R18_131 V18 V131 3080.9137436464353
L18_131 V18 V131 -3.354746302471016e-12
C18_131 V18 V131 -8.962843885205404e-21

R18_132 V18 V132 2694.4081608745564
L18_132 V18 V132 -2.6464276416172446e-12
C18_132 V18 V132 -7.233227219581719e-21

R18_133 V18 V133 -5133.255087721471
L18_133 V18 V133 -5.825607832639135e-12
C18_133 V18 V133 -5.569638684878923e-20

R18_134 V18 V134 1081.9444041045729
L18_134 V18 V134 -4.989784054212681e-12
C18_134 V18 V134 -5.2587266748767334e-20

R18_135 V18 V135 2937.3467998607994
L18_135 V18 V135 -3.0737399760885615e-11
C18_135 V18 V135 4.0288539327602505e-20

R18_136 V18 V136 2050.1761538549536
L18_136 V18 V136 -9.62114846546499e-12
C18_136 V18 V136 -5.980321702180743e-20

R18_137 V18 V137 1309.812362062409
L18_137 V18 V137 -1.1011593723703983e-10
C18_137 V18 V137 -5.129108821770228e-20

R18_138 V18 V138 -1736.0756548344461
L18_138 V18 V138 1.7789920238181562e-12
C18_138 V18 V138 1.1586975635084052e-19

R18_139 V18 V139 -1708.75610216482
L18_139 V18 V139 3.610669852255772e-12
C18_139 V18 V139 5.781330976738375e-22

R18_140 V18 V140 -1416.0828536703707
L18_140 V18 V140 1.991531339331465e-12
C18_140 V18 V140 1.1017964168646338e-19

R18_141 V18 V141 216486.29635857834
L18_141 V18 V141 3.562104379907967e-12
C18_141 V18 V141 1.5181067893344535e-19

R18_142 V18 V142 -666.0215839372856
L18_142 V18 V142 1.3759054845343191e-11
C18_142 V18 V142 -6.40558768683111e-20

R18_143 V18 V143 7601.812706741213
L18_143 V18 V143 -4.7068256663059904e-12
C18_143 V18 V143 -4.9155877736531135e-20

R18_144 V18 V144 -10020.555423604997
L18_144 V18 V144 -3.890563409287711e-12
C18_144 V18 V144 -1.7379018289471796e-20

R18_145 V18 V145 -1204.2024979763796
L18_145 V18 V145 8.604000225866047e-11
C18_145 V18 V145 3.774424297641201e-20

R18_146 V18 V146 538.9266804912912
L18_146 V18 V146 -1.0781113346713742e-12
C18_146 V18 V146 -1.4868423658519466e-20

R18_147 V18 V147 6278.7486015573895
L18_147 V18 V147 -2.236537374008367e-11
C18_147 V18 V147 7.15332445626007e-20

R18_148 V18 V148 1446.9669759689127
L18_148 V18 V148 1.9519453171172483e-11
C18_148 V18 V148 3.983442754137176e-21

R18_149 V18 V149 3362.914391313071
L18_149 V18 V149 -2.907368958257586e-12
C18_149 V18 V149 -5.228471784784234e-20

R18_150 V18 V150 926.2197128226095
L18_150 V18 V150 2.1801070136675452e-12
C18_150 V18 V150 4.609966195493214e-20

R18_151 V18 V151 -1797.53222210484
L18_151 V18 V151 4.0308356485820554e-12
C18_151 V18 V151 4.063109120270797e-21

R18_152 V18 V152 -778.9517806903024
L18_152 V18 V152 5.422908438245987e-12
C18_152 V18 V152 -1.0441917469710079e-20

R18_153 V18 V153 1323.9408733864393
L18_153 V18 V153 7.881872274340081e-12
C18_153 V18 V153 -1.3101888571744562e-19

R18_154 V18 V154 -1034.1878298397146
L18_154 V18 V154 1.499833250159772e-12
C18_154 V18 V154 -1.7088652776973688e-20

R18_155 V18 V155 7317.017343812868
L18_155 V18 V155 -6.4533887545742045e-12
C18_155 V18 V155 -2.1759165509688903e-20

R18_156 V18 V156 750.5938035678081
L18_156 V18 V156 -1.1983932409226318e-11
C18_156 V18 V156 -2.0647098552544272e-20

R18_157 V18 V157 -2161.8412954620867
L18_157 V18 V157 2.9666121549182552e-12
C18_157 V18 V157 -6.918104397949808e-20

R18_158 V18 V158 -1094.444905982792
L18_158 V18 V158 -1.4241193114734784e-12
C18_158 V18 V158 -5.578618666333307e-20

R18_159 V18 V159 887.5475674974587
L18_159 V18 V159 -4.642237769093786e-12
C18_159 V18 V159 -3.304545864764339e-20

R18_160 V18 V160 1462.8373834408626
L18_160 V18 V160 -3.715090506184665e-12
C18_160 V18 V160 1.1428636334221208e-20

R18_161 V18 V161 -1763.5864275964607
L18_161 V18 V161 1.795845391520248e-11
C18_161 V18 V161 1.6363808769453373e-19

R18_162 V18 V162 1501.394401808274
L18_162 V18 V162 -1.8976035100738016e-12
C18_162 V18 V162 -9.544004567986801e-21

R18_163 V18 V163 -1160.9121994298443
L18_163 V18 V163 6.985333166521247e-12
C18_163 V18 V163 -3.5562622921885274e-20

R18_164 V18 V164 -1049.311268895104
L18_164 V18 V164 2.668546082209581e-12
C18_164 V18 V164 2.5511627376479923e-20

R18_165 V18 V165 1664.0961057986763
L18_165 V18 V165 -7.054471616285412e-11
C18_165 V18 V165 8.525694274613374e-20

R18_166 V18 V166 641.6611512671963
L18_166 V18 V166 8.60076993305924e-13
C18_166 V18 V166 2.106492856517734e-20

R18_167 V18 V167 -4911.7775417056655
L18_167 V18 V167 -1.3145857822766364e-11
C18_167 V18 V167 4.3086017818426146e-20

R18_168 V18 V168 -2330.553397746075
L18_168 V18 V168 -2.9739001822800588e-12
C18_168 V18 V168 4.456553813411021e-20

R18_169 V18 V169 1670.4658774036975
L18_169 V18 V169 -2.2200364552283255e-11
C18_169 V18 V169 -9.943429943620716e-20

R18_170 V18 V170 -606.0003751210053
L18_170 V18 V170 -2.9615510256286846e-12
C18_170 V18 V170 7.56048209924525e-20

R18_171 V18 V171 1644.421674586835
L18_171 V18 V171 -1.7056324562614994e-10
C18_171 V18 V171 5.768384394337838e-20

R18_172 V18 V172 1294.1873098195147
L18_172 V18 V172 7.505740015046394e-11
C18_172 V18 V172 8.961723758291426e-21

R18_173 V18 V173 -1494.8159658780828
L18_173 V18 V173 -8.023880925093095e-12
C18_173 V18 V173 -1.4076250226781445e-19

R18_174 V18 V174 -1256.6674443036752
L18_174 V18 V174 -1.090288232210346e-12
C18_174 V18 V174 -1.2826030792151257e-19

R18_175 V18 V175 -21310.15239287967
L18_175 V18 V175 3.383895686551892e-11
C18_175 V18 V175 -1.0862794729204811e-19

R18_176 V18 V176 -201433.37091157725
L18_176 V18 V176 5.489433688240421e-12
C18_176 V18 V176 -1.0341280424499596e-19

R18_177 V18 V177 17231.346485331644
L18_177 V18 V177 1.3817289316468999e-11
C18_177 V18 V177 9.971836716000067e-20

R18_178 V18 V178 634.3827364041589
L18_178 V18 V178 2.0791525117594297e-12
C18_178 V18 V178 5.984539561859425e-22

R18_179 V18 V179 -5015.493638992478
L18_179 V18 V179 2.1073125429049962e-10
C18_179 V18 V179 2.471830342403677e-21

R18_180 V18 V180 -5129.5798886712155
L18_180 V18 V180 -1.5365819889045054e-11
C18_180 V18 V180 2.932818060410326e-20

R18_181 V18 V181 3040.6449420188515
L18_181 V18 V181 -3.29613640925763e-11
C18_181 V18 V181 1.3604397768212616e-19

R18_182 V18 V182 -6770.870467381652
L18_182 V18 V182 5.780956322515363e-12
C18_182 V18 V182 -1.2132114459347887e-20

R18_183 V18 V183 4608.728515034868
L18_183 V18 V183 7.484467443889222e-11
C18_183 V18 V183 9.7746527694851e-21

R18_184 V18 V184 5895.703546898693
L18_184 V18 V184 1.5315059296629416e-11
C18_184 V18 V184 6.181571384297195e-20

R18_185 V18 V185 -5879.435861127811
L18_185 V18 V185 4.368466871439375e-12
C18_185 V18 V185 -1.2423790756554618e-19

R18_186 V18 V186 -1753.6467749028502
L18_186 V18 V186 9.080817522930178e-11
C18_186 V18 V186 9.539384787664422e-20

R18_187 V18 V187 -9755.294352685194
L18_187 V18 V187 5.590452642733743e-12
C18_187 V18 V187 6.67228370310438e-20

R18_188 V18 V188 -2376.2620292805605
L18_188 V18 V188 3.3544295842338903e-12
C18_188 V18 V188 5.976706957868214e-20

R18_189 V18 V189 4247.0294990709535
L18_189 V18 V189 -8.025090858274986e-12
C18_189 V18 V189 -1.8696154379487546e-20

R18_190 V18 V190 1760.4019788051883
L18_190 V18 V190 -3.2501336026614335e-12
C18_190 V18 V190 -3.790059656053348e-20

R18_191 V18 V191 -27493.703346100923
L18_191 V18 V191 -2.821909847865261e-11
C18_191 V18 V191 -4.467647494456239e-21

R18_192 V18 V192 5687.737806894048
L18_192 V18 V192 -7.880394749735249e-12
C18_192 V18 V192 -1.1413707788663734e-19

R18_193 V18 V193 -3879.4622740543205
L18_193 V18 V193 -4.187351313396694e-12
C18_193 V18 V193 -5.2156130010973705e-20

R18_194 V18 V194 -4835.675099656603
L18_194 V18 V194 6.75363249305235e-11
C18_194 V18 V194 -9.461671813663541e-20

R18_195 V18 V195 4548.192708140777
L18_195 V18 V195 -5.833178543878607e-11
C18_195 V18 V195 -7.018070344450582e-20

R18_196 V18 V196 4039.275733165972
L18_196 V18 V196 -5.95893003161798e-12
C18_196 V18 V196 -6.908754772797701e-21

R18_197 V18 V197 -3724.9789608575543
L18_197 V18 V197 4.4886116792286026e-12
C18_197 V18 V197 1.1198062767187517e-19

R18_198 V18 V198 -2952.8897866728084
L18_198 V18 V198 3.171763550048318e-12
C18_198 V18 V198 3.01952506095497e-20

R18_199 V18 V199 -5735.002332457715
L18_199 V18 V199 1.591167716086748e-11
C18_199 V18 V199 -5.441442104238222e-20

R18_200 V18 V200 -2774.6863970767163
L18_200 V18 V200 4.12672126632891e-12
C18_200 V18 V200 9.97121215202212e-20

R19_19 V19 0 -588.243124822847
L19_19 V19 0 -1.997817277229542e-12
C19_19 V19 0 3.4650046259862242e-19

R19_20 V19 V20 -3346.127127092701
L19_20 V19 V20 -1.6870825718591118e-12
C19_20 V19 V20 -5.180466590038366e-19

R19_21 V19 V21 -8472.019059559856
L19_21 V19 V21 -1.4043747708025223e-11
C19_21 V19 V21 1.2346277094262733e-19

R19_22 V19 V22 -4533.771259215443
L19_22 V19 V22 2.6659517505868136e-11
C19_22 V19 V22 7.156013010702088e-20

R19_23 V19 V23 -2949.978249706771
L19_23 V19 V23 1.2589221628253115e-12
C19_23 V19 V23 7.854219254760717e-19

R19_24 V19 V24 -7480.119802280101
L19_24 V19 V24 3.132247854235799e-12
C19_24 V19 V24 2.9152593861577105e-19

R19_25 V19 V25 6140.25547608531
L19_25 V19 V25 2.118996866738976e-12
C19_25 V19 V25 2.070643493768446e-19

R19_26 V19 V26 4101.309022358013
L19_26 V19 V26 2.0059396249254904e-12
C19_26 V19 V26 2.9821223410526244e-19

R19_27 V19 V27 4689.655696047706
L19_27 V19 V27 1.3690456969279706e-12
C19_27 V19 V27 2.3329043716841244e-19

R19_28 V19 V28 6456.322219899964
L19_28 V19 V28 2.4081780856446036e-12
C19_28 V19 V28 1.7005928770184438e-19

R19_29 V19 V29 10276.566426422127
L19_29 V19 V29 -1.6852083926120186e-11
C19_29 V19 V29 -1.5767414602263004e-19

R19_30 V19 V30 10054.361156200497
L19_30 V19 V30 -4.056439922027444e-12
C19_30 V19 V30 -1.9867776660665537e-19

R19_31 V19 V31 904.4565475543039
L19_31 V19 V31 -1.467759849216267e-12
C19_31 V19 V31 -4.461674318901525e-19

R19_32 V19 V32 2752.3908845982437
L19_32 V19 V32 -3.2251802134848247e-12
C19_32 V19 V32 -1.5580080104981125e-19

R19_33 V19 V33 -14480.704167371705
L19_33 V19 V33 1.5052966997425183e-11
C19_33 V19 V33 5.2841180109317904e-20

R19_34 V19 V34 -8505.867836391337
L19_34 V19 V34 -4.943826163102081e-12
C19_34 V19 V34 -1.9457725053108139e-19

R19_35 V19 V35 -2380.181800894843
L19_35 V19 V35 3.12711476038565e-12
C19_35 V19 V35 3.4883957572711296e-19

R19_36 V19 V36 -4620.439510217303
L19_36 V19 V36 -1.0183817491301515e-11
C19_36 V19 V36 4.6969889962141374e-20

R19_37 V19 V37 -10089.769028836465
L19_37 V19 V37 -1.1595593691662654e-11
C19_37 V19 V37 -1.0268086026040016e-20

R19_38 V19 V38 -26896.073515571952
L19_38 V19 V38 3.0680618718449926e-12
C19_38 V19 V38 2.949793845176291e-19

R19_39 V19 V39 -1038.8686595946456
L19_39 V19 V39 -4.1306789287640375e-10
C19_39 V19 V39 -1.3392929142318076e-19

R19_40 V19 V40 -2014.13104280808
L19_40 V19 V40 6.8806823504437794e-12
C19_40 V19 V40 -5.088631184603912e-22

R19_41 V19 V41 9357.48235145551
L19_41 V19 V41 -1.2082721319941424e-11
C19_41 V19 V41 -7.535651633464363e-20

R19_42 V19 V42 12187.924033345776
L19_42 V19 V42 -7.071267073688724e-11
C19_42 V19 V42 -8.365767274436675e-20

R19_43 V19 V43 -16166.328548295232
L19_43 V19 V43 -2.07063052935073e-11
C19_43 V19 V43 4.286530778626358e-20

R19_44 V19 V44 5757.132024244547
L19_44 V19 V44 -1.2427150890609596e-11
C19_44 V19 V44 1.1190662955030151e-20

R19_45 V19 V45 8475.834563163224
L19_45 V19 V45 3.948523142711106e-12
C19_45 V19 V45 1.151364397040761e-19

R19_46 V19 V46 10723.330320748097
L19_46 V19 V46 -3.172418407516895e-12
C19_46 V19 V46 -2.716175928133363e-19

R19_47 V19 V47 1309.0632151083205
L19_47 V19 V47 -6.649002400933397e-12
C19_47 V19 V47 2.5990175501007147e-20

R19_48 V19 V48 3959.4235598103046
L19_48 V19 V48 -1.4942935520554027e-11
C19_48 V19 V48 -6.047742632388638e-20

R19_49 V19 V49 -19412.413529476707
L19_49 V19 V49 -1.930795096196928e-11
C19_49 V19 V49 -5.648389513160345e-20

R19_50 V19 V50 56427.70419224995
L19_50 V19 V50 3.0256138247979105e-12
C19_50 V19 V50 2.8209576903827527e-19

R19_51 V19 V51 3020.5759620743074
L19_51 V19 V51 -3.819391885666681e-12
C19_51 V19 V51 -3.015146881766913e-19

R19_52 V19 V52 -75818.09067369574
L19_52 V19 V52 6.836999095305124e-12
C19_52 V19 V52 1.2816496192809152e-19

R19_53 V19 V53 11050.751296257646
L19_53 V19 V53 -1.0399771664740581e-11
C19_53 V19 V53 -9.046660718835423e-20

R19_54 V19 V54 66721.12302341974
L19_54 V19 V54 -1.409189237276834e-11
C19_54 V19 V54 -5.1229677362565296e-20

R19_55 V19 V55 -3291.8482720109428
L19_55 V19 V55 1.6349432058343928e-12
C19_55 V19 V55 3.8234075102730535e-19

R19_56 V19 V56 -5893.624838512207
L19_56 V19 V56 -8.640852914170723e-12
C19_56 V19 V56 -2.5461571147719218e-20

R19_57 V19 V57 -10695.061079823548
L19_57 V19 V57 6.056594061688584e-12
C19_57 V19 V57 7.033840984018263e-20

R19_58 V19 V58 5524.748944964008
L19_58 V19 V58 -1.695460487354512e-11
C19_58 V19 V58 -1.090887596967781e-19

R19_59 V19 V59 -2136.007599025797
L19_59 V19 V59 -3.119201670280629e-11
C19_59 V19 V59 1.90147461535507e-20

R19_60 V19 V60 -4807.145411646494
L19_60 V19 V60 -2.414822710626794e-11
C19_60 V19 V60 -8.159159895218053e-20

R19_61 V19 V61 19255.78486675937
L19_61 V19 V61 -4.432698238438843e-11
C19_61 V19 V61 -1.1407101633096965e-20

R19_62 V19 V62 -5329.9520716086845
L19_62 V19 V62 5.02678206384572e-12
C19_62 V19 V62 8.284227395429003e-20

R19_63 V19 V63 36952.59874486669
L19_63 V19 V63 -1.5266670495989338e-12
C19_63 V19 V63 -4.532561742251549e-19

R19_64 V19 V64 6976.483497912998
L19_64 V19 V64 8.916608461974533e-12
C19_64 V19 V64 8.974649915839244e-20

R19_65 V19 V65 18220.328206020182
L19_65 V19 V65 -6.288309582091257e-12
C19_65 V19 V65 -1.0499894300660002e-19

R19_66 V19 V66 24223.786791492494
L19_66 V19 V66 -1.122380957408161e-11
C19_66 V19 V66 -4.9884510776972247e-20

R19_67 V19 V67 2330.932250240761
L19_67 V19 V67 4.928496918456087e-12
C19_67 V19 V67 1.2229488434690223e-19

R19_68 V19 V68 5177.146182840147
L19_68 V19 V68 -1.4040843231789903e-11
C19_68 V19 V68 -1.5366479816831265e-20

R19_69 V19 V69 41958.684661522006
L19_69 V19 V69 3.4805579935337566e-12
C19_69 V19 V69 1.7276814830690697e-19

R19_70 V19 V70 12440.227545110038
L19_70 V19 V70 -6.751835649359179e-12
C19_70 V19 V70 -4.1260621042893075e-20

R19_71 V19 V71 2561.0126331484785
L19_71 V19 V71 1.8240675257904245e-12
C19_71 V19 V71 3.4466925648837437e-19

R19_72 V19 V72 9454.135323917788
L19_72 V19 V72 -8.253862336519088e-12
C19_72 V19 V72 -1.2078895104540867e-19

R19_73 V19 V73 7652.967555915913
L19_73 V19 V73 1.1134435545959476e-11
C19_73 V19 V73 -1.4835766328499366e-20

R19_74 V19 V74 -12571.42441554005
L19_74 V19 V74 3.95579773658741e-12
C19_74 V19 V74 7.436078627233993e-20

R19_75 V19 V75 -1876.066507509766
L19_75 V19 V75 -1.9230089034761596e-12
C19_75 V19 V75 -2.743507594949384e-19

R19_76 V19 V76 -4062.7442655503482
L19_76 V19 V76 4.506941952009689e-12
C19_76 V19 V76 1.9948319912214915e-19

R19_77 V19 V77 -4934.969930353417
L19_77 V19 V77 -3.874978356877636e-12
C19_77 V19 V77 -1.5503046408976484e-19

R19_78 V19 V78 8183.6517457783575
L19_78 V19 V78 -7.02045448083509e-11
C19_78 V19 V78 7.839298743057701e-20

R19_79 V19 V79 -2248.551379391099
L19_79 V19 V79 -7.364143269801612e-12
C19_79 V19 V79 -2.031551469405252e-19

R19_80 V19 V80 -5508.047948996732
L19_80 V19 V80 -1.7940908934434385e-11
C19_80 V19 V80 -5.022801599906514e-20

R19_81 V19 V81 9634.263167266994
L19_81 V19 V81 9.689234762465171e-12
C19_81 V19 V81 4.6965768602574374e-20

R19_82 V19 V82 -7728.9082183988885
L19_82 V19 V82 -5.26313597456877e-12
C19_82 V19 V82 -1.6168006437081135e-19

R19_83 V19 V83 4913.131578534801
L19_83 V19 V83 3.049444703921819e-12
C19_83 V19 V83 2.751745980939688e-19

R19_84 V19 V84 8604.718846243835
L19_84 V19 V84 -3.529876827533988e-12
C19_84 V19 V84 -1.4376947646460134e-19

R19_85 V19 V85 -42458.739253763415
L19_85 V19 V85 9.919800913892753e-12
C19_85 V19 V85 5.873659641635157e-20

R19_86 V19 V86 5533.959113111296
L19_86 V19 V86 1.3879406591660977e-11
C19_86 V19 V86 -4.001036069434625e-21

R19_87 V19 V87 1311.7481318044015
L19_87 V19 V87 -4.880912168299725e-12
C19_87 V19 V87 1.1565278065542997e-19

R19_88 V19 V88 7826.059308308078
L19_88 V19 V88 5.753788927247735e-12
C19_88 V19 V88 1.995234907878956e-19

R19_89 V19 V89 8916.06515077794
L19_89 V19 V89 1.5732608826102816e-11
C19_89 V19 V89 7.198434452850934e-20

R19_90 V19 V90 8997.639032010868
L19_90 V19 V90 7.118132214468233e-12
C19_90 V19 V90 1.9395091393569791e-19

R19_91 V19 V91 -3683.3057524375245
L19_91 V19 V91 3.6060019936946127e-12
C19_91 V19 V91 -3.423684649567431e-19

R19_92 V19 V92 29696.004295786814
L19_92 V19 V92 2.5605985725678593e-11
C19_92 V19 V92 -8.801176192923284e-20

R19_93 V19 V93 7606.0526387686705
L19_93 V19 V93 -1.9310689570974213e-11
C19_93 V19 V93 -5.4180110698574647e-20

R19_94 V19 V94 -5398.368518564375
L19_94 V19 V94 -1.134639384441771e-11
C19_94 V19 V94 -6.944835616411042e-20

R19_95 V19 V95 -838.2057149201154
L19_95 V19 V95 7.896991357343407e-12
C19_95 V19 V95 3.509522854056001e-20

R19_96 V19 V96 -2483.0394423676225
L19_96 V19 V96 -9.942489156168614e-12
C19_96 V19 V96 -9.426432391161044e-20

R19_97 V19 V97 -2215.274825557182
L19_97 V19 V97 -5.016532255298033e-11
C19_97 V19 V97 -2.34343293039556e-19

R19_98 V19 V98 14143.348810097203
L19_98 V19 V98 -2.4550678696278782e-11
C19_98 V19 V98 -1.626927335456579e-19

R19_99 V19 V99 831.2952395780704
L19_99 V19 V99 -2.204981788645407e-12
C19_99 V19 V99 2.6766641019278536e-19

R19_100 V19 V100 10377.065586684863
L19_100 V19 V100 -2.0546895052935847e-11
C19_100 V19 V100 1.54905387095239e-19

R19_101 V19 V101 6569.594004407419
L19_101 V19 V101 2.2329400608909655e-11
C19_101 V19 V101 1.4276092521057266e-19

R19_102 V19 V102 -23924.062978507198
L19_102 V19 V102 7.262365726560912e-12
C19_102 V19 V102 6.128137248331035e-20

R19_103 V19 V103 -43946.33942199849
L19_103 V19 V103 3.569172173971074e-12
C19_103 V19 V103 -1.8951400684758771e-19

R19_104 V19 V104 3920.880445409267
L19_104 V19 V104 1.946334215147793e-11
C19_104 V19 V104 -7.660324705632106e-20

R19_105 V19 V105 2245.4944079701036
L19_105 V19 V105 8.032176060364269e-12
C19_105 V19 V105 1.4208480039805746e-19

R19_106 V19 V106 1922.0731241842282
L19_106 V19 V106 -4.947597341304635e-12
C19_106 V19 V106 2.2862208694404956e-19

R19_107 V19 V107 -2278.0881272512083
L19_107 V19 V107 5.885472555887473e-12
C19_107 V19 V107 -2.003807222750636e-20

R19_108 V19 V108 -26283.43185166982
L19_108 V19 V108 4.129653737626941e-11
C19_108 V19 V108 2.3713633450353667e-20

R19_109 V19 V109 -6440.888893339491
L19_109 V19 V109 9.811020038824672e-12
C19_109 V19 V109 -1.8444925646776515e-19

R19_110 V19 V110 -2397.229004950924
L19_110 V19 V110 -2.2942303226121675e-10
C19_110 V19 V110 -1.3238908475736034e-19

R19_111 V19 V111 830.2863957122023
L19_111 V19 V111 -1.6802811541932987e-12
C19_111 V19 V111 -2.4727378904403734e-20

R19_112 V19 V112 3806.5030684272765
L19_112 V19 V112 -6.51297881808339e-12
C19_112 V19 V112 -8.5897277474181e-22

R19_113 V19 V113 -4003.278600936765
L19_113 V19 V113 -4.8661401579704206e-12
C19_113 V19 V113 -1.3682407230526306e-19

R19_114 V19 V114 -1833.846196108887
L19_114 V19 V114 6.5790371113866974e-12
C19_114 V19 V114 -1.9739490407534818e-19

R19_115 V19 V115 -845.1203775907719
L19_115 V19 V115 2.758792159644962e-12
C19_115 V19 V115 1.0930450466153411e-19

R19_116 V19 V116 -1764.3618946378788
L19_116 V19 V116 9.442293486116624e-12
C19_116 V19 V116 -5.535112662205854e-20

R19_117 V19 V117 -3115.9672668791113
L19_117 V19 V117 -5.8623310794043736e-12
C19_117 V19 V117 1.2524040067151446e-19

R19_118 V19 V118 1149.9063887532084
L19_118 V19 V118 -5.078508671724798e-12
C19_118 V19 V118 2.3040465559458604e-19

R19_119 V19 V119 1262.0896821561705
L19_119 V19 V119 3.663763510473688e-12
C19_119 V19 V119 2.0270125184206308e-20

R19_120 V19 V120 2506.690121535446
L19_120 V19 V120 9.103126369682685e-12
C19_120 V19 V120 1.5830786308844116e-19

R19_121 V19 V121 2882.209624313271
L19_121 V19 V121 2.135933026271465e-12
C19_121 V19 V121 4.9429857452586957e-20

R19_122 V19 V122 -303852.4960679218
L19_122 V19 V122 6.381266694802094e-11
C19_122 V19 V122 4.906340190111984e-21

R19_123 V19 V123 1727.6902363234622
L19_123 V19 V123 -1.6321884765998385e-12
C19_123 V19 V123 -2.5374749223520505e-19

R19_124 V19 V124 2371.5101240590825
L19_124 V19 V124 -3.851674004056341e-12
C19_124 V19 V124 -1.4618779094573094e-19

R19_125 V19 V125 1059.2085324816846
L19_125 V19 V125 6.432760783415442e-12
C19_125 V19 V125 3.7161697309686585e-21

R19_126 V19 V126 -3733.042010050291
L19_126 V19 V126 1.3406654544854038e-11
C19_126 V19 V126 -1.0338586424947766e-19

R19_127 V19 V127 -808.0778177981308
L19_127 V19 V127 4.6403400154366115e-12
C19_127 V19 V127 1.9205246802611462e-19

R19_128 V19 V128 -1426.384826026058
L19_128 V19 V128 3.8319848992534514e-11
C19_128 V19 V128 -6.002746183936998e-20

R19_129 V19 V129 -865.8411417262379
L19_129 V19 V129 -2.2934003461051802e-12
C19_129 V19 V129 -9.707572411950046e-20

R19_130 V19 V130 -2914.7569268002167
L19_130 V19 V130 -1.875903884266936e-11
C19_130 V19 V130 4.119772202433305e-20

R19_131 V19 V131 1355.2420823796194
L19_131 V19 V131 7.501276137333683e-11
C19_131 V19 V131 2.5826179680461657e-20

R19_132 V19 V132 1745.0869378617922
L19_132 V19 V132 5.299071407548555e-12
C19_132 V19 V132 1.9795110680168232e-19

R19_133 V19 V133 -1652.2048784787055
L19_133 V19 V133 4.1779604461093215e-11
C19_133 V19 V133 -2.144394677513891e-20

R19_134 V19 V134 3016.4677807925164
L19_134 V19 V134 2.6729206168782448e-11
C19_134 V19 V134 3.597217481765412e-20

R19_135 V19 V135 1708.3350462625176
L19_135 V19 V135 -2.4595692114339223e-12
C19_135 V19 V135 -3.2128913694167146e-19

R19_136 V19 V136 1883.1539730512584
L19_136 V19 V136 -6.963673404738042e-12
C19_136 V19 V136 -1.196861084846749e-19

R19_137 V19 V137 724.741559632058
L19_137 V19 V137 4.758011897353607e-12
C19_137 V19 V137 3.2141774832482684e-20

R19_138 V19 V138 -4276.467976105239
L19_138 V19 V138 -5.283937861695751e-11
C19_138 V19 V138 -6.95130302694806e-20

R19_139 V19 V139 -1238.752134274528
L19_139 V19 V139 1.1751486306646014e-12
C19_139 V19 V139 4.376770353854905e-19

R19_140 V19 V140 -965.8165069530469
L19_140 V19 V140 3.882847157814897e-12
C19_140 V19 V140 1.1290044340924803e-19

R19_141 V19 V141 1775.9577499165425
L19_141 V19 V141 -3.039709056712085e-10
C19_141 V19 V141 -2.370890194078865e-20

R19_142 V19 V142 -1854.0398055702808
L19_142 V19 V142 -1.1018695834416222e-11
C19_142 V19 V142 -7.184388773470317e-21

R19_143 V19 V143 5897.872382043971
L19_143 V19 V143 -1.991845507676859e-12
C19_143 V19 V143 -1.4111456095924476e-19

R19_144 V19 V144 2831.2762086875846
L19_144 V19 V144 -5.581588380672967e-12
C19_144 V19 V144 -1.861940857281019e-20

R19_145 V19 V145 -630.395178041626
L19_145 V19 V145 -3.6458940465267945e-12
C19_145 V19 V145 -5.066894871299751e-20

R19_146 V19 V146 2580.0474160398976
L19_146 V19 V146 -4.156412186474123e-12
C19_146 V19 V146 5.1301159364639263e-20

R19_147 V19 V147 -647.3231805728992
L19_147 V19 V147 -1.5940276140200735e-12
C19_147 V19 V147 -2.2513330099440676e-19

R19_148 V19 V148 -2728.274460963745
L19_148 V19 V148 -7.410005868992841e-12
C19_148 V19 V148 -5.1651406490620294e-20

R19_149 V19 V149 10007.13150279071
L19_149 V19 V149 5.892012457282669e-12
C19_149 V19 V149 1.9225531736689294e-19

R19_150 V19 V150 742.7975706245544
L19_150 V19 V150 3.5431965007630984e-12
C19_150 V19 V150 -7.488352147175516e-20

R19_151 V19 V151 225.13733382025762
L19_151 V19 V151 1.367945328898822e-12
C19_151 V19 V151 1.230552890458118e-19

R19_152 V19 V152 3641.1195217968348
L19_152 V19 V152 1.1868550662712928e-11
C19_152 V19 V152 -1.7279662231222398e-20

R19_153 V19 V153 1228.612485755395
L19_153 V19 V153 2.9183923115357527e-12
C19_153 V19 V153 -6.172676862468898e-20

R19_154 V19 V154 -8619.79829170959
L19_154 V19 V154 2.5967782577330987e-12
C19_154 V19 V154 -4.910377050818451e-21

R19_155 V19 V155 -136.23275512571493
L19_155 V19 V155 1.5614639434892298e-12
C19_155 V19 V155 2.7428954997126315e-19

R19_156 V19 V156 2379.0290733428374
L19_156 V19 V156 6.785036942932351e-12
C19_156 V19 V156 4.925802559105534e-20

R19_157 V19 V157 20861.602971534583
L19_157 V19 V157 1.2306140929787015e-11
C19_157 V19 V157 -2.471073545900036e-19

R19_158 V19 V158 -10169.018520844651
L19_158 V19 V158 -3.1531352839057974e-12
C19_158 V19 V158 4.765791237506822e-20

R19_159 V19 V159 683.9438045965122
L19_159 V19 V159 -9.598133503925956e-13
C19_159 V19 V159 -2.6089794196620996e-19

R19_160 V19 V160 -70788.62505382652
L19_160 V19 V160 -1.524309726019812e-11
C19_160 V19 V160 9.603878169608731e-21

R19_161 V19 V161 -5365.655678133939
L19_161 V19 V161 -6.004975285090729e-12
C19_161 V19 V161 1.601873690307606e-19

R19_162 V19 V162 8937.826512704338
L19_162 V19 V162 -5.934468902584662e-12
C19_162 V19 V162 2.7541072385659376e-20

R19_163 V19 V163 518.3316832242631
L19_163 V19 V163 -1.841764136270132e-12
C19_163 V19 V163 6.258007113751634e-20

R19_164 V19 V164 1675.9337851064734
L19_164 V19 V164 -5.608443001083394e-12
C19_164 V19 V164 3.695944429066453e-20

R19_165 V19 V165 3942.4719737684886
L19_165 V19 V165 3.9303302921913307e-11
C19_165 V19 V165 8.226059005007856e-20

R19_166 V19 V166 2592.0420803016655
L19_166 V19 V166 2.949924765485251e-12
C19_166 V19 V166 -3.352118480991676e-20

R19_167 V19 V167 1315.171681001376
L19_167 V19 V167 7.965329093224191e-13
C19_167 V19 V167 3.849920410334006e-20

R19_168 V19 V168 -1020.8605619708261
L19_168 V19 V168 -1.0853213863348935e-11
C19_168 V19 V168 3.995133406831425e-20

R19_169 V19 V169 1763.721910611405
L19_169 V19 V169 -3.2452978137733773e-10
C19_169 V19 V169 -1.7331365945135615e-19

R19_170 V19 V170 8119.723115991244
L19_170 V19 V170 -3.811671807595743e-12
C19_170 V19 V170 4.788613705095478e-20

R19_171 V19 V171 -308.536138360978
L19_171 V19 V171 -7.793075275526378e-12
C19_171 V19 V171 4.6721960261130197e-20

R19_172 V19 V172 -5256.425894580979
L19_172 V19 V172 1.3705948336121002e-11
C19_172 V19 V172 -1.056622805144965e-20

R19_173 V19 V173 -1991.0712109309018
L19_173 V19 V173 -1.0241730182164742e-11
C19_173 V19 V173 -2.288904711239592e-20

R19_174 V19 V174 -1128.373323086392
L19_174 V19 V174 -3.9024494268026533e-11
C19_174 V19 V174 -9.102407680310465e-20

R19_175 V19 V175 544.7500716043625
L19_175 V19 V175 -1.3387899167343635e-12
C19_175 V19 V175 6.541791999653625e-20

R19_176 V19 V176 -32727.8064120871
L19_176 V19 V176 -1.1620323478293658e-11
C19_176 V19 V176 -2.4758246985472625e-20

R19_177 V19 V177 1965.3270445086391
L19_177 V19 V177 2.037715596530271e-11
C19_177 V19 V177 4.926936001843145e-20

R19_178 V19 V178 1553.3627481151234
L19_178 V19 V178 6.947145894848556e-11
C19_178 V19 V178 -2.389822085465247e-20

R19_179 V19 V179 -881.2672695578945
L19_179 V19 V179 2.8062408809095763e-12
C19_179 V19 V179 -1.4415709153473365e-19

R19_180 V19 V180 2161.5769985277166
L19_180 V19 V180 2.5012116602311957e-10
C19_180 V19 V180 -5.92439889826697e-20

R19_181 V19 V181 -6022.38613324515
L19_181 V19 V181 -2.374987810360677e-11
C19_181 V19 V181 6.316361538337372e-20

R19_182 V19 V182 -2080.3271252465106
L19_182 V19 V182 1.0919204960436489e-11
C19_182 V19 V182 7.495557422075091e-20

R19_183 V19 V183 922.9276350036283
L19_183 V19 V183 1.4287321725571041e-11
C19_183 V19 V183 -2.4607161977183768e-20

R19_184 V19 V184 50786.52101385591
L19_184 V19 V184 2.7525498995917008e-11
C19_184 V19 V184 2.2389655832664836e-20

R19_185 V19 V185 -7559.487158614388
L19_185 V19 V185 4.376671310627127e-12
C19_185 V19 V185 -4.862683692584345e-20

R19_186 V19 V186 -3338.8917901966856
L19_186 V19 V186 3.965425798945139e-12
C19_186 V19 V186 2.053570709712125e-20

R19_187 V19 V187 23619.18753292182
L19_187 V19 V187 -1.0744704143946645e-11
C19_187 V19 V187 1.9020275488108019e-19

R19_188 V19 V188 -913.5060343057409
L19_188 V19 V188 3.69238381912794e-12
C19_188 V19 V188 1.1226561222245048e-19

R19_189 V19 V189 2470.234369988435
L19_189 V19 V189 -1.3474272304835312e-11
C19_189 V19 V189 -3.6537722647082787e-20

R19_190 V19 V190 1916.2598696881287
L19_190 V19 V190 -5.225081416677542e-12
C19_190 V19 V190 -6.9480507044008e-20

R19_191 V19 V191 -2348.3573925929545
L19_191 V19 V191 9.326909887245542e-12
C19_191 V19 V191 -9.011833288955921e-20

R19_192 V19 V192 3127.9710258708446
L19_192 V19 V192 -1.1549690826448403e-11
C19_192 V19 V192 -1.1057854790976746e-19

R19_193 V19 V193 -5529.498569701025
L19_193 V19 V193 -3.8039647318385366e-12
C19_193 V19 V193 -6.055917788172962e-20

R19_194 V19 V194 -8492.477702806284
L19_194 V19 V194 -1.3609128702456988e-11
C19_194 V19 V194 -1.1094775798870872e-19

R19_195 V19 V195 3063.346845722032
L19_195 V19 V195 4.3205699161186854e-11
C19_195 V19 V195 9.375701893656345e-20

R19_196 V19 V196 678.732244861575
L19_196 V19 V196 -5.36310324860023e-12
C19_196 V19 V196 -5.032780923218579e-20

R19_197 V19 V197 7892.240151879522
L19_197 V19 V197 8.224963874483607e-12
C19_197 V19 V197 8.952347752242984e-20

R19_198 V19 V198 4254.599924390306
L19_198 V19 V198 8.701471973930764e-12
C19_198 V19 V198 -2.6883654316138236e-21

R19_199 V19 V199 -4216.373098851086
L19_199 V19 V199 -9.572290533167978e-12
C19_199 V19 V199 -2.9030791864117895e-20

R19_200 V19 V200 -1481.9548241756502
L19_200 V19 V200 8.575986814645709e-12
C19_200 V19 V200 1.0839251223460768e-19

R20_20 V20 0 -186.8636109392712
L20_20 V20 0 -9.556287398282664e-13
C20_20 V20 0 9.797172235557469e-19

R20_21 V20 V21 -4505.14162193042
L20_21 V20 V21 -8.069139044747687e-12
C20_21 V20 V21 1.487180866043261e-19

R20_22 V20 V22 -3300.547406890804
L20_22 V20 V22 1.3281089114225222e-11
C20_22 V20 V22 1.0664108285885549e-19

R20_23 V20 V23 -5298.860540694987
L20_23 V20 V23 2.832979158768278e-12
C20_23 V20 V23 3.628545334824423e-19

R20_24 V20 V24 -2522.3149775225347
L20_24 V20 V24 9.307696328081135e-13
C20_24 V20 V24 1.0013261183520355e-18

R20_25 V20 V25 3956.1318125414446
L20_25 V20 V25 1.4765656301965315e-12
C20_25 V20 V25 2.8508266120290154e-19

R20_26 V20 V26 3244.480457878515
L20_26 V20 V26 1.5506203092912742e-12
C20_26 V20 V26 3.5665583373362675e-19

R20_27 V20 V27 4801.647420590304
L20_27 V20 V27 2.2054509682570892e-12
C20_27 V20 V27 1.3498630753342637e-19

R20_28 V20 V28 3125.786836380703
L20_28 V20 V28 9.43284483518962e-13
C20_28 V20 V28 3.507526318675886e-19

R20_29 V20 V29 5637.179088181525
L20_29 V20 V29 -2.2108061170884005e-11
C20_29 V20 V29 -1.9834109051703972e-19

R20_30 V20 V30 6925.075303372591
L20_30 V20 V30 -3.121218712818585e-12
C20_30 V20 V30 -2.5206390406334227e-19

R20_31 V20 V31 2229.9259921318394
L20_31 V20 V31 -3.09254514832376e-12
C20_31 V20 V31 -2.435616921434171e-19

R20_32 V20 V32 729.3567129093997
L20_32 V20 V32 -1.1050743321803287e-12
C20_32 V20 V32 -4.87512318198355e-19

R20_33 V20 V33 -7800.874638258469
L20_33 V20 V33 5.8463974695865e-11
C20_33 V20 V33 2.7589561243008015e-20

R20_34 V20 V34 -4332.78591087883
L20_34 V20 V34 -3.2048270059517645e-12
C20_34 V20 V34 -2.848738306800627e-19

R20_35 V20 V35 -4855.058175075743
L20_35 V20 V35 -2.5875528118924515e-11
C20_35 V20 V35 3.747659252769219e-21

R20_36 V20 V36 -1434.072885119824
L20_36 V20 V36 7.617687903682314e-12
C20_36 V20 V36 4.357661146706583e-19

R20_37 V20 V37 -5800.9295464215775
L20_37 V20 V37 -7.354974839890556e-12
C20_37 V20 V37 -8.794552402758523e-21

R20_38 V20 V38 -11306.658848220093
L20_38 V20 V38 2.3838445070299756e-12
C20_38 V20 V38 3.9111563090015607e-19

R20_39 V20 V39 -2122.055630976318
L20_39 V20 V39 4.9191538911462185e-12
C20_39 V20 V39 6.542002113151879e-20

R20_40 V20 V40 -737.0201484600402
L20_40 V20 V40 5.4972764776431985e-12
C20_40 V20 V40 -1.4775673407806145e-20

R20_41 V20 V41 6691.392113588552
L20_41 V20 V41 -1.0305121124415514e-11
C20_41 V20 V41 -1.0653973824741632e-19

R20_42 V20 V42 10149.965730501212
L20_42 V20 V42 -3.243864125533687e-11
C20_42 V20 V42 -1.4208885479986887e-19

R20_43 V20 V43 5404.049137308236
L20_43 V20 V43 -9.087284572571365e-12
C20_43 V20 V43 -7.479409402748789e-20

R20_44 V20 V44 9921.03381205688
L20_44 V20 V44 -6.449514138136698e-12
C20_44 V20 V44 1.6741372790086558e-20

R20_45 V20 V45 4841.196979328451
L20_45 V20 V45 2.55482221663809e-12
C20_45 V20 V45 1.688564768858169e-19

R20_46 V20 V46 5822.465754847726
L20_46 V20 V46 -2.7295127126202442e-12
C20_46 V20 V46 -3.4523914110272224e-19

R20_47 V20 V47 2921.3358087101706
L20_47 V20 V47 -9.504157564676076e-12
C20_47 V20 V47 -7.639733689288995e-20

R20_48 V20 V48 856.2212387133084
L20_48 V20 V48 -6.0999577450202735e-12
C20_48 V20 V48 -4.6770457161847595e-20

R20_49 V20 V49 -11186.943080686371
L20_49 V20 V49 -1.2567170886504962e-11
C20_49 V20 V49 -8.793945259739824e-20

R20_50 V20 V50 -32623.88771966463
L20_50 V20 V50 2.4447274704287543e-12
C20_50 V20 V50 3.475006361425701e-19

R20_51 V20 V51 8933.594723478593
L20_51 V20 V51 4.2117037373042345e-12
C20_51 V20 V51 1.2127281360706969e-19

R20_52 V20 V52 11079.871186723707
L20_52 V20 V52 -7.555553820379746e-12
C20_52 V20 V52 -1.0096561570403874e-19

R20_53 V20 V53 10171.920061225746
L20_53 V20 V53 -4.864892417085406e-12
C20_53 V20 V53 -1.7125202271853674e-19

R20_54 V20 V54 -16304.111222730595
L20_54 V20 V54 -6.608312776131393e-12
C20_54 V20 V54 -9.24684248561624e-20

R20_55 V20 V55 -22192.516238485314
L20_55 V20 V55 -1.2645964716877753e-11
C20_55 V20 V55 -6.141912519649809e-20

R20_56 V20 V56 -1364.0476128921073
L20_56 V20 V56 2.0682735693435157e-12
C20_56 V20 V56 4.509179914733444e-19

R20_57 V20 V57 -7023.89589290389
L20_57 V20 V57 4.569953109850119e-12
C20_57 V20 V57 9.532756840801351e-20

R20_58 V20 V58 3606.295191906977
L20_58 V20 V58 -9.768686518006425e-12
C20_58 V20 V58 -1.8043592478265086e-19

R20_59 V20 V59 -4873.516689128897
L20_59 V20 V59 -3.010051606672247e-11
C20_59 V20 V59 -1.5174837914489668e-19

R20_60 V20 V60 -1601.8410549122636
L20_60 V20 V60 -6.595749677616024e-12
C20_60 V20 V60 -1.956267396945151e-20

R20_61 V20 V61 10432.909884045166
L20_61 V20 V61 2.3560002653129105e-11
C20_61 V20 V61 2.93926452876928e-20

R20_62 V20 V62 -4308.106908729176
L20_62 V20 V62 3.318271445118461e-12
C20_62 V20 V62 1.352710857351078e-19

R20_63 V20 V63 10419.68095858973
L20_63 V20 V63 8.126108853020219e-12
C20_63 V20 V63 1.2695994760327224e-19

R20_64 V20 V64 3379.1093573466887
L20_64 V20 V64 -1.8560520657141617e-12
C20_64 V20 V64 -3.926460032654868e-19

R20_65 V20 V65 10359.018912070142
L20_65 V20 V65 -3.989941669215632e-12
C20_65 V20 V65 -1.8061011929455825e-19

R20_66 V20 V66 138246.43726748537
L20_66 V20 V66 -7.784980829041444e-12
C20_66 V20 V66 -8.365375990962493e-20

R20_67 V20 V67 28426.19983215426
L20_67 V20 V67 -6.974547818743053e-12
C20_67 V20 V67 -3.872518131011259e-20

R20_68 V20 V68 1630.385983399896
L20_68 V20 V68 4.7590439510181185e-12
C20_68 V20 V68 9.071023933141452e-20

R20_69 V20 V69 -29133.74441312788
L20_69 V20 V69 2.8012706812502876e-12
C20_69 V20 V69 2.3047189289592006e-19

R20_70 V20 V70 9466.96324854681
L20_70 V20 V70 -4.224832603895763e-12
C20_70 V20 V70 -6.537743660885165e-20

R20_71 V20 V71 8277.67714520951
L20_71 V20 V71 -1.8993458268223918e-11
C20_71 V20 V71 -9.573393698896147e-20

R20_72 V20 V72 2057.536429942009
L20_72 V20 V72 1.9582905136145023e-12
C20_72 V20 V72 3.7345979438629925e-19

R20_73 V20 V73 6814.816229227582
L20_73 V20 V73 6.0100599588215746e-12
C20_73 V20 V73 6.7538055911352836e-21

R20_74 V20 V74 -7703.160354417724
L20_74 V20 V74 2.765114371463823e-12
C20_74 V20 V74 1.2360720008933024e-19

R20_75 V20 V75 15816.416608319456
L20_75 V20 V75 5.0845827347367875e-12
C20_75 V20 V75 8.443632082409171e-20

R20_76 V20 V76 -865.9131355541415
L20_76 V20 V76 -2.2217013611786033e-12
C20_76 V20 V76 -1.226531284587553e-19

R20_77 V20 V77 -4519.783006915029
L20_77 V20 V77 -2.804208303618226e-12
C20_77 V20 V77 -2.146729852791009e-19

R20_78 V20 V78 3905.704338659329
L20_78 V20 V78 -6.971823062791608e-11
C20_78 V20 V78 8.649412131996016e-20

R20_79 V20 V79 -2870.6606064454554
L20_79 V20 V79 -3.516887388766797e-11
C20_79 V20 V79 2.435262324742605e-21

R20_80 V20 V80 -9411.99289015767
L20_80 V20 V80 -4.406774752282804e-12
C20_80 V20 V80 -3.0129749337246114e-19

R20_81 V20 V81 3665.5286004739946
L20_81 V20 V81 8.067589392375681e-12
C20_81 V20 V81 4.264742656899789e-21

R20_82 V20 V82 -5875.510727223822
L20_82 V20 V82 -3.5942181973209363e-12
C20_82 V20 V82 -2.2798774247110466e-19

R20_83 V20 V83 8502.452226665528
L20_83 V20 V83 -5.199574384171532e-12
C20_83 V20 V83 -1.335086333632819e-19

R20_84 V20 V84 2792.699762922316
L20_84 V20 V84 5.068354271872161e-12
C20_84 V20 V84 2.1463319449469182e-19

R20_85 V20 V85 -17216.64385077763
L20_85 V20 V85 6.821017960319819e-12
C20_85 V20 V85 9.533021684941835e-20

R20_86 V20 V86 7083.195942032181
L20_86 V20 V86 8.742485525242028e-12
C20_86 V20 V86 1.2085652108675984e-21

R20_87 V20 V87 4414.671566373206
L20_87 V20 V87 1.2941542029041291e-11
C20_87 V20 V87 1.4609457458346454e-19

R20_88 V20 V88 1275.711760714575
L20_88 V20 V88 -9.147717711213696e-12
C20_88 V20 V88 2.246642131398908e-19

R20_89 V20 V89 19978.207435711414
L20_89 V20 V89 1.548997432885795e-11
C20_89 V20 V89 8.716675334108525e-20

R20_90 V20 V90 9358.028059078004
L20_90 V20 V90 5.486890744395033e-12
C20_90 V20 V90 2.161323965878164e-19

R20_91 V20 V91 3544.224247809616
L20_91 V20 V91 7.533760846180418e-12
C20_91 V20 V91 -1.4706984470280657e-19

R20_92 V20 V92 -1734.0957968396713
L20_92 V20 V92 3.3781223805761104e-12
C20_92 V20 V92 -3.252447344790385e-19

R20_93 V20 V93 3492.262308860766
L20_93 V20 V93 -1.0722082696850229e-11
C20_93 V20 V93 -9.816678291017847e-20

R20_94 V20 V94 -7429.940768585762
L20_94 V20 V94 -5.977082203941533e-12
C20_94 V20 V94 -1.174808509804383e-19

R20_95 V20 V95 -2096.837823419643
L20_95 V20 V95 -1.2122295419023506e-11
C20_95 V20 V95 -6.608232899591562e-20

R20_96 V20 V96 -603.3289370668346
L20_96 V20 V96 1.1281402862018925e-11
C20_96 V20 V96 -1.0083283391980211e-20

R20_97 V20 V97 -1704.3364105617861
L20_97 V20 V97 -9.721363819327857e-11
C20_97 V20 V97 -3.0770725043692102e-19

R20_98 V20 V98 13624.131575049007
L20_98 V20 V98 -1.13289993357264e-09
C20_98 V20 V98 -1.915110005172167e-19

R20_99 V20 V99 16227.635322433864
L20_99 V20 V99 -1.3138209090245047e-11
C20_99 V20 V99 1.3473989362784677e-19

R20_100 V20 V100 486.29133101030504
L20_100 V20 V100 -1.6202496520919306e-12
C20_100 V20 V100 3.2255689587756856e-19

R20_101 V20 V101 4656.87747583171
L20_101 V20 V101 1.4152531932746906e-11
C20_101 V20 V101 1.7553584668741692e-19

R20_102 V20 V102 -11029.770652622647
L20_102 V20 V102 4.826103974371017e-12
C20_102 V20 V102 8.961542772833111e-20

R20_103 V20 V103 3001.79543935433
L20_103 V20 V103 7.357966836647105e-12
C20_103 V20 V103 -6.625296621141587e-20

R20_104 V20 V104 -69074.47985367438
L20_104 V20 V104 3.0210352129469044e-12
C20_104 V20 V104 -2.1348452238678108e-19

R20_105 V20 V105 1635.0473464832546
L20_105 V20 V105 7.515922290032081e-12
C20_105 V20 V105 1.628135178943912e-19

R20_106 V20 V106 1314.9175412959685
L20_106 V20 V106 -2.773684837281653e-12
C20_106 V20 V106 2.3476430348361947e-19

R20_107 V20 V107 37696.579473093974
L20_107 V20 V107 -2.5363753997832586e-11
C20_107 V20 V107 -6.426758587419605e-20

R20_108 V20 V108 -966.3761044594938
L20_108 V20 V108 3.1004918197949713e-12
C20_108 V20 V108 8.778476996033855e-20

R20_109 V20 V109 -2045.822809801646
L20_109 V20 V109 5.056083365484639e-12
C20_109 V20 V109 -2.4092208840508946e-19

R20_110 V20 V110 -1363.6095049594674
L20_110 V20 V110 1.424689253317227e-11
C20_110 V20 V110 -1.0933331384704093e-19

R20_111 V20 V111 2372.035770547667
L20_111 V20 V111 -4.040983852968764e-12
C20_111 V20 V111 6.315254271269016e-20

R20_112 V20 V112 816.2246121241695
L20_112 V20 V112 -1.379027034790358e-12
C20_112 V20 V112 -2.2299911170769503e-19

R20_113 V20 V113 -8302.468241884082
L20_113 V20 V113 -3.152969695207194e-12
C20_113 V20 V113 -1.7197349591319528e-19

R20_114 V20 V114 -1538.3871320675157
L20_114 V20 V114 4.9959797179579074e-12
C20_114 V20 V114 -2.1967517839434565e-19

R20_115 V20 V115 -900.6130765159284
L20_115 V20 V115 4.459956480040363e-12
C20_115 V20 V115 1.304588085885103e-20

R20_116 V20 V116 -997.4600969324187
L20_116 V20 V116 5.35430291210581e-12
C20_116 V20 V116 8.189990294155081e-20

R20_117 V20 V117 -2772.917737407257
L20_117 V20 V117 -3.5163490232732826e-12
C20_117 V20 V117 1.7332037986693922e-19

R20_118 V20 V118 774.9697679527695
L20_118 V20 V118 -2.9839912494812487e-12
C20_118 V20 V118 2.436237524433006e-19

R20_119 V20 V119 1594.1129609786424
L20_119 V20 V119 1.069279440903797e-11
C20_119 V20 V119 1.481299623785165e-19

R20_120 V20 V120 788.8443963467531
L20_120 V20 V120 2.0701488093960283e-12
C20_120 V20 V120 2.7108372514143806e-19

R20_121 V20 V121 4664.570948368066
L20_121 V20 V121 1.473935036696625e-12
C20_121 V20 V121 5.3676096978182627e-20

R20_122 V20 V122 -5953.744604372242
L20_122 V20 V122 1.1385120635197474e-11
C20_122 V20 V122 3.885198493695853e-20

R20_123 V20 V123 1795.9819377564622
L20_123 V20 V123 -3.057515021749661e-12
C20_123 V20 V123 -1.1884928381539703e-19

R20_124 V20 V124 -17040.54732562016
L20_124 V20 V124 -1.334446681090658e-12
C20_124 V20 V124 -5.378919827997976e-19

R20_125 V20 V125 796.2123197233956
L20_125 V20 V125 4.042254780496949e-12
C20_125 V20 V125 -1.9918461141802313e-20

R20_126 V20 V126 -2708.933081300956
L20_126 V20 V126 6.212613192051665e-12
C20_126 V20 V126 -8.867529058547567e-20

R20_127 V20 V127 -925.3303009120103
L20_127 V20 V127 1.0415211793029827e-11
C20_127 V20 V127 -1.1161150959018787e-19

R20_128 V20 V128 -635.4714881609517
L20_128 V20 V128 6.2435680491650305e-12
C20_128 V20 V128 1.3406918703831205e-19

R20_129 V20 V129 -643.3765393964513
L20_129 V20 V129 -1.6751592049844234e-12
C20_129 V20 V129 -1.038079067944041e-19

R20_130 V20 V130 -2859.7876923300505
L20_130 V20 V130 -6.81496312602708e-12
C20_130 V20 V130 4.948829319480227e-20

R20_131 V20 V131 1020.1166007266274
L20_131 V20 V131 1.7360989715437654e-11
C20_131 V20 V131 1.6145889781014772e-19

R20_132 V20 V132 572.5016455729591
L20_132 V20 V132 6.104153236622673e-12
C20_132 V20 V132 2.2234193078261636e-19

R20_133 V20 V133 -1885.4979326373382
L20_133 V20 V133 -6.47905543258354e-11
C20_133 V20 V133 1.604718196772613e-20

R20_134 V20 V134 1351.577004734572
L20_134 V20 V134 1.3908302400116126e-11
C20_134 V20 V134 1.1132168282036008e-19

R20_135 V20 V135 4080.3673392682535
L20_135 V20 V135 -6.4677543194427654e-12
C20_135 V20 V135 1.0521510423244527e-20

R20_136 V20 V136 1369.2063273881824
L20_136 V20 V136 -2.1139037850066287e-12
C20_136 V20 V136 -4.631726507169141e-19

R20_137 V20 V137 642.6313841805751
L20_137 V20 V137 3.917587443570387e-12
C20_137 V20 V137 -1.689578297535409e-21

R20_138 V20 V138 -1589.2786897805227
L20_138 V20 V138 1.3461032846761647e-10
C20_138 V20 V138 -1.0274126472214712e-19

R20_139 V20 V139 -714.5324150425765
L20_139 V20 V139 2.687739521624921e-12
C20_139 V20 V139 3.731835576379631e-20

R20_140 V20 V140 -1252.6789743517697
L20_140 V20 V140 1.1532903576508354e-12
C20_140 V20 V140 5.031232362499915e-19

R20_141 V20 V141 1775.2089068212433
L20_141 V20 V141 1.246828681574865e-11
C20_141 V20 V141 -1.1836749737552901e-20

R20_142 V20 V142 -1035.4959970935654
L20_142 V20 V142 -7.1582653333568576e-12
C20_142 V20 V142 -1.8464529910614843e-20

R20_143 V20 V143 1237.6598233620255
L20_143 V20 V143 -2.5218489312839396e-12
C20_143 V20 V143 -8.731739938155771e-20

R20_144 V20 V144 -469.14796673978304
L20_144 V20 V144 -1.6734632040527167e-12
C20_144 V20 V144 -3.9059417530726836e-20

R20_145 V20 V145 -522.3883927277109
L20_145 V20 V145 -2.8764998228450697e-12
C20_145 V20 V145 -4.141966626918488e-20

R20_146 V20 V146 1869.1955489013246
L20_146 V20 V146 -2.6004993799214202e-12
C20_146 V20 V146 5.876659963987119e-20

R20_147 V20 V147 -1246.7961142999736
L20_147 V20 V147 -3.23358421376861e-12
C20_147 V20 V147 -7.608637090360315e-20

R20_148 V20 V148 265.5580995787442
L20_148 V20 V148 -2.3625765786525318e-12
C20_148 V20 V148 -3.3145121479662464e-19

R20_149 V20 V149 6626.95976123052
L20_149 V20 V149 2.133712019469028e-11
C20_149 V20 V149 1.9282756213180074e-19

R20_150 V20 V150 505.81020124800466
L20_150 V20 V150 2.6727085577168485e-12
C20_150 V20 V150 -1.22622314858374e-19

R20_151 V20 V151 1128.8076883412155
L20_151 V20 V151 2.3085919971028935e-12
C20_151 V20 V151 5.509084718132439e-20

R20_152 V20 V152 -3388.29459330371
L20_152 V20 V152 1.8113291392025346e-12
C20_152 V20 V152 1.0294886190332475e-19

R20_153 V20 V153 1516.932893403617
L20_153 V20 V153 1.86541333208124e-12
C20_153 V20 V153 -6.521577309605076e-20

R20_154 V20 V154 -866.5053310027125
L20_154 V20 V154 1.6342772123990022e-12
C20_154 V20 V154 1.086779960947883e-20

R20_155 V20 V155 -413.88318845940677
L20_155 V20 V155 3.0478101256361384e-12
C20_155 V20 V155 9.879311554665346e-20

R20_156 V20 V156 1884.0523286639504
L20_156 V20 V156 1.1615765485363086e-12
C20_156 V20 V156 2.1052554190047783e-19

R20_157 V20 V157 1509.9475498290897
L20_157 V20 V157 4.564891439796989e-12
C20_157 V20 V157 -3.469050725158755e-19

R20_158 V20 V158 1720.4356771814173
L20_158 V20 V158 -2.109637841318793e-12
C20_158 V20 V158 2.640039442535361e-20

R20_159 V20 V159 458.6539764410025
L20_159 V20 V159 -4.212167910185695e-12
C20_159 V20 V159 -8.167134367188442e-20

R20_160 V20 V160 -329.08620138870907
L20_160 V20 V160 -8.939881316349018e-13
C20_160 V20 V160 -1.3207410857996628e-19

R20_161 V20 V161 -1582.9898179907232
L20_161 V20 V161 -5.959522341892257e-12
C20_161 V20 V161 1.9050663374676868e-19

R20_162 V20 V162 11725.358452656545
L20_162 V20 V162 -4.106695277152315e-12
C20_162 V20 V162 5.4004799525893386e-21

R20_163 V20 V163 4670.811996415769
L20_163 V20 V163 -4.623189464345908e-12
C20_163 V20 V163 -5.942656083089567e-20

R20_164 V20 V164 225.85747086944963
L20_164 V20 V164 -2.0965784300177473e-12
C20_164 V20 V164 7.824047558741879e-20

R20_165 V20 V165 976.3956924837771
L20_165 V20 V165 3.517615516319044e-11
C20_165 V20 V165 9.269442577343785e-20

R20_166 V20 V166 1225.8348297280927
L20_166 V20 V166 1.7968438126378577e-12
C20_166 V20 V166 -7.219589276246328e-20

R20_167 V20 V167 1034.9675384036566
L20_167 V20 V167 1.4278053142970217e-11
C20_167 V20 V167 4.5787601956519184e-20

R20_168 V20 V168 -347.18847895750474
L20_168 V20 V168 7.527911941701065e-13
C20_168 V20 V168 9.041420077793827e-20

R20_169 V20 V169 2016.6387890734409
L20_169 V20 V169 3.091606058221976e-11
C20_169 V20 V169 -2.2981668465670105e-19

R20_170 V20 V170 -5741.405787582882
L20_170 V20 V170 -3.8190281320567374e-12
C20_170 V20 V170 6.261776992637435e-20

R20_171 V20 V171 -784.1504755001093
L20_171 V20 V171 4.829817464121162e-12
C20_171 V20 V171 5.84564249736077e-20

R20_172 V20 V172 -829.3769410669764
L20_172 V20 V172 -3.3477609333246277e-12
C20_172 V20 V172 -4.1302907622105365e-21

R20_173 V20 V173 -1374.3596398743093
L20_173 V20 V173 -8.445791044974092e-12
C20_173 V20 V173 -3.228651143636456e-20

R20_174 V20 V174 -847.8623547667083
L20_174 V20 V174 -5.00125181213796e-12
C20_174 V20 V174 -1.0522525899780596e-19

R20_175 V20 V175 3306.4929436297243
L20_175 V20 V175 -1.0850369865800064e-11
C20_175 V20 V175 -3.1965723504191135e-20

R20_176 V20 V176 571.233453815431
L20_176 V20 V176 -1.1806069587841383e-12
C20_176 V20 V176 1.140067992542238e-19

R20_177 V20 V177 1338.3236922919205
L20_177 V20 V177 4.8017865719546115e-11
C20_177 V20 V177 4.6980456219683076e-20

R20_178 V20 V178 1081.3343318840941
L20_178 V20 V178 -3.7092008019599327e-09
C20_178 V20 V178 -3.000461065415974e-20

R20_179 V20 V179 -6063.602048469798
L20_179 V20 V179 -6.6994672508090016e-12
C20_179 V20 V179 -1.0243000132000915e-19

R20_180 V20 V180 19425.075052789558
L20_180 V20 V180 2.4175965767421544e-12
C20_180 V20 V180 -1.9846121001186713e-19

R20_181 V20 V181 -3745.18731622965
L20_181 V20 V181 -1.306727660176195e-11
C20_181 V20 V181 8.486819405152134e-20

R20_182 V20 V182 -1327.1952021659029
L20_182 V20 V182 6.839000295602889e-12
C20_182 V20 V182 7.402201162688113e-20

R20_183 V20 V183 2028.5754020730478
L20_183 V20 V183 -1.9062186128375996e-11
C20_183 V20 V183 -2.7638521332575405e-20

R20_184 V20 V184 -28587.260011895953
L20_184 V20 V184 5.307992966324121e-12
C20_184 V20 V184 7.322134461754945e-20

R20_185 V20 V185 -9170.851500816274
L20_185 V20 V185 2.6250096293201573e-12
C20_185 V20 V185 -5.640613532836384e-20

R20_186 V20 V186 -7591.595182148966
L20_186 V20 V186 3.1393704022435606e-12
C20_186 V20 V186 7.219439999231975e-20

R20_187 V20 V187 -3038.4573017418547
L20_187 V20 V187 3.0263189949004854e-12
C20_187 V20 V187 1.6124984100485374e-19

R20_188 V20 V188 -602.3825580113726
L20_188 V20 V188 1.1138225156348932e-11
C20_188 V20 V188 1.7434469080594008e-19

R20_189 V20 V189 3325.8673905259684
L20_189 V20 V189 -1.133530917963828e-11
C20_189 V20 V189 -3.229089517275955e-20

R20_190 V20 V190 1203.52465533315
L20_190 V20 V190 -4.355405572127528e-12
C20_190 V20 V190 -1.0624446738208056e-19

R20_191 V20 V191 -3270.195053644851
L20_191 V20 V191 8.446205479014708e-12
C20_191 V20 V191 -1.6388981836527092e-20

R20_192 V20 V192 3025.32862310752
L20_192 V20 V192 -7.72559642099033e-12
C20_192 V20 V192 -2.221923673424052e-19

R20_193 V20 V193 -1745.8706884030362
L20_193 V20 V193 -2.4002555430838908e-12
C20_193 V20 V193 -9.493281456024636e-20

R20_194 V20 V194 13072.247566533208
L20_194 V20 V194 -6.132043577189356e-12
C20_194 V20 V194 -1.946371170325059e-19

R20_195 V20 V195 1295.693080842117
L20_195 V20 V195 -4.745706906605619e-12
C20_195 V20 V195 -1.7402305929000237e-19

R20_196 V20 V196 648.8103174502522
L20_196 V20 V196 1.4776941880167497e-11
C20_196 V20 V196 2.307048158594635e-19

R20_197 V20 V197 -6369.863784541721
L20_197 V20 V197 6.0530005832396354e-12
C20_197 V20 V197 1.3448868157534103e-19

R20_198 V20 V198 1895.3601502031108
L20_198 V20 V198 5.754021034172124e-12
C20_198 V20 V198 -5.641204906170508e-20

R20_199 V20 V199 634.8475911154115
L20_199 V20 V199 -8.662436312092303e-11
C20_199 V20 V199 -6.980679446857453e-20

R20_200 V20 V200 -459.48835321567674
L20_200 V20 V200 -2.0982923108531676e-11
C20_200 V20 V200 6.773862378502045e-20

R21_21 V21 0 -54.20559197772121
L21_21 V21 0 -1.2539726191172493e-13
C21_21 V21 0 -5.056124282907885e-19

R21_22 V21 V22 -767.1678700755002
L21_22 V21 V22 -1.9230112438215915e-12
C21_22 V21 V22 -8.931179758426822e-21

R21_23 V21 V23 -1267.821015552542
L21_23 V21 V23 -1.6763889217255361e-12
C21_23 V21 V23 -9.867533754481891e-20

R21_24 V21 V24 -914.3792199848646
L21_24 V21 V24 -1.3046780360721923e-12
C21_24 V21 V24 -1.091132172190106e-19

R21_25 V21 V25 221.23782008006935
L21_25 V21 V25 5.908276997713637e-13
C21_25 V21 V25 7.935890079295058e-20

R21_26 V21 V26 1423.2271108418554
L21_26 V21 V26 2.840596749425934e-12
C21_26 V21 V26 -2.5882033480702098e-20

R21_27 V21 V27 2866.3208138936416
L21_27 V21 V27 1.6446382518951735e-12
C21_27 V21 V27 5.607739170896019e-20

R21_28 V21 V28 1667.60085185814
L21_28 V21 V28 1.0567722813221938e-12
C21_28 V21 V28 6.264498023071121e-20

R21_29 V21 V29 231.79546813472143
L21_29 V21 V29 7.108041325629309e-13
C21_29 V21 V29 2.179236468099174e-19

R21_30 V21 V30 2593.627213126951
L21_30 V21 V30 3.0649097006907866e-12
C21_30 V21 V30 1.1379654561202856e-20

R21_31 V21 V31 2804.1220689112492
L21_31 V21 V31 3.5398693396538256e-12
C21_31 V21 V31 -3.3589118704768483e-21

R21_32 V21 V32 1647.775658370974
L21_32 V21 V32 2.6825699620549097e-12
C21_32 V21 V32 -5.118330770074629e-21

R21_33 V21 V33 497.43231520880454
L21_33 V21 V33 1.0514479188877174e-11
C21_33 V21 V33 -2.510707598271851e-19

R21_34 V21 V34 -18720.6717593394
L21_34 V21 V34 6.3104305171336676e-12
C21_34 V21 V34 5.3326881449313096e-20

R21_35 V21 V35 -2618.087350108683
L21_35 V21 V35 -6.950003955769042e-12
C21_35 V21 V35 -4.8360362286263446e-20

R21_36 V21 V36 -1552.850623745096
L21_36 V21 V36 -4.025214330769363e-12
C21_36 V21 V36 -6.365446201673419e-20

R21_37 V21 V37 -607.2215638112775
L21_37 V21 V37 -7.814766502714782e-13
C21_37 V21 V37 9.675647064280884e-20

R21_38 V21 V38 -3498.060796562111
L21_38 V21 V38 -1.6787208519839758e-12
C21_38 V21 V38 -6.233993260328185e-20

R21_39 V21 V39 -3006.5437055758057
L21_39 V21 V39 -2.857411085655103e-12
C21_39 V21 V39 7.53999622604547e-20

R21_40 V21 V40 -1817.3467711601686
L21_40 V21 V40 -2.016802873706457e-12
C21_40 V21 V40 9.910540489971949e-20

R21_41 V21 V41 -2013.6064311054552
L21_41 V21 V41 -4.2575183677643584e-12
C21_41 V21 V41 -7.379672110835947e-20

R21_42 V21 V42 -2558.638985542568
L21_42 V21 V42 -7.017988966081209e-12
C21_42 V21 V42 -4.327129630665458e-20

R21_43 V21 V43 -1748.1013529579689
L21_43 V21 V43 -3.1435177771279704e-12
C21_43 V21 V43 -9.67955005729089e-20

R21_44 V21 V44 -1358.7842597990946
L21_44 V21 V44 -2.8917935365775532e-12
C21_44 V21 V44 -1.2322548716946494e-19

R21_45 V21 V45 487.280540533955
L21_45 V21 V45 8.435655364938576e-13
C21_45 V21 V45 6.351643541774375e-20

R21_46 V21 V46 1024488.5600847317
L21_46 V21 V46 5.3725875351105495e-12
C21_46 V21 V46 8.83979982117588e-20

R21_47 V21 V47 -60952.93857284766
L21_47 V21 V47 3.944817142448353e-12
C21_47 V21 V47 2.1644393185646666e-20

R21_48 V21 V48 4234.36310123097
L21_48 V21 V48 2.100894763289449e-12
C21_48 V21 V48 2.678018406006273e-20

R21_49 V21 V49 405.1867874930351
L21_49 V21 V49 2.2558709929781287e-12
C21_49 V21 V49 1.7919024998810805e-19

R21_50 V21 V50 -6125.291111328188
L21_50 V21 V50 7.184921147062119e-12
C21_50 V21 V50 -8.044920711934601e-21

R21_51 V21 V51 -16245.38595634557
L21_51 V21 V51 2.5425116822161783e-12
C21_51 V21 V51 6.196247925436334e-20

R21_52 V21 V52 -3559.4351795753855
L21_52 V21 V52 2.7751938837279395e-12
C21_52 V21 V52 7.918611050464618e-20

R21_53 V21 V53 683.89790285069
L21_53 V21 V53 5.024809398904506e-12
C21_53 V21 V53 -1.5672301406926724e-19

R21_54 V21 V54 2503.0030719115243
L21_54 V21 V54 6.958160973343731e-12
C21_54 V21 V54 3.05310400747524e-21

R21_55 V21 V55 2125.6745679846977
L21_55 V21 V55 8.361160328727209e-12
C21_55 V21 V55 -2.9332338700818595e-20

R21_56 V21 V56 3239.8127411795185
L21_56 V21 V56 -3.506636379593655e-11
C21_56 V21 V56 -2.980056850901665e-20

R21_57 V21 V57 360635.54729723884
L21_57 V21 V57 -8.117783397165424e-13
C21_57 V21 V57 -9.597742562044318e-20

R21_58 V21 V58 -1978.3820944045929
L21_58 V21 V58 -2.0280084719225362e-12
C21_58 V21 V58 -1.0827842017804065e-19

R21_59 V21 V59 -1269.9336432264765
L21_59 V21 V59 -1.6336958687247595e-12
C21_59 V21 V59 -3.979823887072117e-20

R21_60 V21 V60 -868.7645299034191
L21_60 V21 V60 -1.1177003964295034e-12
C21_60 V21 V60 -6.636285789713712e-20

R21_61 V21 V61 -2118.9723434416765
L21_61 V21 V61 1.3318892984739147e-12
C21_61 V21 V61 1.3780411871116235e-19

R21_62 V21 V62 -22761.254126925316
L21_62 V21 V62 -6.913003862357746e-12
C21_62 V21 V62 1.3377119012835196e-20

R21_63 V21 V63 -10355.031221475623
L21_63 V21 V63 -3.3939129595102333e-12
C21_63 V21 V63 -4.8163521580232676e-20

R21_64 V21 V64 31679.704565845517
L21_64 V21 V64 -8.284253340352172e-12
C21_64 V21 V64 -5.2388769325559286e-20

R21_65 V21 V65 614.9351906686562
L21_65 V21 V65 1.5577126835215538e-12
C21_65 V21 V65 1.1428076703377798e-19

R21_66 V21 V66 -4389.747592223757
L21_66 V21 V66 3.391620802864006e-12
C21_66 V21 V66 1.3131526889434965e-19

R21_67 V21 V67 -5056.525694180982
L21_67 V21 V67 2.1286976852301702e-12
C21_67 V21 V67 1.1884510162138687e-19

R21_68 V21 V68 -10322.042897836476
L21_68 V21 V68 1.1178714531280148e-12
C21_68 V21 V68 1.7603282925436087e-19

R21_69 V21 V69 875.6073886678491
L21_69 V21 V69 5.854465884088259e-12
C21_69 V21 V69 -6.656166745759834e-20

R21_70 V21 V70 -15058.803520560854
L21_70 V21 V70 1.2154007242338252e-11
C21_70 V21 V70 -6.435615300196246e-20

R21_71 V21 V71 27320.268287321403
L21_71 V21 V71 2.8635606007821327e-12
C21_71 V21 V71 3.241174366212949e-20

R21_72 V21 V72 14998.771816029059
L21_72 V21 V72 3.3433294479016356e-12
C21_72 V21 V72 2.58371077834542e-20

R21_73 V21 V73 1267.6667823540165
L21_73 V21 V73 -5.066816744386487e-12
C21_73 V21 V73 -2.192984724711688e-19

R21_74 V21 V74 3860.1764543206064
L21_74 V21 V74 -2.2300376744068496e-12
C21_74 V21 V74 -1.535385627680009e-19

R21_75 V21 V75 8142.714674383721
L21_75 V21 V75 -1.676507358788732e-12
C21_75 V21 V75 -1.8492877142439113e-19

R21_76 V21 V76 -5851.521973494526
L21_76 V21 V76 -9.844669512928437e-13
C21_76 V21 V76 -2.4088701535851785e-19

R21_77 V21 V77 -3480.967971210418
L21_77 V21 V77 -1.507006338711786e-12
C21_77 V21 V77 1.3195352581645783e-19

R21_78 V21 V78 11410.458251819215
L21_78 V21 V78 9.969500380884622e-12
C21_78 V21 V78 1.767107199333698e-20

R21_79 V21 V79 -8930.793561790226
L21_79 V21 V79 -2.9617970555330045e-11
C21_79 V21 V79 8.209625751546438e-20

R21_80 V21 V80 -8672.432124517129
L21_80 V21 V80 5.497410572459521e-12
C21_80 V21 V80 1.382013934080461e-19

R21_81 V21 V81 337.7289295007715
L21_81 V21 V81 7.507440270748875e-13
C21_81 V21 V81 2.340297348273141e-19

R21_82 V21 V82 -2224.539324479333
L21_82 V21 V82 3.2918036370088133e-12
C21_82 V21 V82 2.218590480480906e-19

R21_83 V21 V83 -1246.1150257878862
L21_83 V21 V83 1.322526502999935e-11
C21_83 V21 V83 9.627537582257296e-20

R21_84 V21 V84 -1187.4093361261396
L21_84 V21 V84 3.442873705458656e-12
C21_84 V21 V84 1.647901952097731e-19

R21_85 V21 V85 -15674.116617858872
L21_85 V21 V85 -4.917709182782512e-12
C21_85 V21 V85 -2.819380368518586e-19

R21_86 V21 V86 -988.924090920413
L21_86 V21 V86 -1.0277398901758602e-11
C21_86 V21 V86 -5.949971391741364e-20

R21_87 V21 V87 -3073.404242186522
L21_87 V21 V87 -5.448257527222079e-12
C21_87 V21 V87 -1.2054973058396458e-19

R21_88 V21 V88 -3140.917323744373
L21_88 V21 V88 -5.939779759179663e-12
C21_88 V21 V88 -1.529917125799299e-19

R21_89 V21 V89 1049.9351040494155
L21_89 V21 V89 1.61800078882653e-12
C21_89 V21 V89 6.157882814923276e-20

R21_90 V21 V90 1784.236587804292
L21_90 V21 V90 -2.364408445080762e-12
C21_90 V21 V90 -2.3199838650711458e-19

R21_91 V21 V91 2788.169611224883
L21_91 V21 V91 1.6158895961090364e-12
C21_91 V21 V91 1.0482520526537054e-19

R21_92 V21 V92 12013.461999807841
L21_92 V21 V92 2.862141692797697e-12
C21_92 V21 V92 3.616341501153243e-20

R21_93 V21 V93 728.8010675565936
L21_93 V21 V93 -5.374681184173344e-12
C21_93 V21 V93 1.141767391970395e-19

R21_94 V21 V94 1550.5380291338035
L21_94 V21 V94 4.828672317908685e-12
C21_94 V21 V94 1.3553198157285405e-19

R21_95 V21 V95 5377.177345517726
L21_95 V21 V95 -5.900699849104735e-12
C21_95 V21 V95 4.698650192443038e-20

R21_96 V21 V96 3938.1336976733214
L21_96 V21 V96 -3.786956830921105e-12
C21_96 V21 V96 6.771376092418879e-20

R21_97 V21 V97 611.4070506515877
L21_97 V21 V97 -1.9816343103696686e-12
C21_97 V21 V97 -6.86249805745662e-20

R21_98 V21 V98 -612.9247842362275
L21_98 V21 V98 4.332617679480409e-12
C21_98 V21 V98 1.1050580423940419e-19

R21_99 V21 V99 -642.8854016276946
L21_99 V21 V99 -1.8147448070217992e-12
C21_99 V21 V99 -1.1873550529855358e-19

R21_100 V21 V100 -609.1674227453308
L21_100 V21 V100 -3.237363364767855e-12
C21_100 V21 V100 -3.671556636113729e-20

R21_101 V21 V101 -1973.960117534973
L21_101 V21 V101 1.6026148109299219e-12
C21_101 V21 V101 2.744308796005978e-20

R21_102 V21 V102 -6560.919936785099
L21_102 V21 V102 -2.4714309640709944e-12
C21_102 V21 V102 -1.431486784687167e-19

R21_103 V21 V103 -48619.81450466003
L21_103 V21 V103 5.0075117030528964e-11
C21_103 V21 V103 -3.24861813819447e-20

R21_104 V21 V104 -3346.4760848736637
L21_104 V21 V104 5.7628106942177534e-11
C21_104 V21 V104 -3.6668062633736257e-20

R21_105 V21 V105 283.0998827744617
L21_105 V21 V105 1.3271259668983317e-12
C21_105 V21 V105 -7.216284361098095e-20

R21_106 V21 V106 -3862.9943566782636
L21_106 V21 V106 -1.0808655289572298e-11
C21_106 V21 V106 -2.921028320896199e-20

R21_107 V21 V107 15872.894770645602
L21_107 V21 V107 3.949924679234536e-12
C21_107 V21 V107 9.782806872830936e-20

R21_108 V21 V108 2935.2697799863877
L21_108 V21 V108 4.738744896164737e-12
C21_108 V21 V108 1.388271312425855e-21

R21_109 V21 V109 -2645.2633938228473
L21_109 V21 V109 -2.0762597248116923e-11
C21_109 V21 V109 7.045981803196898e-20

R21_110 V21 V110 38638.22580398529
L21_110 V21 V110 6.624675830229976e-12
C21_110 V21 V110 6.538126047003362e-20

R21_111 V21 V111 -10557.466946473467
L21_111 V21 V111 2.9125609414233023e-12
C21_111 V21 V111 5.935668116539e-20

R21_112 V21 V112 -3956.0794958350416
L21_112 V21 V112 8.161824049764538e-12
C21_112 V21 V112 6.307882481610981e-20

R21_113 V21 V113 1121.716209329127
L21_113 V21 V113 -2.355255870104851e-12
C21_113 V21 V113 1.2335918286979372e-19

R21_114 V21 V114 -4351.3743598568935
L21_114 V21 V114 -9.446122367998425e-12
C21_114 V21 V114 5.768053595388258e-20

R21_115 V21 V115 -2810.074634264547
L21_115 V21 V115 -1.6735506154542697e-12
C21_115 V21 V115 -1.2657952967179598e-19

R21_116 V21 V116 -4297.66444886619
L21_116 V21 V116 -2.080446582232861e-12
C21_116 V21 V116 -3.5021730104076425e-20

R21_117 V21 V117 777.0764045261913
L21_117 V21 V117 -2.2959254156966266e-12
C21_117 V21 V117 -2.0328433943173496e-19

R21_118 V21 V118 -14441.816999293402
L21_118 V21 V118 2.351069235129235e-11
C21_118 V21 V118 -9.356943973451453e-20

R21_119 V21 V119 -3079.9220338625355
L21_119 V21 V119 2.872129046648375e-11
C21_119 V21 V119 -2.3824571862734142e-20

R21_120 V21 V120 -1850.0980123431434
L21_120 V21 V120 -2.430033885372599e-11
C21_120 V21 V120 -8.586015285302907e-20

R21_121 V21 V121 10917.46375507747
L21_121 V21 V121 9.922614142079727e-13
C21_121 V21 V121 1.0763734328688853e-19

R21_122 V21 V122 -3582.6456877998726
L21_122 V21 V122 8.308576371314609e-11
C21_122 V21 V122 1.9107381916831537e-20

R21_123 V21 V123 3618.3278189940556
L21_123 V21 V123 3.934978604762836e-12
C21_123 V21 V123 9.478263749387455e-20

R21_124 V21 V124 2954.0226119649014
L21_124 V21 V124 2.5407223409223514e-12
C21_124 V21 V124 1.099685754838063e-19

R21_125 V21 V125 408.08909755207634
L21_125 V21 V125 1.0468805483405947e-12
C21_125 V21 V125 1.3981451750314833e-19

R21_126 V21 V126 -6264.082468501174
L21_126 V21 V126 4.4361184729007035e-12
C21_126 V21 V126 8.287673151226153e-20

R21_127 V21 V127 -6713.517369230263
L21_127 V21 V127 -1.133572256344168e-11
C21_127 V21 V127 1.0612561379634253e-21

R21_128 V21 V128 4173.853367959192
L21_128 V21 V128 3.720558575681701e-11
C21_128 V21 V128 4.620640938487116e-20

R21_129 V21 V129 -5919.177179973137
L21_129 V21 V129 -1.4839973373184569e-12
C21_129 V21 V129 -1.7909818441570993e-19

R21_130 V21 V130 7124.501399216654
L21_130 V21 V130 -2.6763499860326426e-12
C21_130 V21 V130 -9.733457531533122e-20

R21_131 V21 V131 33266.09332853975
L21_131 V21 V131 -1.0257164762537199e-10
C21_131 V21 V131 -5.1989951220888084e-20

R21_132 V21 V132 -1664.4950450323017
L21_132 V21 V132 -3.287687240879945e-12
C21_132 V21 V132 -1.5053185284566359e-19

R21_133 V21 V133 -714.5524935169466
L21_133 V21 V133 -1.634104647812265e-12
C21_133 V21 V133 7.341480083534172e-20

R21_134 V21 V134 -1153.0710911244093
L21_134 V21 V134 -7.783517491853364e-12
C21_134 V21 V134 6.221648133722236e-20

R21_135 V21 V135 8422.472503438026
L21_135 V21 V135 3.1438997851981375e-10
C21_135 V21 V135 5.993632058847651e-20

R21_136 V21 V136 2228.72377355156
L21_136 V21 V136 1.1051831436056123e-11
C21_136 V21 V136 7.232967687755949e-20

R21_137 V21 V137 538.1576549701189
L21_137 V21 V137 -4.3245467829673806e-12
C21_137 V21 V137 -4.086792347713373e-20

R21_138 V21 V138 834.757920408798
L21_138 V21 V138 2.41380631361789e-12
C21_138 V21 V138 1.5919141714041547e-20

R21_139 V21 V139 -2309.59628692122
L21_139 V21 V139 -2.247483614961716e-11
C21_139 V21 V139 -8.889852481487928e-20

R21_140 V21 V140 -2492.11710437322
L21_140 V21 V140 -5.383660309886618e-12
C21_140 V21 V140 -5.995496749177112e-20

R21_141 V21 V141 -1029.2722711364138
L21_141 V21 V141 9.905690796366318e-13
C21_141 V21 V141 1.0576088368956969e-19

R21_142 V21 V142 -972.8234293092165
L21_142 V21 V142 -5.8498675167262146e-12
C21_142 V21 V142 -3.2188795805349874e-20

R21_143 V21 V143 -2420.0675572733685
L21_143 V21 V143 -5.794871277260496e-12
C21_143 V21 V143 5.0683117304197964e-20

R21_144 V21 V144 -1029.8556471918828
L21_144 V21 V144 1.897483527773778e-10
C21_144 V21 V144 3.1411390266592076e-20

R21_145 V21 V145 367.13766027667566
L21_145 V21 V145 1.1003323442617588e-12
C21_145 V21 V145 1.359461419450545e-19

R21_146 V21 V146 -1907.8653035408972
L21_146 V21 V146 -7.85968291793547e-12
C21_146 V21 V146 -2.0010956139271348e-20

R21_147 V21 V147 4678.831502547894
L21_147 V21 V147 2.2816324661040026e-12
C21_147 V21 V147 1.0119639872503234e-19

R21_148 V21 V148 748.6716229203886
L21_148 V21 V148 1.830967825096432e-12
C21_148 V21 V148 7.070724093301555e-20

R21_149 V21 V149 -256.84890887360973
L21_149 V21 V149 -1.4170403282796138e-12
C21_149 V21 V149 -2.9264099191743334e-19

R21_150 V21 V150 795.7346299308597
L21_150 V21 V150 2.0106899992440153e-12
C21_150 V21 V150 1.0789745127834288e-19

R21_151 V21 V151 831.5662094248828
L21_151 V21 V151 3.0023175558712027e-12
C21_151 V21 V151 -5.951677393876714e-20

R21_152 V21 V152 -1826.1896384003073
L21_152 V21 V152 -1.0655163609784934e-11
C21_152 V21 V152 -1.7719225799961577e-20

R21_153 V21 V153 385.929523178971
L21_153 V21 V153 -9.250877366429288e-13
C21_153 V21 V153 -9.754161604238889e-20

R21_154 V21 V154 -2566.845933008867
L21_154 V21 V154 -2.4307425582595867e-12
C21_154 V21 V154 -8.054741303169843e-20

R21_155 V21 V155 -548.7713974694066
L21_155 V21 V155 -1.7663586464934376e-12
C21_155 V21 V155 -6.359778311706426e-20

R21_156 V21 V156 5171.454292178732
L21_156 V21 V156 -3.470246422192733e-12
C21_156 V21 V156 -7.79702362763055e-20

R21_157 V21 V157 329.1907517351417
L21_157 V21 V157 4.622753091982764e-12
C21_157 V21 V157 2.582021090001004e-19

R21_158 V21 V158 -1579.7446723977932
L21_158 V21 V158 -6.206720017867192e-12
C21_158 V21 V158 -4.770549528440899e-21

R21_159 V21 V159 37006.34615578718
L21_159 V21 V159 -3.1535585120026052e-12
C21_159 V21 V159 -3.51773045266204e-21

R21_160 V21 V160 -970.8927895449555
L21_160 V21 V160 -2.4717835952940668e-12
C21_160 V21 V160 4.8760027357295526e-21

R21_161 V21 V161 2999.837632170369
L21_161 V21 V161 1.1148794789000973e-12
C21_161 V21 V161 3.870263962835357e-20

R21_162 V21 V162 -12728.481692770789
L21_162 V21 V162 -8.160305931104839e-12
C21_162 V21 V162 -6.256551932992745e-20

R21_163 V21 V163 -848.7190003880701
L21_163 V21 V163 -5.012641808352814e-12
C21_163 V21 V163 -1.1595568067972699e-20

R21_164 V21 V164 -9764.02095640195
L21_164 V21 V164 4.4191343854469055e-12
C21_164 V21 V164 -3.397951908051401e-20

R21_165 V21 V165 381.23254937421325
L21_165 V21 V165 7.519267112234391e-13
C21_165 V21 V165 -5.1223545581788414e-20

R21_166 V21 V166 -1417.9064203501598
L21_166 V21 V166 1.458639366123879e-12
C21_166 V21 V166 5.746048488530313e-20

R21_167 V21 V167 3189.9168462511575
L21_167 V21 V167 1.9362677894601686e-12
C21_167 V21 V167 3.7266391856661377e-20

R21_168 V21 V168 -734.2787794951114
L21_168 V21 V168 2.059765071938403e-12
C21_168 V21 V168 8.283963742498376e-20

R21_169 V21 V169 15722.029924692853
L21_169 V21 V169 -9.49907067665778e-13
C21_169 V21 V169 -2.3794028304439707e-20

R21_170 V21 V170 514.513692638447
L21_170 V21 V170 7.616463208419745e-12
C21_170 V21 V170 -3.381190416352945e-20

R21_171 V21 V171 576.3639408975621
L21_171 V21 V171 2.7400203980001448e-12
C21_171 V21 V171 -4.468627533480954e-20

R21_172 V21 V172 698.1676082660284
L21_172 V21 V172 1.0716065960657364e-11
C21_172 V21 V172 -4.245243104807048e-20

R21_173 V21 V173 615.3498505013372
L21_173 V21 V173 -1.532541998735003e-12
C21_173 V21 V173 -1.006067364746116e-20

R21_174 V21 V174 -554.2616423278033
L21_174 V21 V174 -7.190524895923665e-13
C21_174 V21 V174 -2.5788025687735842e-20

R21_175 V21 V175 -519.3346590901494
L21_175 V21 V175 -7.982865382286454e-13
C21_175 V21 V175 -8.792607278679812e-20

R21_176 V21 V176 -644.603656802646
L21_176 V21 V176 -6.67523731825321e-13
C21_176 V21 V176 -9.747419652469767e-20

R21_177 V21 V177 -1628.9366458533582
L21_177 V21 V177 1.4992200463710936e-12
C21_177 V21 V177 -4.640763252140059e-20

R21_178 V21 V178 3382.956434895707
L21_178 V21 V178 4.316037157794106e-12
C21_178 V21 V178 4.4486935029861915e-20

R21_179 V21 V179 -9352.906832555422
L21_179 V21 V179 2.877593645421307e-12
C21_179 V21 V179 1.2456045106363507e-19

R21_180 V21 V180 2488.5668131741045
L21_180 V21 V180 1.6535376824481048e-12
C21_180 V21 V180 1.150516724791648e-19

R21_181 V21 V181 -476.87783327895545
L21_181 V21 V181 1.7676586953355257e-12
C21_181 V21 V181 1.7301533531809166e-19

R21_182 V21 V182 1146.518136377269
L21_182 V21 V182 2.323735133444314e-12
C21_182 V21 V182 -4.0005735885117465e-20

R21_183 V21 V183 1304.3641721747397
L21_183 V21 V183 2.292418956175596e-12
C21_183 V21 V183 7.305069631225416e-21

R21_184 V21 V184 1051.3121156425989
L21_184 V21 V184 1.308462682653403e-12
C21_184 V21 V184 3.3507080360616096e-22

R21_185 V21 V185 216.92252201804982
L21_185 V21 V185 -7.839756493655785e-12
C21_185 V21 V185 -6.647395336847117e-20

R21_186 V21 V186 -780.1258834488399
L21_186 V21 V186 1.2174951273574678e-12
C21_186 V21 V186 2.637018762212034e-20

R21_187 V21 V187 -13088.73340224571
L21_187 V21 V187 7.455822159829443e-12
C21_187 V21 V187 -8.576691797933652e-20

R21_188 V21 V188 -4048.033587574571
L21_188 V21 V188 1.9536501753140562e-11
C21_188 V21 V188 -4.8584058262107934e-20

R21_189 V21 V189 -245.4315525965428
L21_189 V21 V189 -9.63680216058398e-13
C21_189 V21 V189 -8.289893823238077e-20

R21_190 V21 V190 10114.760709650936
L21_190 V21 V190 -2.2713325105198544e-12
C21_190 V21 V190 4.4967256914142726e-20

R21_191 V21 V191 888.0460452453832
L21_191 V21 V191 -2.4400674530677934e-12
C21_191 V21 V191 -1.632924828158839e-20

R21_192 V21 V192 1519.330421607977
L21_192 V21 V192 -1.2166670547578466e-12
C21_192 V21 V192 -3.6926048957277315e-20

R21_193 V21 V193 -3126.343814670188
L21_193 V21 V193 1.9868714633473484e-12
C21_193 V21 V193 4.9583535679857654e-20

R21_194 V21 V194 1101.729960548528
L21_194 V21 V194 -7.922505643950702e-13
C21_194 V21 V194 -3.3659135349204446e-20

R21_195 V21 V195 -4302.476915173451
L21_195 V21 V195 9.53800514512335e-12
C21_195 V21 V195 5.117834157638027e-20

R21_196 V21 V196 -3900.140795681506
L21_196 V21 V196 -2.8500601063327354e-12
C21_196 V21 V196 2.2301292269092892e-20

R21_197 V21 V197 474.08495173667814
L21_197 V21 V197 2.0177957312791015e-12
C21_197 V21 V197 1.8430446390206518e-20

R21_198 V21 V198 -1331.4789894767916
L21_198 V21 V198 1.7500943684662546e-12
C21_198 V21 V198 -1.6302272318960273e-20

R21_199 V21 V199 -718.0843788965793
L21_199 V21 V199 2.7944061657357292e-12
C21_199 V21 V199 -1.4954270718062094e-20

R21_200 V21 V200 -795.2408270769921
L21_200 V21 V200 9.561221736624296e-13
C21_200 V21 V200 3.409388241044031e-20

R22_22 V22 0 -120.76590120969006
L22_22 V22 0 -2.9012991332148693e-13
C22_22 V22 0 -3.456673205152099e-19

R22_23 V22 V23 -2777.7296468979584
L22_23 V22 V23 -3.0175666490447543e-12
C22_23 V22 V23 -1.0061217421753774e-19

R22_24 V22 V24 -2466.281675127059
L22_24 V22 V24 -2.4754170526419324e-12
C22_24 V22 V24 -1.2182501387254747e-19

R22_25 V22 V25 1000.5997336068407
L22_25 V22 V25 2.6618482492806043e-12
C22_25 V22 V25 -1.142351615255285e-19

R22_26 V22 V26 1054.2436429072527
L22_26 V22 V26 1.6137164959775993e-12
C22_26 V22 V26 1.630955512671302e-19

R22_27 V22 V27 4594.642502231246
L22_27 V22 V27 4.870966875259135e-12
C22_27 V22 V27 6.885473813653678e-23

R22_28 V22 V28 3658.354685037227
L22_28 V22 V28 3.929990364690065e-12
C22_28 V22 V28 -2.384901086497728e-20

R22_29 V22 V29 1176.1905411764694
L22_29 V22 V29 5.783361997143822e-12
C22_29 V22 V29 -4.6404092746218053e-20

R22_30 V22 V30 872.4716744081081
L22_30 V22 V30 1.01717396823088e-12
C22_30 V22 V30 4.1880853025031256e-19

R22_31 V22 V31 2020.016137687428
L22_31 V22 V31 7.872154757649707e-12
C22_31 V22 V31 4.088615585782917e-20

R22_32 V22 V32 1696.1686667442307
L22_32 V22 V32 8.79324218736354e-12
C22_32 V22 V32 2.6728905762345014e-20

R22_33 V22 V33 2780.225748801049
L22_33 V22 V33 2.3300302949457525e-12
C22_33 V22 V33 1.5038515252434954e-19

R22_34 V22 V34 -3295.2053226358194
L22_34 V22 V34 -1.7017348346159355e-12
C22_34 V22 V34 -4.557883728746161e-19

R22_35 V22 V35 -3156.2984698501973
L22_35 V22 V35 1.9198522318291702e-11
C22_35 V22 V35 5.232993445528008e-20

R22_36 V22 V36 -1919.0000947407034
L22_36 V22 V36 3.0953818235533883e-11
C22_36 V22 V36 6.658998555783448e-20

R22_37 V22 V37 -3212.4169710661527
L22_37 V22 V37 -3.1140348697264007e-12
C22_37 V22 V37 3.770982125162178e-20

R22_38 V22 V38 -2470.947856620777
L22_38 V22 V38 -1.4235957989925238e-12
C22_38 V22 V38 -1.567854275754139e-19

R22_39 V22 V39 -2391.646747788563
L22_39 V22 V39 -5.516827872832711e-12
C22_39 V22 V39 -4.6912480117624126e-20

R22_40 V22 V40 -1723.8244641957435
L22_40 V22 V40 -4.295816488764556e-12
C22_40 V22 V40 -4.6347534552518946e-20

R22_41 V22 V41 32263.84598977232
L22_41 V22 V41 -3.6237454000510885e-12
C22_41 V22 V41 -1.0665219112916647e-19

R22_42 V22 V42 -2319.708719854778
L22_42 V22 V42 3.2604884796244985e-12
C22_42 V22 V42 2.0698238108949276e-19

R22_43 V22 V43 -8416.22464479947
L22_43 V22 V43 -8.716576580864577e-12
C22_43 V22 V43 3.4553821954052086e-21

R22_44 V22 V44 -9388.814243840296
L22_44 V22 V44 -5.512373372897224e-12
C22_44 V22 V44 -2.351593487129987e-20

R22_45 V22 V45 1982.767157916794
L22_45 V22 V45 5.664941341352406e-12
C22_45 V22 V45 -5.770502739709024e-20

R22_46 V22 V46 2001.9674478564032
L22_46 V22 V46 1.7011061755426778e-12
C22_46 V22 V46 3.9614703996090387e-19

R22_47 V22 V47 4156.059729313375
L22_47 V22 V47 -7.348020771302418e-10
C22_47 V22 V47 5.395473950086066e-21

R22_48 V22 V48 2370.120401865209
L22_48 V22 V48 2.253076614471685e-11
C22_48 V22 V48 -3.12261074741064e-21

R22_49 V22 V49 2576.1738582412104
L22_49 V22 V49 4.3953295470226354e-12
C22_49 V22 V49 3.2960716871488427e-20

R22_50 V22 V50 2788.3329004833477
L22_50 V22 V50 -5.265967240013314e-12
C22_50 V22 V50 -2.718249414941629e-19

R22_51 V22 V51 11027.117679810644
L22_51 V22 V51 1.1741425494996845e-11
C22_51 V22 V51 -9.872274458252126e-20

R22_52 V22 V52 -12773.546909373052
L22_52 V22 V52 2.060055188602853e-11
C22_52 V22 V52 -1.174746239878023e-19

R22_53 V22 V53 2575.5100742196028
L22_53 V22 V53 1.9769000807263806e-12
C22_53 V22 V53 1.8149547599057533e-19

R22_54 V22 V54 -16599.532462328778
L22_54 V22 V54 -1.361577494491907e-12
C22_54 V22 V54 -3.6083337298638696e-19

R22_55 V22 V55 -34529.42480644592
L22_55 V22 V55 4.7637084634364085e-12
C22_55 V22 V55 1.3090965686433375e-19

R22_56 V22 V56 -3399.1519985890686
L22_56 V22 V56 5.415523893760678e-12
C22_56 V22 V56 1.4354951761995955e-19

R22_57 V22 V57 56399.22187088645
L22_57 V22 V57 -1.6200686782749688e-12
C22_57 V22 V57 -9.40467008406848e-20

R22_58 V22 V58 20517.099518512132
L22_58 V22 V58 1.2779716826195276e-12
C22_58 V22 V58 4.794933504344849e-19

R22_59 V22 V59 -3343.9543769267398
L22_59 V22 V59 -7.576398238808954e-12
C22_59 V22 V59 5.99253203103117e-20

R22_60 V22 V60 -2355.1666894419204
L22_60 V22 V60 -4.7587572285757675e-12
C22_60 V22 V60 8.872175271099953e-20

R22_61 V22 V61 -10266.644918416448
L22_61 V22 V61 -2.04628869011784e-10
C22_61 V22 V61 -1.2499908081166679e-19

R22_62 V22 V62 -2721.6304283844374
L22_62 V22 V62 5.6751087484593354e-12
C22_62 V22 V62 3.518016236330077e-20

R22_63 V22 V63 48589.91729601762
L22_63 V22 V63 -3.4513903877531856e-12
C22_63 V22 V63 -1.557639462109527e-19

R22_64 V22 V64 6129.375583763839
L22_64 V22 V64 -3.217929413477581e-12
C22_64 V22 V64 -2.2748025414300513e-19

R22_65 V22 V65 2738.8225532094716
L22_65 V22 V65 2.52130872389733e-12
C22_65 V22 V65 1.6807235163140879e-19

R22_66 V22 V66 2730.926623497733
L22_66 V22 V66 -1.920771005925481e-12
C22_66 V22 V66 -2.401029947989498e-19

R22_67 V22 V67 24942.288887713916
L22_67 V22 V67 5.9062834061978685e-12
C22_67 V22 V67 5.676527282945297e-20

R22_68 V22 V68 5335.288240654009
L22_68 V22 V68 3.340600591476078e-12
C22_68 V22 V68 7.393519785717816e-20

R22_69 V22 V69 5341.325197310517
L22_69 V22 V69 5.708744147248764e-12
C22_69 V22 V69 -2.937270631187488e-20

R22_70 V22 V70 3678.1747252325304
L22_70 V22 V70 1.7650704474682765e-12
C22_70 V22 V70 1.6616935869458413e-19

R22_71 V22 V71 7017.033583982855
L22_71 V22 V71 4.974397743768555e-12
C22_71 V22 V71 5.098136814080554e-20

R22_72 V22 V72 6834.39259093408
L22_72 V22 V72 3.5483539471999433e-12
C22_72 V22 V72 1.1656741265945072e-19

R22_73 V22 V73 2545.842543453286
L22_73 V22 V73 -2.448969761850591e-11
C22_73 V22 V73 -9.791696912713005e-20

R22_74 V22 V74 -2600.6762374691643
L22_74 V22 V74 7.374135502479389e-12
C22_74 V22 V74 -6.784083117725697e-21

R22_75 V22 V75 -26532.566885806038
L22_75 V22 V75 -5.130532016213946e-12
C22_75 V22 V75 -7.325077531420038e-20

R22_76 V22 V76 -2285.7225979241894
L22_76 V22 V76 -2.8554642369703205e-12
C22_76 V22 V76 -1.4143740560242617e-19

R22_77 V22 V77 -4949.144271994512
L22_77 V22 V77 -4.0638520558654625e-12
C22_77 V22 V77 1.1108945774363503e-19

R22_78 V22 V78 2367.0666139775053
L22_78 V22 V78 -3.2926946984219826e-12
C22_78 V22 V78 -8.65222421591741e-21

R22_79 V22 V79 -4738.717211255931
L22_79 V22 V79 -2.6430969967124925e-11
C22_79 V22 V79 1.97773416561352e-20

R22_80 V22 V80 -67919.38518187744
L22_80 V22 V80 -4.46303785478996e-11
C22_80 V22 V80 4.272137055128527e-20

R22_81 V22 V81 1226.6861377357488
L22_81 V22 V81 2.719036379171646e-12
C22_81 V22 V81 2.2449960529407097e-20

R22_82 V22 V82 -5993.338268280081
L22_82 V22 V82 5.92442285307713e-12
C22_82 V22 V82 6.063976272943102e-20

R22_83 V22 V83 -7384.60213693979
L22_83 V22 V83 1.8961292805364788e-11
C22_83 V22 V83 5.974881243249424e-20

R22_84 V22 V84 -16854.841154688027
L22_84 V22 V84 1.4570682066223085e-11
C22_84 V22 V84 8.602991629924856e-20

R22_85 V22 V85 -6932.893933119997
L22_85 V22 V85 2.9000169530816783e-10
C22_85 V22 V85 -7.241514985734047e-20

R22_86 V22 V86 16018.853154748436
L22_86 V22 V86 7.769879617325574e-12
C22_86 V22 V86 -1.1957618467958417e-19

R22_87 V22 V87 11860.864701931798
L22_87 V22 V87 -1.155853406091879e-11
C22_87 V22 V87 -4.173074437129834e-20

R22_88 V22 V88 21373.70484461189
L22_88 V22 V88 -1.3739598761540685e-11
C22_88 V22 V88 -7.625514288626901e-20

R22_89 V22 V89 7103.7929772006255
L22_89 V22 V89 5.367924456487236e-12
C22_89 V22 V89 -3.7814310187542684e-20

R22_90 V22 V90 8042.936343628383
L22_90 V22 V90 3.829131694903335e-11
C22_90 V22 V90 4.6335261199190574e-20

R22_91 V22 V91 7013.053048214312
L22_91 V22 V91 5.489565125747286e-12
C22_91 V22 V91 1.4082413788733703e-20

R22_92 V22 V92 -6947.712938714409
L22_92 V22 V92 5.231899003271892e-12
C22_92 V22 V92 2.3558337044488443e-20

R22_93 V22 V93 1678.646762443582
L22_93 V22 V93 -9.466235128516293e-12
C22_93 V22 V93 6.887118664707179e-20

R22_94 V22 V94 -1879.6181498219012
L22_94 V22 V94 -6.276399027832603e-12
C22_94 V22 V94 1.0059876837453408e-19

R22_95 V22 V95 -3311.50740705217
L22_95 V22 V95 -1.1531219391582708e-11
C22_95 V22 V95 3.632386472932707e-21

R22_96 V22 V96 -2617.636110249413
L22_96 V22 V96 -6.8424035973357285e-12
C22_96 V22 V96 1.3104969885252618e-20

R22_97 V22 V97 -10144.743304432794
L22_97 V22 V97 -5.402232843437207e-12
C22_97 V22 V97 7.523864577770584e-20

R22_98 V22 V98 2471.8271798654678
L22_98 V22 V98 2.7174621787859e-12
C22_98 V22 V98 -1.2645648847537927e-20

R22_99 V22 V99 -2513.6099608061154
L22_99 V22 V99 -5.363038430226443e-12
C22_99 V22 V99 1.1681801698303336e-20

R22_100 V22 V100 -9715.620192235501
L22_100 V22 V100 -3.706806141114036e-12
C22_100 V22 V100 -3.0927166935834086e-21

R22_101 V22 V101 11411.39457943363
L22_101 V22 V101 3.745065332322838e-12
C22_101 V22 V101 -7.641235160542911e-20

R22_102 V22 V102 72521.45140178966
L22_102 V22 V102 -2.283913061613863e-12
C22_102 V22 V102 -1.9261489236970087e-19

R22_103 V22 V103 3664.3213651984393
L22_103 V22 V103 5.5196359131796235e-12
C22_103 V22 V103 -1.0300245206307778e-22

R22_104 V22 V104 4763.422679330024
L22_104 V22 V104 4.287299802783503e-12
C22_104 V22 V104 2.3558012144928072e-20

R22_105 V22 V105 964.0768972912292
L22_105 V22 V105 3.469609306038749e-12
C22_105 V22 V105 -4.912337451141498e-20

R22_106 V22 V106 2890.5198922808263
L22_106 V22 V106 8.001489486461952e-12
C22_106 V22 V106 9.694564504972053e-20

R22_107 V22 V107 9967.771843315142
L22_107 V22 V107 -9.24797512001342e-12
C22_107 V22 V107 -3.3358019488443255e-20

R22_108 V22 V108 -8082.52683356105
L22_108 V22 V108 -2.946580079792873e-11
C22_108 V22 V108 -6.110625994803362e-20

R22_109 V22 V109 -2634.4891096469014
L22_109 V22 V109 -5.8649463300812294e-12
C22_109 V22 V109 5.226409326474e-20

R22_110 V22 V110 -1631.3822722397608
L22_110 V22 V110 1.9983777434278664e-12
C22_110 V22 V110 2.9048225503624167e-19

R22_111 V22 V111 5678.719919614242
L22_111 V22 V111 -1.713996481094247e-11
C22_111 V22 V111 -9.643924032876046e-21

R22_112 V22 V112 7706.751037176479
L22_112 V22 V112 -7.618902380816552e-12
C22_112 V22 V112 -1.1587976539645867e-20

R22_113 V22 V113 3002.616875833405
L22_113 V22 V113 -4.452340241655885e-12
C22_113 V22 V113 7.132657139262445e-20

R22_114 V22 V114 -2758.6266584606788
L22_114 V22 V114 -1.5570887000533251e-12
C22_114 V22 V114 -3.1103917427135204e-19

R22_115 V22 V115 -1470.4907609010468
L22_115 V22 V115 2.3633379400177788e-11
C22_115 V22 V115 2.0128630002271436e-20

R22_116 V22 V116 -2571.414984410204
L22_116 V22 V116 -2.2129946260259688e-11
C22_116 V22 V116 5.840107021802967e-20

R22_117 V22 V117 -15338.625226502108
L22_117 V22 V117 1.9371888303338043e-11
C22_117 V22 V117 -2.750602624855368e-20

R22_118 V22 V118 1248.8337363684475
L22_118 V22 V118 1.3112911187638753e-11
C22_118 V22 V118 -9.270237668871865e-20

R22_119 V22 V119 3528.652622317349
L22_119 V22 V119 1.3983459755075035e-10
C22_119 V22 V119 -1.0017974292622169e-20

R22_120 V22 V120 4713.9608419992155
L22_120 V22 V120 6.387089589197204e-11
C22_120 V22 V120 -2.759855196787391e-20

R22_121 V22 V121 3609.9523889790353
L22_121 V22 V121 3.0075046743924432e-12
C22_121 V22 V121 -8.115571673804253e-20

R22_122 V22 V122 35997.013032737326
L22_122 V22 V122 6.121000609160268e-12
C22_122 V22 V122 2.747752797110148e-19

R22_123 V22 V123 2061.8101394046034
L22_123 V22 V123 -2.402826577108049e-11
C22_123 V22 V123 -3.5853716202203714e-20

R22_124 V22 V124 2443.045001316018
L22_124 V22 V124 4.251506558367525e-11
C22_124 V22 V124 -4.4607412268592515e-20

R22_125 V22 V125 888.085683198577
L22_125 V22 V125 1.2899899166390024e-11
C22_125 V22 V125 4.686794088870217e-20

R22_126 V22 V126 11961.86263956517
L22_126 V22 V126 -4.156884471886299e-11
C22_126 V22 V126 -1.189454024468002e-19

R22_127 V22 V127 -1857.6809972908284
L22_127 V22 V127 -2.0417728071361362e-11
C22_127 V22 V127 1.2407120588320306e-20

R22_128 V22 V128 -2147.051123080068
L22_128 V22 V128 -1.675358801622696e-11
C22_128 V22 V128 1.6451186289976617e-20

R22_129 V22 V129 -1176.6877694979694
L22_129 V22 V129 -4.33944234944544e-12
C22_129 V22 V129 2.9950952612488705e-20

R22_130 V22 V130 -1354.211047235788
L22_130 V22 V130 3.044987027962631e-11
C22_130 V22 V130 -5.692866529936815e-20

R22_131 V22 V131 3315.137321803454
L22_131 V22 V131 1.0736456744680269e-11
C22_131 V22 V131 2.8009317435401305e-20

R22_132 V22 V132 4343.42094410397
L22_132 V22 V132 7.698256084890808e-12
C22_132 V22 V132 4.3485811000951566e-20

R22_133 V22 V133 -1846.3490323052383
L22_133 V22 V133 7.844500538063014e-12
C22_133 V22 V133 -2.528192897141185e-20

R22_134 V22 V134 1938.2185068290062
L22_134 V22 V134 -2.383491863626295e-12
C22_134 V22 V134 7.934021580184237e-20

R22_135 V22 V135 4992.190488779
L22_135 V22 V135 -1.8803709232948715e-11
C22_135 V22 V135 -3.217683538337906e-20

R22_136 V22 V136 2486.4143058258223
L22_136 V22 V136 -2.2069374789136784e-11
C22_136 V22 V136 -1.72400050308637e-21

R22_137 V22 V137 670.994652064347
L22_137 V22 V137 -3.4852328585293324e-12
C22_137 V22 V137 5.718889435816575e-21

R22_138 V22 V138 2731.141293235278
L22_138 V22 V138 3.4775682828901648e-12
C22_138 V22 V138 -3.2071287365213563e-20

R22_139 V22 V139 -2038.8537779576195
L22_139 V22 V139 -8.819212542314061e-11
C22_139 V22 V139 -4.462086337366596e-21

R22_140 V22 V140 -10153.714796833505
L22_140 V22 V140 -6.499647747561123e-12
C22_140 V22 V140 -4.9440165457387284e-20

R22_141 V22 V141 -5096.3605554090755
L22_141 V22 V141 1.1031959086010732e-11
C22_141 V22 V141 1.0125015729839291e-20

R22_142 V22 V142 -700.6803646780529
L22_142 V22 V142 1.4121296677899714e-12
C22_142 V22 V142 4.408540142926375e-20

R22_143 V22 V143 3585.4663973618194
L22_143 V22 V143 -4.047806515799847e-11
C22_143 V22 V143 3.6182163866138776e-20

R22_144 V22 V144 -1105.7837208949836
L22_144 V22 V144 7.527439016657415e-12
C22_144 V22 V144 2.4485686440365533e-20

R22_145 V22 V145 -1942.7485395017125
L22_145 V22 V145 1.3890418313333204e-12
C22_145 V22 V145 -4.9731045061355244e-21

R22_146 V22 V146 1062.9116382082614
L22_146 V22 V146 -2.690598303337623e-12
C22_146 V22 V146 -6.904383812253419e-20

R22_147 V22 V147 -1139.3030234770677
L22_147 V22 V147 7.118175715009363e-12
C22_147 V22 V147 -2.8829273180414264e-20

R22_148 V22 V148 622.1942869255737
L22_148 V22 V148 4.975227149280497e-12
C22_148 V22 V148 9.158139337959614e-21

R22_149 V22 V149 -1418.8625876681754
L22_149 V22 V149 -7.767852361256518e-12
C22_149 V22 V149 -2.0985101923323663e-20

R22_150 V22 V150 1175.8931442769679
L22_150 V22 V150 -1.4283539291109347e-12
C22_150 V22 V150 1.074415571629803e-20

R22_151 V22 V151 748.9635020406313
L22_151 V22 V151 4.362174720592098e-12
C22_151 V22 V151 -7.938411174891265e-21

R22_152 V22 V152 -770.4690095058277
L22_152 V22 V152 2.754615267608032e-11
C22_152 V22 V152 -8.550739700085512e-21

R22_153 V22 V153 664.0446635838894
L22_153 V22 V153 -1.530713769890121e-12
C22_153 V22 V153 2.3188613750454554e-20

R22_154 V22 V154 55304.33655451482
L22_154 V22 V154 -6.764699268837487e-11
C22_154 V22 V154 2.2239585446376937e-20

R22_155 V22 V155 -367.9641581500397
L22_155 V22 V155 -7.814847389251985e-12
C22_155 V22 V155 3.283846774388119e-22

R22_156 V22 V156 529.0137074265759
L22_156 V22 V156 -9.342710117571566e-12
C22_156 V22 V156 1.3350106448697308e-20

R22_157 V22 V157 1292.0302321748652
L22_157 V22 V157 -1.469084004914031e-11
C22_157 V22 V157 4.53328365635507e-20

R22_158 V22 V158 -2097.1430618980603
L22_158 V22 V158 7.493209511403202e-13
C22_158 V22 V158 4.4644207650381553e-20

R22_159 V22 V159 530.6034496344782
L22_159 V22 V159 -3.2058844929431847e-12
C22_159 V22 V159 3.1051879095920115e-21

R22_160 V22 V160 -1271.2319244601574
L22_160 V22 V160 -3.0832202705473668e-12
C22_160 V22 V160 -1.60051506151364e-20

R22_161 V22 V161 -1801.2972746270816
L22_161 V22 V161 2.5796154556728835e-12
C22_161 V22 V161 -4.900616570067064e-20

R22_162 V22 V162 -3472.841996401216
L22_162 V22 V162 -3.949695317133149e-12
C22_162 V22 V162 -5.859572817596185e-20

R22_163 V22 V163 -2985.89458201225
L22_163 V22 V163 -1.1904439139645346e-11
C22_163 V22 V163 1.5899503944325126e-20

R22_164 V22 V164 1221.2686527901171
L22_164 V22 V164 6.099120038664709e-12
C22_164 V22 V164 -1.1855644708269976e-20

R22_165 V22 V165 924.4361071648029
L22_165 V22 V165 1.5381643880272651e-12
C22_165 V22 V165 2.609676378523648e-21

R22_166 V22 V166 630.9414359700717
L22_166 V22 V166 -7.834573320446506e-13
C22_166 V22 V166 -7.823759064841397e-21

R22_167 V22 V167 2987.2555713082484
L22_167 V22 V167 1.6468214865472011e-12
C22_167 V22 V167 2.1685950478069026e-21

R22_168 V22 V168 -506.8256248685498
L22_168 V22 V168 1.6842111733415792e-12
C22_168 V22 V168 7.533198625202218e-21

R22_169 V22 V169 1961.423505602395
L22_169 V22 V169 -2.165629289639615e-12
C22_169 V22 V169 7.334909144288732e-21

R22_170 V22 V170 -2435.5413970109826
L22_170 V22 V170 7.8928452233798e-13
C22_170 V22 V170 1.1010511509402274e-20

R22_171 V22 V171 -2419.507524864112
L22_171 V22 V171 7.387606015187576e-12
C22_171 V22 V171 -4.651862832595393e-20

R22_172 V22 V172 1640.820581811539
L22_172 V22 V172 -1.2351027579919958e-11
C22_172 V22 V172 -1.542734563968285e-20

R22_173 V22 V173 5529.214886870631
L22_173 V22 V173 -1.1240004046713311e-11
C22_173 V22 V173 3.014411215325049e-20

R22_174 V22 V174 -430.6087039896637
L22_174 V22 V174 4.624167762428663e-12
C22_174 V22 V174 -1.8395934592185093e-21

R22_175 V22 V175 7029.421332165656
L22_175 V22 V175 -1.5951528741277083e-12
C22_175 V22 V175 1.8642802014021515e-20

R22_176 V22 V176 2008.0423670781365
L22_176 V22 V176 -1.236004384995837e-12
C22_176 V22 V176 5.321092439182072e-21

R22_177 V22 V177 1802.7731534112545
L22_177 V22 V177 2.6783809605945255e-12
C22_177 V22 V177 -3.65738913783187e-20

R22_178 V22 V178 608.7766532371688
L22_178 V22 V178 -1.075930477540277e-12
C22_178 V22 V178 4.609010746559534e-20

R22_179 V22 V179 -2125.465746311745
L22_179 V22 V179 3.769907696564691e-12
C22_179 V22 V179 3.2990718525501405e-20

R22_180 V22 V180 -71619.10960005662
L22_180 V22 V180 1.8738363488201564e-12
C22_180 V22 V180 1.9936457358402033e-20

R22_181 V22 V181 -1055.1759736462736
L22_181 V22 V181 -8.259931901802037e-12
C22_181 V22 V181 -2.7404310794784714e-21

R22_182 V22 V182 14299.913621252143
L22_182 V22 V182 3.010109359739496e-12
C22_182 V22 V182 -3.243193685278077e-20

R22_183 V22 V183 1011.3999946837524
L22_183 V22 V183 7.799853902314013e-12
C22_183 V22 V183 1.5480088567806227e-20

R22_184 V22 V184 2482.892328472938
L22_184 V22 V184 4.1078856083459e-12
C22_184 V22 V184 -1.2114807050261137e-21

R22_185 V22 V185 1199.4244514897132
L22_185 V22 V185 7.68795078146578e-12
C22_185 V22 V185 3.8526810685475007e-20

R22_186 V22 V186 -851.7211523474858
L22_186 V22 V186 2.9658958990625384e-12
C22_186 V22 V186 -6.522833352523577e-20

R22_187 V22 V187 -2156.092086933363
L22_187 V22 V187 1.4769930930347173e-11
C22_187 V22 V187 -3.5790191779360926e-20

R22_188 V22 V188 -779.0118610243451
L22_188 V22 V188 -6.583223357046493e-11
C22_188 V22 V188 -1.9759423823818284e-20

R22_189 V22 V189 -7793.048068514954
L22_189 V22 V189 -1.3176771027281028e-11
C22_189 V22 V189 -3.6195374787887127e-20

R22_190 V22 V190 1660.2506522960166
L22_190 V22 V190 -2.3040380453423843e-11
C22_190 V22 V190 7.036398271604743e-20

R22_191 V22 V191 -3764.0077362519432
L22_191 V22 V191 7.704088245323337e-12
C22_191 V22 V191 -3.180008143096881e-20

R22_192 V22 V192 2173.4956588044192
L22_192 V22 V192 -3.7828389574517714e-11
C22_192 V22 V192 -2.0268543670012603e-20

R22_193 V22 V193 -1673.2222890640423
L22_193 V22 V193 -7.873801104430205e-12
C22_193 V22 V193 2.5219525563201815e-20

R22_194 V22 V194 103481.60173409777
L22_194 V22 V194 -3.656823107008924e-12
C22_194 V22 V194 -6.4586887008269035e-21

R22_195 V22 V195 1451.834563502256
L22_195 V22 V195 -5.436270341989821e-12
C22_195 V22 V195 6.243596802352826e-20

R22_196 V22 V196 995.183942513414
L22_196 V22 V196 -2.701802917507546e-12
C22_196 V22 V196 5.460105122512427e-20

R22_197 V22 V197 3380.4509946534417
L22_197 V22 V197 6.888654477510026e-12
C22_197 V22 V197 -4.833209895146168e-21

R22_198 V22 V198 -3272.955359814472
L22_198 V22 V198 -3.6144743170985795e-11
C22_198 V22 V198 1.7879278677792526e-21

R22_199 V22 V199 4323.831378291755
L22_199 V22 V199 -5.891786663783632e-11
C22_199 V22 V199 4.378704032055385e-20

R22_200 V22 V200 -1015.4657231559944
L22_200 V22 V200 3.3934585828311733e-12
C22_200 V22 V200 5.8032726622371245e-21

R23_23 V23 0 -266.91035951070864
L23_23 V23 0 -3.275146266032805e-13
C23_23 V23 0 -5.554074669240575e-19

R23_24 V23 V24 -3011.929857892638
L23_24 V23 V24 -1.5373560389693868e-12
C23_24 V23 V24 -2.944399992424588e-19

R23_25 V23 V25 1711.9228418608366
L23_25 V23 V25 4.070348969849827e-12
C23_25 V23 V25 -1.1265549598442436e-19

R23_26 V23 V26 3851.1837102092063
L23_26 V23 V26 -1.5225683380964136e-11
C23_26 V23 V26 -1.368135114196957e-19

R23_27 V23 V27 1705.0788715203494
L23_27 V23 V27 1.1063771124587073e-12
C23_27 V23 V27 3.3624164247566254e-19

R23_28 V23 V28 3823.455187512121
L23_28 V23 V28 2.7123217783838805e-12
C23_28 V23 V28 2.90061050598883e-20

R23_29 V23 V29 1948.6849245970145
L23_29 V23 V29 2.512039058000562e-12
C23_29 V23 V29 7.565008942840923e-20

R23_30 V23 V30 5182.161112202354
L23_30 V23 V30 3.5984697759298346e-12
C23_30 V23 V30 1.30046778482681e-19

R23_31 V23 V31 1347.603727731476
L23_31 V23 V31 1.1256785977376714e-12
C23_31 V23 V31 4.537217536137693e-19

R23_32 V23 V32 2744.9906002833995
L23_32 V23 V32 3.1180125027373993e-12
C23_32 V23 V32 9.464285477724125e-20

R23_33 V23 V33 5507.947990245435
L23_33 V23 V33 1.0207408226880991e-11
C23_33 V23 V33 2.8361252380995574e-20

R23_34 V23 V34 -12006.717427654574
L23_34 V23 V34 8.104938963186677e-12
C23_34 V23 V34 1.0056733380003339e-19

R23_35 V23 V35 -3212.7794281699266
L23_35 V23 V35 -8.762761066455029e-13
C23_35 V23 V35 -7.875126550770088e-19

R23_36 V23 V36 -3109.3914442410405
L23_36 V23 V36 -5.0116382687980935e-12
C23_36 V23 V36 -1.00102446284718e-19

R23_37 V23 V37 -4853.1572871027
L23_37 V23 V37 -2.4055404676174645e-12
C23_37 V23 V37 -4.8161625609767883e-20

R23_38 V23 V38 -10214.988975225408
L23_38 V23 V38 -2.13709856681152e-12
C23_38 V23 V38 -2.263675711652444e-19

R23_39 V23 V39 -2203.678351996852
L23_39 V23 V39 -4.1556906483203835e-12
C23_39 V23 V39 1.7880806976434638e-19

R23_40 V23 V40 -2608.207844310276
L23_40 V23 V40 -4.834392157867214e-12
C23_40 V23 V40 4.627861199247782e-20

R23_41 V23 V41 167363.75590658392
L23_41 V23 V41 -1.1459305398723812e-11
C23_41 V23 V41 -3.779184813951212e-22

R23_42 V23 V42 351920.5645590528
L23_42 V23 V42 -4.898630823646532e-11
C23_42 V23 V42 5.521350486123629e-20

R23_43 V23 V43 -3333.6813477140417
L23_43 V23 V43 7.319306427829006e-12
C23_43 V23 V43 1.2589981371913877e-19

R23_44 V23 V44 -10910.134242394393
L23_44 V23 V44 -7.52680763571412e-12
C23_44 V23 V44 -4.879466094393601e-20

R23_45 V23 V45 3284.2872925333986
L23_45 V23 V45 4.146071970923327e-12
C23_45 V23 V45 -3.231818412626438e-20

R23_46 V23 V46 6515.736855903477
L23_46 V23 V46 2.634496503969195e-12
C23_46 V23 V46 2.1377946039930186e-19

R23_47 V23 V47 2940.871051765003
L23_47 V23 V47 1.7523308231931501e-12
C23_47 V23 V47 1.1745476159147485e-19

R23_48 V23 V48 3539.4081210880095
L23_48 V23 V48 3.4742708940518008e-12
C23_48 V23 V48 6.185250343060338e-20

R23_49 V23 V49 4295.675482761553
L23_49 V23 V49 4.9621323060856305e-12
C23_49 V23 V49 6.988858872663812e-20

R23_50 V23 V50 19518.635263334265
L23_50 V23 V50 -6.444953869480145e-12
C23_50 V23 V50 -1.862103636322921e-19

R23_51 V23 V51 3420.6532311286787
L23_51 V23 V51 6.8089335167208286e-12
C23_51 V23 V51 1.8068708502663588e-19

R23_52 V23 V52 -207850.4541375071
L23_52 V23 V52 2.601459600253679e-10
C23_52 V23 V52 -5.538212496461202e-20

R23_53 V23 V53 4183.222873931258
L23_53 V23 V53 3.2085052572130668e-12
C23_53 V23 V53 1.053778390347596e-19

R23_54 V23 V54 65442.86100036051
L23_54 V23 V54 3.0530584361561826e-11
C23_54 V23 V54 3.4925919996875933e-20

R23_55 V23 V55 10364.089175759478
L23_55 V23 V55 -1.0683954861241012e-12
C23_55 V23 V55 -5.697838643193763e-19

R23_56 V23 V56 -7433.882625878379
L23_56 V23 V56 -6.258573081054337e-11
C23_56 V23 V56 7.294257620212988e-21

R23_57 V23 V57 -61340.859114890925
L23_57 V23 V57 -1.6126186166594162e-12
C23_57 V23 V57 -1.5569511375569225e-19

R23_58 V23 V58 13515.927946207046
L23_58 V23 V58 -1.0047346749681103e-09
C23_58 V23 V58 4.4346330600961324e-20

R23_59 V23 V59 -1968.9331258426716
L23_59 V23 V59 4.202764791157595e-12
C23_59 V23 V59 1.644140543201714e-19

R23_60 V23 V60 -3096.5740295000237
L23_60 V23 V60 -5.879609089644936e-12
C23_60 V23 V60 2.3351213312324703e-20

R23_61 V23 V61 -19366.852260813408
L23_61 V23 V61 5.9061488709392714e-12
C23_61 V23 V61 2.551857835704443e-20

R23_62 V23 V62 -7382.616299561719
L23_62 V23 V62 -6.224948493528867e-12
C23_62 V23 V62 -5.319726054687426e-20

R23_63 V23 V63 11243.779997094127
L23_63 V23 V63 1.5764960303456997e-12
C23_63 V23 V63 4.481099240379294e-19

R23_64 V23 V64 9742.48662106964
L23_64 V23 V64 -6.520321257956443e-12
C23_64 V23 V64 -9.424549996891241e-20

R23_65 V23 V65 5483.825059798628
L23_65 V23 V65 2.8206190671618054e-12
C23_65 V23 V65 1.5240084963827333e-19

R23_66 V23 V66 10943.600076686233
L23_66 V23 V66 6.252743284462184e-12
C23_66 V23 V66 6.0904115844776e-20

R23_67 V23 V67 9341.129671294228
L23_67 V23 V67 -1.8925823489951942e-12
C23_67 V23 V67 -2.640992509365399e-19

R23_68 V23 V68 7363.066682515721
L23_68 V23 V68 3.803216799086842e-12
C23_68 V23 V68 5.738806063959478e-20

R23_69 V23 V69 5251.09270371391
L23_69 V23 V69 -1.1733809841344524e-11
C23_69 V23 V69 -1.4891181043204716e-19

R23_70 V23 V70 21918.90348671875
L23_70 V23 V70 8.519291031270233e-12
C23_70 V23 V70 1.3509790499665291e-20

R23_71 V23 V71 3819.463460473941
L23_71 V23 V71 4.748952738444253e-12
C23_71 V23 V71 -1.0027020579663643e-19

R23_72 V23 V72 6468.832430455454
L23_72 V23 V72 3.67302642213777e-12
C23_72 V23 V72 8.944361654038401e-20

R23_73 V23 V73 5233.572115258647
L23_73 V23 V73 3.813555128296361e-11
C23_73 V23 V73 5.158938133952434e-21

R23_74 V23 V74 -10546.854812156314
L23_74 V23 V74 -5.723059484448693e-12
C23_74 V23 V74 -3.1871019832707206e-20

R23_75 V23 V75 -5053.591913815299
L23_75 V23 V75 5.504991684626713e-12
C23_75 V23 V75 1.8500840204618134e-19

R23_76 V23 V76 -3064.364512838356
L23_76 V23 V76 -2.0553203341237347e-12
C23_76 V23 V76 -1.7881636483037442e-19

R23_77 V23 V77 -5582.418547298451
L23_77 V23 V77 -6.139450732884501e-12
C23_77 V23 V77 7.665903083614372e-20

R23_78 V23 V78 8908.67914981143
L23_78 V23 V78 -1.3231870169795577e-11
C23_78 V23 V78 -1.2196982137015312e-19

R23_79 V23 V79 -7125.33665240825
L23_79 V23 V79 -6.679592079917691e-12
C23_79 V23 V79 5.345579310460071e-20

R23_80 V23 V80 -16892.67872294295
L23_80 V23 V80 2.2326009677777456e-11
C23_80 V23 V80 3.5597559255127953e-20

R23_81 V23 V81 2280.776126360939
L23_81 V23 V81 3.3577912629631403e-12
C23_81 V23 V81 3.328181326905459e-20

R23_82 V23 V82 -10483.19347902811
L23_82 V23 V82 3.956806638875386e-12
C23_82 V23 V82 1.6931088201642435e-19

R23_83 V23 V83 -30733.772120402737
L23_83 V23 V83 -6.9908678599481515e-12
C23_83 V23 V83 -1.3532992056362693e-19

R23_84 V23 V84 -64284.54813195857
L23_84 V23 V84 5.028760387706439e-12
C23_84 V23 V84 1.0899754064944653e-19

R23_85 V23 V85 -48619.395704865245
L23_85 V23 V85 9.567499089921497e-12
C23_85 V23 V85 -3.2122548848078468e-21

R23_86 V23 V86 9569.638945663
L23_86 V23 V86 5.643507034831547e-12
C23_86 V23 V86 9.419621001185584e-20

R23_87 V23 V87 -6484.477424489938
L23_87 V23 V87 -3.226090711002988e-11
C23_87 V23 V87 -1.4465530211602062e-19

R23_88 V23 V88 57358.156155938326
L23_88 V23 V88 -6.544402817851432e-12
C23_88 V23 V88 -1.3685468674481229e-19

R23_89 V23 V89 16771.449401105896
L23_89 V23 V89 -1.6618548367024437e-11
C23_89 V23 V89 -1.1189423485281384e-19

R23_90 V23 V90 -14671.649518588945
L23_90 V23 V90 -1.7358255491716987e-12
C23_90 V23 V90 -3.009314914665745e-19

R23_91 V23 V91 1322.9319030059341
L23_91 V23 V91 2.3110362425633903e-12
C23_91 V23 V91 3.490956162359954e-19

R23_92 V23 V92 31312.554139621505
L23_92 V23 V92 4.438172696997422e-12
C23_92 V23 V92 9.814235759468568e-20

R23_93 V23 V93 3303.1163938309633
L23_93 V23 V93 -8.113455670593331e-12
C23_93 V23 V93 1.331240930444153e-20

R23_94 V23 V94 -11484.445155337453
L23_94 V23 V94 8.800553921558944e-12
C23_94 V23 V94 6.046626870564287e-20

R23_95 V23 V95 -2238.7789589652107
L23_95 V23 V95 1.6395747810882055e-10
C23_95 V23 V95 7.574446898790547e-20

R23_96 V23 V96 -3500.0959551083497
L23_96 V23 V96 -1.0183990864969808e-11
C23_96 V23 V96 3.639107670453746e-20

R23_97 V23 V97 44649.93954872682
L23_97 V23 V97 1.1819980717952686e-11
C23_97 V23 V97 2.3358732115764895e-19

R23_98 V23 V98 12634.783398117932
L23_98 V23 V98 2.4390545802288106e-12
C23_98 V23 V98 2.3439921305520535e-19

R23_99 V23 V99 -2303.827083446854
L23_99 V23 V99 -3.086210425738361e-12
C23_99 V23 V99 -3.857718117220554e-19

R23_100 V23 V100 -16601.169871877737
L23_100 V23 V100 -4.415579794789784e-12
C23_100 V23 V100 -1.6357612962738972e-19

R23_101 V23 V101 843280.0187731973
L23_101 V23 V101 9.597724671066653e-12
C23_101 V23 V101 -1.3316861260585373e-19

R23_102 V23 V102 -48719.3244905357
L23_102 V23 V102 -3.862671016422778e-12
C23_102 V23 V102 -8.574844293575861e-20

R23_103 V23 V103 2020.2295432549313
L23_103 V23 V103 -2.176504130462917e-12
C23_103 V23 V103 -2.3031378797453583e-20

R23_104 V23 V104 5974.444390110014
L23_104 V23 V104 6.12990005955147e-12
C23_104 V23 V104 1.3053301991559235e-19

R23_105 V23 V105 1598.1449031737106
L23_105 V23 V105 1.2193487728969686e-11
C23_105 V23 V105 -9.003713310958152e-20

R23_106 V23 V106 39502.40805471882
L23_106 V23 V106 -5.5312561748368126e-12
C23_106 V23 V106 -2.5780471995503457e-19

R23_107 V23 V107 17536.432771035565
L23_107 V23 V107 1.5283435597649547e-12
C23_107 V23 V107 3.2972711978713637e-19

R23_108 V23 V108 -19908.182565409894
L23_108 V23 V108 -1.5379897907258447e-11
C23_108 V23 V108 -6.407159207736814e-20

R23_109 V23 V109 -5775.64926102984
L23_109 V23 V109 -1.3754684104998654e-10
C23_109 V23 V109 1.936476133632831e-19

R23_110 V23 V110 -4220.008596759483
L23_110 V23 V110 5.4385668257056046e-12
C23_110 V23 V110 1.6678225115932735e-19

R23_111 V23 V111 -43784.43283274792
L23_111 V23 V111 1.3668939405489755e-12
C23_111 V23 V111 1.489189652093524e-19

R23_112 V23 V112 19055.588264949605
L23_112 V23 V112 1.0647528106821994e-11
C23_112 V23 V112 -2.96977697681107e-20

R23_113 V23 V113 7122.240931367149
L23_113 V23 V113 -3.564188314241305e-11
C23_113 V23 V113 3.442697590414458e-20

R23_114 V23 V114 -11590.299314682235
L23_114 V23 V114 2.1223632476062526e-11
C23_114 V23 V114 2.0870518572659096e-19

R23_115 V23 V115 -2076.9096171669316
L23_115 V23 V115 -1.0088789532978676e-12
C23_115 V23 V115 -3.9264346760118495e-19

R23_116 V23 V116 -4235.599585539772
L23_116 V23 V116 -5.6568604994725795e-12
C23_116 V23 V116 8.133920642973908e-20

R23_117 V23 V117 -12712.509910752497
L23_117 V23 V117 -3.629363327831753e-11
C23_117 V23 V117 -1.1666854505719648e-19

R23_118 V23 V118 3881.9155867817503
L23_118 V23 V118 -1.8892168180694374e-11
C23_118 V23 V118 -2.1387498425005634e-19

R23_119 V23 V119 1509.5610019322748
L23_119 V23 V119 -3.231709753280082e-12
C23_119 V23 V119 -1.2772455003197625e-20

R23_120 V23 V120 4150.524152638387
L23_120 V23 V120 -6.220726148154752e-12
C23_120 V23 V120 -1.34057829524236e-19

R23_121 V23 V121 4647.254566864862
L23_121 V23 V121 2.2064222282483522e-10
C23_121 V23 V121 4.143266296156561e-20

R23_122 V23 V122 -17382.28062681358
L23_122 V23 V122 8.920907391553503e-10
C23_122 V23 V122 -2.6939239671231393e-20

R23_123 V23 V123 -14124.524461825682
L23_123 V23 V123 9.298751927640848e-13
C23_123 V23 V123 4.490169256342569e-19

R23_124 V23 V124 12797.411555768014
L23_124 V23 V124 2.6070562383739557e-12
C23_124 V23 V124 9.510100307264087e-20

R23_125 V23 V125 1426.8781418321669
L23_125 V23 V125 2.87788062728898e-11
C23_125 V23 V125 1.2144473408448099e-20

R23_126 V23 V126 -12536.263627211549
L23_126 V23 V126 6.027466334999537e-12
C23_126 V23 V126 1.3501189648019898e-19

R23_127 V23 V127 -2727.056305332636
L23_127 V23 V127 7.014255745065915e-11
C23_127 V23 V127 -1.9659253375451836e-19

R23_128 V23 V128 -3247.9004123636264
L23_128 V23 V128 1.9897632092960952e-11
C23_128 V23 V128 5.723669261925244e-20

R23_129 V23 V129 -1558.3692310015008
L23_129 V23 V129 2.696009302098654e-12
C23_129 V23 V129 5.1441452296460063e-20

R23_130 V23 V130 -5523.751899924645
L23_130 V23 V130 -6.4337073289427226e-12
C23_130 V23 V130 -6.24937520107158e-20

R23_131 V23 V131 5457.664096237291
L23_131 V23 V131 -1.7634990726276997e-12
C23_131 V23 V131 -1.622619670562978e-19

R23_132 V23 V132 3252.7294956058836
L23_132 V23 V132 -2.2836325629447658e-12
C23_132 V23 V132 -1.940760591572824e-19

R23_133 V23 V133 -4997.115077819924
L23_133 V23 V133 -4.734426151962204e-12
C23_133 V23 V133 -2.1943658863767697e-20

R23_134 V23 V134 13374.923696351922
L23_134 V23 V134 -4.171162259117389e-12
C23_134 V23 V134 -4.9350902985729714e-20

R23_135 V23 V135 -4624.397179723117
L23_135 V23 V135 4.061757491101213e-12
C23_135 V23 V135 4.023973244414708e-19

R23_136 V23 V136 10234.166724151804
L23_136 V23 V136 -3.126448509781723e-11
C23_136 V23 V136 9.746642381882841e-20

R23_137 V23 V137 1518.254795187443
L23_137 V23 V137 -1.4021780875150117e-12
C23_137 V23 V137 -3.719193163731867e-20

R23_138 V23 V138 20529.79162226504
L23_138 V23 V138 3.377200890481667e-12
C23_138 V23 V138 1.0113601323153122e-19

R23_139 V23 V139 2566.721424654835
L23_139 V23 V139 -1.9113815639755953e-12
C23_139 V23 V139 -4.247119640353506e-19

R23_140 V23 V140 -14892.991012041868
L23_140 V23 V140 2.0027895916601493e-11
C23_140 V23 V140 -8.632174833996125e-20

R23_141 V23 V141 23115.68147032421
L23_141 V23 V141 1.7065067104265578e-12
C23_141 V23 V141 1.0984645871875566e-19

R23_142 V23 V142 -2421.521283652809
L23_142 V23 V142 2.7437957318814387e-12
C23_142 V23 V142 1.4546063018098995e-20

R23_143 V23 V143 2976.2880857262444
L23_143 V23 V143 1.1642922962112834e-12
C23_143 V23 V143 8.383481270739491e-20

R23_144 V23 V144 -5874.423265969815
L23_144 V23 V144 5.899158478408156e-12
C23_144 V23 V144 1.3119697605875309e-20

R23_145 V23 V145 -3969.406882623209
L23_145 V23 V145 9.204657809315395e-13
C23_145 V23 V145 6.540439157953434e-20

R23_146 V23 V146 6212.623205992908
L23_146 V23 V146 -9.93243572609982e-12
C23_146 V23 V146 -9.279160112339823e-20

R23_147 V23 V147 -533.8338759735411
L23_147 V23 V147 8.179543524023772e-11
C23_147 V23 V147 2.4534429578917343e-19

R23_148 V23 V148 4648.2986533130625
L23_148 V23 V148 2.859935770373902e-12
C23_148 V23 V148 7.392139493746252e-20

R23_149 V23 V149 -2280.3897476690545
L23_149 V23 V149 -1.0010210318621168e-12
C23_149 V23 V149 -2.1709726481910424e-19

R23_150 V23 V150 1843.0483822919364
L23_150 V23 V150 -3.5333184397181325e-12
C23_150 V23 V150 7.614691491973626e-20

R23_151 V23 V151 536.5535327983939
L23_151 V23 V151 -1.0728008816507847e-12
C23_151 V23 V151 -7.178309266791147e-20

R23_152 V23 V152 -11868.584038122832
L23_152 V23 V152 -6.410474151516401e-11
C23_152 V23 V152 4.394652336392125e-21

R23_153 V23 V153 1752.5733681059123
L23_153 V23 V153 -1.1061888359371106e-12
C23_153 V23 V153 2.3391482402779868e-20

R23_154 V23 V154 5631.075686083072
L23_154 V23 V154 -2.988580714325697e-12
C23_154 V23 V154 2.2191722146749298e-20

R23_155 V23 V155 -398.53695826716364
L23_155 V23 V155 -2.8963634823506177e-12
C23_155 V23 V155 -2.730950749708437e-19

R23_156 V23 V156 2050.9503552596093
L23_156 V23 V156 -3.468449951749689e-12
C23_156 V23 V156 -5.07406021908489e-20

R23_157 V23 V157 1238.7630914080169
L23_157 V23 V157 2.21100699546054e-12
C23_157 V23 V157 1.746686238070884e-19

R23_158 V23 V158 -3616.6530389623977
L23_158 V23 V158 3.5956438005962276e-12
C23_158 V23 V158 -4.796746801185358e-20

R23_159 V23 V159 950.76447258138
L23_159 V23 V159 7.104999993460091e-13
C23_159 V23 V159 2.174557531175832e-19

R23_160 V23 V160 -2443.624653474142
L23_160 V23 V160 -3.141993991845305e-12
C23_160 V23 V160 -9.351469551657993e-21

R23_161 V23 V161 -2598.0397228694765
L23_161 V23 V161 2.274122246982356e-12
C23_161 V23 V161 -7.328557883031998e-20

R23_162 V23 V162 -7247.4473888527245
L23_162 V23 V162 -8.091702097362955e-12
C23_162 V23 V162 -7.323447070246849e-20

R23_163 V23 V163 -1737.686184447021
L23_163 V23 V163 -2.231074159196962e-12
C23_163 V23 V163 -1.3592093994040108e-19

R23_164 V23 V164 2338.4648727725585
L23_164 V23 V164 3.0454745668789796e-12
C23_164 V23 V164 -4.9900067275204613e-20

R23_165 V23 V165 3445.2114877938693
L23_165 V23 V165 3.678877484568305e-12
C23_165 V23 V165 1.6558907029586625e-20

R23_166 V23 V166 3789.9323040540635
L23_166 V23 V166 4.942496362555427e-11
C23_166 V23 V166 7.806484725776765e-20

R23_167 V23 V167 778.2989759847364
L23_167 V23 V167 -1.1736442210887894e-12
C23_167 V23 V167 3.905330579134677e-20

R23_168 V23 V168 -966.4658625817272
L23_168 V23 V168 4.151023097238612e-12
C23_168 V23 V168 -9.298958844968344e-21

R23_169 V23 V169 2874.3712115037456
L23_169 V23 V169 -3.2046599203498573e-12
C23_169 V23 V169 9.793075906113858e-20

R23_170 V23 V170 5581.515385759742
L23_170 V23 V170 4.501227049207391e-12
C23_170 V23 V170 -4.7030483331641575e-20

R23_171 V23 V171 -1298.0308797539185
L23_171 V23 V171 1.069969816130354e-12
C23_171 V23 V171 6.707637191458386e-21

R23_172 V23 V172 4315.734728359527
L23_172 V23 V172 2.0865799112696562e-10
C23_172 V23 V172 2.757572458330776e-20

R23_173 V23 V173 11215.631301683734
L23_173 V23 V173 -7.63729195858805e-12
C23_173 V23 V173 -7.395281883107125e-20

R23_174 V23 V174 -1332.2648782986198
L23_174 V23 V174 -1.9420018190903186e-12
C23_174 V23 V174 4.07454961912037e-20

R23_175 V23 V175 -2418.1615682650636
L23_175 V23 V175 -3.3219334236236944e-12
C23_175 V23 V175 -1.6540933213177083e-19

R23_176 V23 V176 -113260.87588825755
L23_176 V23 V176 -1.905235358552361e-12
C23_176 V23 V176 -4.9767745823352896e-20

R23_177 V23 V177 3262.083287586569
L23_177 V23 V177 5.003929993164991e-12
C23_177 V23 V177 1.3331639306949948e-20

R23_178 V23 V178 1907.4804709079583
L23_178 V23 V178 5.085942452484594e-12
C23_178 V23 V178 1.1095851079267766e-20

R23_179 V23 V179 -2112.6413347006583
L23_179 V23 V179 -2.320409412846458e-12
C23_179 V23 V179 1.5492969111932606e-19

R23_180 V23 V180 5093.334126391867
L23_180 V23 V180 2.919788015333053e-12
C23_180 V23 V180 6.744893012606474e-20

R23_181 V23 V181 -1701.5828202817534
L23_181 V23 V181 1.678235584276392e-11
C23_181 V23 V181 3.7901104811348194e-20

R23_182 V23 V182 -2862.905492560036
L23_182 V23 V182 -3.322755482869282e-11
C23_182 V23 V182 -3.4542803184412875e-20

R23_183 V23 V183 721.0074798213271
L23_183 V23 V183 1.8168186872448978e-12
C23_183 V23 V183 -1.3299389002016873e-21

R23_184 V23 V184 2748.3585019602892
L23_184 V23 V184 2.899792510305964e-12
C23_184 V23 V184 8.8464388520152e-21

R23_185 V23 V185 1860.0606986440425
L23_185 V23 V185 1.40634221751547e-11
C23_185 V23 V185 -3.1820616063107564e-20

R23_186 V23 V186 -5814.666191397931
L23_186 V23 V186 6.462799059033094e-12
C23_186 V23 V186 5.23876333557661e-20

R23_187 V23 V187 -1469.31273483015
L23_187 V23 V187 -6.639202734447168e-12
C23_187 V23 V187 -1.8539652093150048e-19

R23_188 V23 V188 -1185.5822366300642
L23_188 V23 V188 -3.24503407575093e-12
C23_188 V23 V188 -8.919367097474056e-20

R23_189 V23 V189 -8101.475942835165
L23_189 V23 V189 -4.531470384670638e-12
C23_189 V23 V189 1.7962822155818925e-20

R23_190 V23 V190 3663.6338839672717
L23_190 V23 V190 -2.1487948040498226e-11
C23_190 V23 V190 1.830082160940671e-20

R23_191 V23 V191 -1836.9416771679112
L23_191 V23 V191 -4.6230559445878614e-12
C23_191 V23 V191 1.5627793982135256e-19

R23_192 V23 V192 16246.904621222224
L23_192 V23 V192 -5.946659185379368e-12
C23_192 V23 V192 5.96185824551613e-20

R23_193 V23 V193 -3725.825568533599
L23_193 V23 V193 -3.206481073871276e-11
C23_193 V23 V193 2.1360740644327865e-20

R23_194 V23 V194 -7732.108044433437
L23_194 V23 V194 -3.840395748364682e-12
C23_194 V23 V194 8.102660395926887e-20

R23_195 V23 V195 1117.3640247623796
L23_195 V23 V195 2.9686423825703197e-12
C23_195 V23 V195 -1.4184326297070529e-19

R23_196 V23 V196 1091.8469095022958
L23_196 V23 V196 9.012545120911147e-12
C23_196 V23 V196 4.9472547800387647e-20

R23_197 V23 V197 3416.0320041415434
L23_197 V23 V197 3.619081320296775e-12
C23_197 V23 V197 -2.1159704782236342e-20

R23_198 V23 V198 9866.27469988499
L23_198 V23 V198 4.471951592095348e-11
C23_198 V23 V198 7.3241646687016e-22

R23_199 V23 V199 -341158.52466844866
L23_199 V23 V199 3.905770333167361e-11
C23_199 V23 V199 -4.509429485362441e-20

R23_200 V23 V200 -2329.365662025315
L23_200 V23 V200 4.1947069470213835e-12
C23_200 V23 V200 -7.438326176154487e-20

R24_24 V24 0 -167.63421766945385
L24_24 V24 0 -2.2022397284321856e-13
C24_24 V24 0 -1.2852437218304825e-18

R24_25 V24 V25 1242.92877954492
L24_25 V24 V25 3.1872040407710267e-12
C24_25 V24 V25 -1.3915374667508383e-19

R24_26 V24 V26 3586.856449783964
L24_26 V24 V26 -1.3679912583251991e-11
C24_26 V24 V26 -1.4616609738557548e-19

R24_27 V24 V27 4172.682640130067
L24_27 V24 V27 3.4062870573972217e-12
C24_27 V24 V27 2.4657332744385147e-20

R24_28 V24 V28 1467.6877860596608
L24_28 V24 V28 8.304257252186763e-13
C24_28 V24 V28 3.4277949374598466e-19

R24_29 V24 V29 1354.392065706396
L24_29 V24 V29 1.880496160655407e-12
C24_29 V24 V29 8.675585973798185e-20

R24_30 V24 V30 4538.187437551223
L24_30 V24 V30 2.9289304196701505e-12
C24_30 V24 V30 1.3987046891836193e-19

R24_31 V24 V31 2691.366327915766
L24_31 V24 V31 3.0112240205638474e-12
C24_31 V24 V31 1.4417664691114023e-19

R24_32 V24 V32 1283.8712082318343
L24_32 V24 V32 9.811282750914233e-13
C24_32 V24 V32 4.723446452858054e-19

R24_33 V24 V33 4151.357147401567
L24_33 V24 V33 8.296464890365367e-12
C24_33 V24 V33 5.722693929918086e-20

R24_34 V24 V34 -6825.484908390382
L24_34 V24 V34 6.848603601209749e-12
C24_34 V24 V34 1.429490274177554e-19

R24_35 V24 V35 -5456.165669977316
L24_35 V24 V35 -4.454676877738492e-12
C24_35 V24 V35 -8.654762239929302e-20

R24_36 V24 V36 -1621.5074531244363
L24_36 V24 V36 -7.464272936402864e-13
C24_36 V24 V36 -9.00644567842548e-19

R24_37 V24 V37 -3193.2944376528712
L24_37 V24 V37 -1.7523882533903185e-12
C24_37 V24 V37 -7.986482526806359e-20

R24_38 V24 V38 -6879.3682987384345
L24_38 V24 V38 -1.6122636713554498e-12
C24_38 V24 V38 -2.8849289106043723e-19

R24_39 V24 V39 -3489.644094130444
L24_39 V24 V39 -4.552047669571387e-12
C24_39 V24 V39 -2.1234460860735692e-20

R24_40 V24 V40 -1765.791268692471
L24_40 V24 V40 -2.7052562965449853e-12
C24_40 V24 V40 1.1807834086044593e-19

R24_41 V24 V41 -99277.07416686123
L24_41 V24 V41 -1.1452955802608096e-11
C24_41 V24 V41 9.196555789632629e-21

R24_42 V24 V42 -51449.477732333915
L24_42 V24 V42 -1.3470016986969532e-10
C24_42 V24 V42 8.10893252987209e-20

R24_43 V24 V43 -17285.644452794957
L24_43 V24 V43 -6.8613217524119325e-12
C24_43 V24 V43 1.1115241189055762e-20

R24_44 V24 V44 -2878.699659526365
L24_44 V24 V44 1.142961091067198e-11
C24_44 V24 V44 1.529313764469657e-19

R24_45 V24 V45 2295.866721982406
L24_45 V24 V45 2.9420413957884607e-12
C24_45 V24 V45 -4.0864381301161015e-20

R24_46 V24 V46 4823.528980503108
L24_46 V24 V46 1.8616248416368178e-12
C24_46 V24 V46 2.727334235963471e-19

R24_47 V24 V47 4606.245404601631
L24_47 V24 V47 3.12922365463976e-12
C24_47 V24 V47 8.968802033681738e-20

R24_48 V24 V48 1829.2359185148039
L24_48 V24 V48 1.0724269297988424e-12
C24_48 V24 V48 2.196448744924318e-19

R24_49 V24 V49 3051.36688741351
L24_49 V24 V49 4.055108668456308e-12
C24_49 V24 V49 9.503207387105297e-20

R24_50 V24 V50 58282.19333389446
L24_50 V24 V50 -4.598799725346651e-12
C24_50 V24 V50 -2.191117586615748e-19

R24_51 V24 V51 7687.4929307210405
L24_51 V24 V51 1.5315302839056452e-11
C24_51 V24 V51 -6.855744023061782e-20

R24_52 V24 V52 14931.92459320387
L24_52 V24 V52 -5.936344765546962e-12
C24_52 V24 V52 6.1731534329687616e-21

R24_53 V24 V53 3446.352388578908
L24_53 V24 V53 2.4080823292880624e-12
C24_53 V24 V53 1.6432357152112468e-19

R24_54 V24 V54 -36598.12087249614
L24_54 V24 V54 9.72699347240464e-11
C24_54 V24 V54 4.6090929627694073e-20

R24_55 V24 V55 17355.67181823237
L24_55 V24 V55 1.4001894585984675e-11
C24_55 V24 V55 4.97259208557866e-20

R24_56 V24 V56 -7101.890209882037
L24_56 V24 V56 -9.046946707300624e-13
C24_56 V24 V56 -6.646197293269272e-19

R24_57 V24 V57 -29870.004797331276
L24_57 V24 V57 -1.2520753171697934e-12
C24_57 V24 V57 -2.1556677617458463e-19

R24_58 V24 V58 17836.959762266153
L24_58 V24 V58 2.0109387210147277e-11
C24_58 V24 V58 8.353515283134583e-20

R24_59 V24 V59 -4169.364400059487
L24_59 V24 V59 -2.1059532482517936e-11
C24_59 V24 V59 9.900347896118979e-20

R24_60 V24 V60 -1385.3281830195142
L24_60 V24 V60 8.214739237550583e-12
C24_60 V24 V60 1.9357235039180815e-19

R24_61 V24 V61 -17263.96982187435
L24_61 V24 V61 4.703639461743609e-12
C24_61 V24 V61 1.9085222395947318e-20

R24_62 V24 V62 -7226.110805377345
L24_62 V24 V62 -5.74214895813012e-12
C24_62 V24 V62 -7.395864054132467e-20

R24_63 V24 V63 48836.33465201648
L24_63 V24 V63 -3.0083942633077115e-12
C24_63 V24 V63 -1.5287005734802259e-19

R24_64 V24 V64 4827.014013664084
L24_64 V24 V64 1.2953191022662144e-12
C24_64 V24 V64 4.370454855683657e-19

R24_65 V24 V65 3852.266963679847
L24_65 V24 V65 1.904754109269867e-12
C24_65 V24 V65 2.3681778084374694e-19

R24_66 V24 V66 12267.421235309774
L24_66 V24 V66 4.879016028299769e-12
C24_66 V24 V66 9.42917269056298e-20

R24_67 V24 V67 29914.30514050007
L24_67 V24 V67 5.570262963078849e-12
C24_67 V24 V67 4.939908159621919e-20

R24_68 V24 V68 3932.2021292302743
L24_68 V24 V68 -4.98601546115623e-12
C24_68 V24 V68 -2.0335232938488875e-19

R24_69 V24 V69 4614.857757318631
L24_69 V24 V69 -5.669485251287407e-12
C24_69 V24 V69 -2.042971573374956e-19

R24_70 V24 V70 39722.43144125313
L24_70 V24 V70 8.862452903971405e-12
C24_70 V24 V70 1.6821414870078625e-20

R24_71 V24 V71 9651.962837248762
L24_71 V24 V71 2.7201496234688835e-12
C24_71 V24 V71 1.203617514731702e-19

R24_72 V24 V72 6258.496710139719
L24_72 V24 V72 1.737331885972093e-11
C24_72 V24 V72 -1.5434489758041685e-19

R24_73 V24 V73 5108.014971328352
L24_73 V24 V73 -3.329145889058583e-11
C24_73 V24 V73 -3.09538562157362e-20

R24_74 V24 V74 -7857.797475437605
L24_74 V24 V74 -3.6224364566275763e-12
C24_74 V24 V74 -8.925133894362665e-20

R24_75 V24 V75 -39476.049611579125
L24_75 V24 V75 -3.965295058150158e-12
C24_75 V24 V75 -4.7454010650970885e-20

R24_76 V24 V76 -2312.5800388278767
L24_76 V24 V76 -5.050319328616788e-12
C24_76 V24 V76 2.747080755078001e-20

R24_77 V24 V77 -5117.108290307997
L24_77 V24 V77 -5.8463024285076126e-12
C24_77 V24 V77 1.0507651343425741e-19

R24_78 V24 V78 5338.251369154625
L24_78 V24 V78 -2.7511117975431566e-11
C24_78 V24 V78 -9.660381009015094e-20

R24_79 V24 V79 -7137.159956024223
L24_79 V24 V79 -8.531805393091326e-12
C24_79 V24 V79 -5.906401008405144e-20

R24_80 V24 V80 -50629.30362085417
L24_80 V24 V80 -1.246821643262016e-11
C24_80 V24 V80 1.4618118882496178e-19

R24_81 V24 V81 1519.6642831036177
L24_81 V24 V81 1.9884478706840636e-12
C24_81 V24 V81 1.2535264473888777e-19

R24_82 V24 V82 -7268.406316769432
L24_82 V24 V82 2.733693546664193e-12
C24_82 V24 V82 2.2880314805225366e-19

R24_83 V24 V83 -34762.119834920835
L24_83 V24 V83 1.0406260191989752e-11
C24_83 V24 V83 9.50921001265188e-20

R24_84 V24 V84 -37613.13972474909
L24_84 V24 V84 4.077783911413733e-12
C24_84 V24 V84 -3.587230220478949e-20

R24_85 V24 V85 -44908.77642813692
L24_85 V24 V85 9.24750115252049e-12
C24_85 V24 V85 -3.0511971666058325e-20

R24_86 V24 V86 17202.834537284587
L24_86 V24 V86 5.088698822316712e-12
C24_86 V24 V86 7.712075546104397e-20

R24_87 V24 V87 -881999.3014904852
L24_87 V24 V87 -1.0238884378442793e-11
C24_87 V24 V87 -7.333728259745735e-20

R24_88 V24 V88 -4533.7325325537195
L24_88 V24 V88 -5.384965890749655e-12
C24_88 V24 V88 -2.0792976588497341e-19

R24_89 V24 V89 18425.325307127743
L24_89 V24 V89 -9.60026685657208e-12
C24_89 V24 V89 -1.5018677478706182e-19

R24_90 V24 V90 -24539.098753726626
L24_90 V24 V90 -1.3425551550093865e-12
C24_90 V24 V90 -3.369113721783271e-19

R24_91 V24 V91 3664.4299491478528
L24_91 V24 V91 2.21450422489236e-12
C24_91 V24 V91 1.3665017304295612e-19

R24_92 V24 V92 1593.9813329716337
L24_92 V24 V92 4.046164208018563e-12
C24_92 V24 V92 2.1443852344295033e-19

R24_93 V24 V93 2658.8586002995767
L24_93 V24 V93 -7.344225960007941e-12
C24_93 V24 V93 4.856089385868701e-20

R24_94 V24 V94 -9756.401885043524
L24_94 V24 V94 4.735848356654817e-12
C24_94 V24 V94 1.1109877609385288e-19

R24_95 V24 V95 -4490.382249189946
L24_95 V24 V95 -1.4360254544991768e-11
C24_95 V24 V95 2.9292354648053946e-20

R24_96 V24 V96 -2277.5180321817957
L24_96 V24 V96 1.542735879981557e-11
C24_96 V24 V96 1.2567486766944188e-19

R24_97 V24 V97 11112.257391154952
L24_97 V24 V97 6.470265010971674e-12
C24_97 V24 V97 2.7102825314896005e-19

R24_98 V24 V98 20232.268084952964
L24_98 V24 V98 1.9208810566901087e-12
C24_98 V24 V98 2.617004731170328e-19

R24_99 V24 V99 -3543.3498498992262
L24_99 V24 V99 -1.999728127016865e-12
C24_99 V24 V99 -1.6226856485935675e-19

R24_100 V24 V100 -1749.965761713475
L24_100 V24 V100 -4.747653388543721e-12
C24_100 V24 V100 -3.2310494420843754e-19

R24_101 V24 V101 -36594.785729579686
L24_101 V24 V101 5.46321834861852e-12
C24_101 V24 V101 -1.23678735656913e-19

R24_102 V24 V102 139066.27902402403
L24_102 V24 V102 -2.377221130573792e-12
C24_102 V24 V102 -1.3973672405856e-19

R24_103 V24 V103 3960.716976368678
L24_103 V24 V103 6.898834628686706e-12
C24_103 V24 V103 7.145115433966712e-20

R24_104 V24 V104 2083.8920568227113
L24_104 V24 V104 -2.7071519260844113e-12
C24_104 V24 V104 -2.9740752285992685e-20

R24_105 V24 V105 1317.2758281116267
L24_105 V24 V105 1.8692961637941734e-11
C24_105 V24 V105 -1.0365531024509402e-19

R24_106 V24 V106 -10311.865028366801
L24_106 V24 V106 -5.9089084157469295e-12
C24_106 V24 V106 -2.2357356908306974e-19

R24_107 V24 V107 132719.59308303404
L24_107 V24 V107 3.274414341085744e-12
C24_107 V24 V107 9.92485089169794e-20

R24_108 V24 V108 13558.089699308563
L24_108 V24 V108 3.308544245512123e-12
C24_108 V24 V108 1.9110374076938244e-19

R24_109 V24 V109 -5949.375598471083
L24_109 V24 V109 5.429583991441808e-11
C24_109 V24 V109 2.2740303442885653e-19

R24_110 V24 V110 -6046.39687023987
L24_110 V24 V110 5.464441998923486e-12
C24_110 V24 V110 1.4188606389214552e-19

R24_111 V24 V111 96738.11877608288
L24_111 V24 V111 4.8687403891549545e-12
C24_111 V24 V111 -4.683690719576868e-20

R24_112 V24 V112 -7473.298515279756
L24_112 V24 V112 1.100606342653198e-12
C24_112 V24 V112 3.0734556905709196e-19

R24_113 V24 V113 5229.373265836714
L24_113 V24 V113 -3.9630574637086797e-11
C24_113 V24 V113 4.660772098601267e-20

R24_114 V24 V114 -21169.264055815023
L24_114 V24 V114 3.582936324903049e-11
C24_114 V24 V114 1.844454404630861e-19

R24_115 V24 V115 -2584.1737814137286
L24_115 V24 V115 -1.8388913638630725e-12
C24_115 V24 V115 -4.469973728748796e-20

R24_116 V24 V116 -2263.4704523848336
L24_116 V24 V116 -1.0780785280167943e-12
C24_116 V24 V116 -3.534584721703844e-19

R24_117 V24 V117 -12390.05229886769
L24_117 V24 V117 -1.6115904583884356e-11
C24_117 V24 V117 -1.6373256469816393e-19

R24_118 V24 V118 7190.959409700758
L24_118 V24 V118 -1.435297591176161e-11
C24_118 V24 V118 -2.1279924235912923e-19

R24_119 V24 V119 5142.985062458724
L24_119 V24 V119 -8.617860436858167e-12
C24_119 V24 V119 -1.0114137494922196e-19

R24_120 V24 V120 1286.8263874256718
L24_120 V24 V120 -1.6648105554632006e-12
C24_120 V24 V120 -2.1143355673529994e-19

R24_121 V24 V121 3935.6460828469812
L24_121 V24 V121 -4.1336319952805463e-10
C24_121 V24 V121 7.047752139849983e-20

R24_122 V24 V122 -40930.148110910675
L24_122 V24 V122 -3.5568920654942975e-11
C24_122 V24 V122 -2.5361829338120308e-20

R24_123 V24 V123 6154.273487028217
L24_123 V24 V123 2.255269374518686e-12
C24_123 V24 V123 5.1512151730289874e-20

R24_124 V24 V124 -2960.5202985898823
L24_124 V24 V124 6.828141861353903e-13
C24_124 V24 V124 6.831208265702561e-19

R24_125 V24 V125 1175.917416528483
L24_125 V24 V125 1.3926677107329289e-11
C24_125 V24 V125 5.241894456798212e-20

R24_126 V24 V126 58120.42196311855
L24_126 V24 V126 5.020757646209488e-12
C24_126 V24 V126 1.1079322802754886e-19

R24_127 V24 V127 -3637.057173352485
L24_127 V24 V127 -2.979647117269899e-11
C24_127 V24 V127 1.190515307077171e-19

R24_128 V24 V128 -3253.519401830141
L24_128 V24 V128 1.2402211724216959e-11
C24_128 V24 V128 -1.4787690774060173e-19

R24_129 V24 V129 -1433.9372686446861
L24_129 V24 V129 1.994893452070544e-12
C24_129 V24 V129 4.565528187854967e-20

R24_130 V24 V130 -4484.663367814149
L24_130 V24 V130 -4.6969335827803295e-12
C24_130 V24 V130 -9.86923683819498e-20

R24_131 V24 V131 3370.590288823165
L24_131 V24 V131 -6.157828416780339e-12
C24_131 V24 V131 -1.3253639773286529e-19

R24_132 V24 V132 3832.258606871783
L24_132 V24 V132 -9.853701435032628e-13
C24_132 V24 V132 -3.3170455121825485e-19

R24_133 V24 V133 -4298.303850327253
L24_133 V24 V133 -2.5326709772926887e-12
C24_133 V24 V133 -1.0540845929443344e-19

R24_134 V24 V134 15806.67337339523
L24_134 V24 V134 -2.6114276056260998e-12
C24_134 V24 V134 -8.800668567561511e-20

R24_135 V24 V135 -5876.40807829094
L24_135 V24 V135 -7.92293936226795e-12
C24_135 V24 V135 -5.842934027618942e-20

R24_136 V24 V136 -4406.739345081534
L24_136 V24 V136 2.9819021734454567e-12
C24_136 V24 V136 4.732526379562436e-19

R24_137 V24 V137 1481.9951730396313
L24_137 V24 V137 -1.2134853214627833e-12
C24_137 V24 V137 -1.95416773347872e-20

R24_138 V24 V138 7095.774961020255
L24_138 V24 V138 2.319461128192577e-12
C24_138 V24 V138 1.1193673887121727e-19

R24_139 V24 V139 -8725.43210305499
L24_139 V24 V139 -2.2076767851953726e-11
C24_139 V24 V139 4.220537315190624e-20

R24_140 V24 V140 1236.7998303919424
L24_140 V24 V140 -2.0966454237408677e-12
C24_140 V24 V140 -4.362554997535244e-19

R24_141 V24 V141 -11129.39836852838
L24_141 V24 V141 1.3344110903217663e-12
C24_141 V24 V141 1.761754291321107e-19

R24_142 V24 V142 -2011.8941217610413
L24_142 V24 V142 2.4095837633031803e-12
C24_142 V24 V142 1.7327833749557594e-20

R24_143 V24 V143 5894.134175641588
L24_143 V24 V143 3.2747004364662315e-12
C24_143 V24 V143 3.733892989072284e-20

R24_144 V24 V144 -1066.7168144317002
L24_144 V24 V144 1.2657241636379167e-12
C24_144 V24 V144 4.032292907511799e-20

R24_145 V24 V145 32484.04110267901
L24_145 V24 V145 7.646051662838785e-13
C24_145 V24 V145 5.82542828402898e-20

R24_146 V24 V146 -25081.421944996775
L24_146 V24 V146 -1.1933210454384774e-11
C24_146 V24 V146 -9.31624339380732e-20

R24_147 V24 V147 -1352.5657783212998
L24_147 V24 V147 2.9520380745425717e-12
C24_147 V24 V147 8.019709624216039e-20

R24_148 V24 V148 1198.8661170406924
L24_148 V24 V148 3.680427666572436e-12
C24_148 V24 V148 2.944014318654306e-19

R24_149 V24 V149 -1167.5775463818466
L24_149 V24 V149 -8.77890431714832e-13
C24_149 V24 V149 -2.2851960262150744e-19

R24_150 V24 V150 1893.914856163162
L24_150 V24 V150 -3.672962474927498e-12
C24_150 V24 V150 1.6179669279002675e-19

R24_151 V24 V151 1116.3118312611734
L24_151 V24 V151 -1.283019630822973e-11
C24_151 V24 V151 -2.893565530495698e-20

R24_152 V24 V152 -1096.3604091005323
L24_152 V24 V152 -8.987297283079404e-13
C24_152 V24 V152 -8.133410709646662e-20

R24_153 V24 V153 1375.5403422382944
L24_153 V24 V153 -7.957822155099154e-13
C24_153 V24 V153 -5.298945732738804e-20

R24_154 V24 V154 17451.35282463703
L24_154 V24 V154 -1.8220644245823737e-12
C24_154 V24 V154 -3.477300174904618e-20

R24_155 V24 V155 -674.4039877023476
L24_155 V24 V155 -1.5557641463188377e-12
C24_155 V24 V155 -5.813189420736813e-20

R24_156 V24 V156 460.0032233908014
L24_156 V24 V156 -1.5785406458405813e-11
C24_156 V24 V156 -2.0932145069422191e-19

R24_157 V24 V157 797.9911320876415
L24_157 V24 V157 1.4348334532680305e-12
C24_157 V24 V157 3.176749253757758e-19

R24_158 V24 V158 -8527.450678624391
L24_158 V24 V158 2.2036771188186797e-12
C24_158 V24 V158 -2.151790832601834e-20

R24_159 V24 V159 1035.2143000294864
L24_159 V24 V159 -1.0082383027036138e-11
C24_159 V24 V159 7.057769469686061e-21

R24_160 V24 V160 -852.2135245643717
L24_160 V24 V160 7.987108753879131e-13
C24_160 V24 V160 9.116242186859067e-20

R24_161 V24 V161 -2398.3260114355785
L24_161 V24 V161 1.8422259742517824e-12
C24_161 V24 V161 -4.6453290462781205e-20

R24_162 V24 V162 -5488.082599097591
L24_162 V24 V162 -1.0834800983852268e-11
C24_162 V24 V162 -5.942559555380402e-20

R24_163 V24 V163 -11746.28492711343
L24_163 V24 V163 6.816495200127973e-12
C24_163 V24 V163 3.279761828769293e-20

R24_164 V24 V164 4474.359441522508
L24_164 V24 V164 -6.510839028822826e-12
C24_164 V24 V164 -9.741687585951785e-20

R24_165 V24 V165 1845.2231084475336
L24_165 V24 V165 2.8475391717074816e-12
C24_165 V24 V165 -1.7191176324693978e-20

R24_166 V24 V166 2905.02872981667
L24_166 V24 V166 -3.294210851104375e-11
C24_166 V24 V166 1.297932052860842e-19

R24_167 V24 V167 3981.031364070831
L24_167 V24 V167 2.577120760705714e-12
C24_167 V24 V167 2.584914001356768e-21

R24_168 V24 V168 -2173.4894239233245
L24_168 V24 V168 -9.742720310056768e-13
C24_168 V24 V168 4.078875632786886e-20

R24_169 V24 V169 3782.4476071649174
L24_169 V24 V169 -2.5062777881092472e-12
C24_169 V24 V169 1.1016688844420631e-19

R24_170 V24 V170 4392.018336117017
L24_170 V24 V170 4.335368887816551e-12
C24_170 V24 V170 -5.579404036247265e-20

R24_171 V24 V171 -3427.8923072620732
L24_171 V24 V171 -8.658103561769302e-12
C24_171 V24 V171 -3.1279534652032896e-20

R24_172 V24 V172 2370.604455714337
L24_172 V24 V172 1.1982553057956796e-12
C24_172 V24 V172 -2.291983981111306e-20

R24_173 V24 V173 3602.353794206803
L24_173 V24 V173 -6.137321972997272e-12
C24_173 V24 V173 -6.855216087423255e-20

R24_174 V24 V174 -1074.9506922814994
L24_174 V24 V174 -1.6369911422301252e-12
C24_174 V24 V174 1.9619712272164133e-20

R24_175 V24 V175 20122.267560985347
L24_175 V24 V175 -1.6333476186492226e-12
C24_175 V24 V175 -4.692824406277105e-20

R24_176 V24 V176 -2144.1822701692827
L24_176 V24 V176 -3.3671165205387035e-12
C24_176 V24 V176 -2.2639980818868877e-19

R24_177 V24 V177 3747.7922632133495
L24_177 V24 V177 3.1708707242091897e-12
C24_177 V24 V177 1.676398029121712e-20

R24_178 V24 V178 1777.7814616290932
L24_178 V24 V178 3.251608796393157e-12
C24_178 V24 V178 2.727837030044755e-20

R24_179 V24 V179 -6724.73155013471
L24_179 V24 V179 1.7037311060006936e-12
C24_179 V24 V179 1.0658083009079042e-19

R24_180 V24 V180 71443.39764998673
L24_180 V24 V180 -3.202469182916133e-12
C24_180 V24 V180 2.399709984917528e-19

R24_181 V24 V181 -1415.36586248465
L24_181 V24 V181 8.356067175302273e-12
C24_181 V24 V181 6.8499751801874e-20

R24_182 V24 V182 -3326.5810831193144
L24_182 V24 V182 -1.8692226303164888e-11
C24_182 V24 V182 -3.201230332346481e-20

R24_183 V24 V183 1824.2631915111363
L24_183 V24 V183 3.57321163568315e-12
C24_183 V24 V183 4.992917618763769e-20

R24_184 V24 V184 949.1020949941138
L24_184 V24 V184 1.2464931709593967e-12
C24_184 V24 V184 -6.074450421175414e-20

R24_185 V24 V185 1201.5007429918464
L24_185 V24 V185 1.9679929657196397e-11
C24_185 V24 V185 -4.6864100980975086e-20

R24_186 V24 V186 -20525.088150962943
L24_186 V24 V186 4.0327916791558156e-12
C24_186 V24 V186 9.325531578722606e-21

R24_187 V24 V187 -9801.41651695462
L24_187 V24 V187 -3.4005027988242955e-12
C24_187 V24 V187 -1.2857715783566624e-19

R24_188 V24 V188 -617.6928315484782
L24_188 V24 V188 -2.0070213086831197e-12
C24_188 V24 V188 -1.2932489702213627e-19

R24_189 V24 V189 -2866.5084817965035
L24_189 V24 V189 -3.417544939963095e-12
C24_189 V24 V189 -1.38534906672582e-20

R24_190 V24 V190 3762.7699061292556
L24_190 V24 V190 -1.1779561652813176e-10
C24_190 V24 V190 7.029167877245316e-20

R24_191 V24 V191 -2857.702299970988
L24_191 V24 V191 -2.8684226022293914e-12
C24_191 V24 V191 -3.44474009266665e-20

R24_192 V24 V192 27801.419817963288
L24_192 V24 V192 -7.59919458664365e-12
C24_192 V24 V192 1.4953152125180964e-19

R24_193 V24 V193 -2185.578402413524
L24_193 V24 V193 -6.988251755973728e-11
C24_193 V24 V193 4.208669309064197e-20

R24_194 V24 V194 -10535.401195588574
L24_194 V24 V194 -3.4488211548937504e-12
C24_194 V24 V194 1.1763000983642374e-19

R24_195 V24 V195 1931.8063957878612
L24_195 V24 V195 2.1084246297198533e-12
C24_195 V24 V195 2.1191190140549585e-19

R24_196 V24 V196 758.7254404575692
L24_196 V24 V196 6.719288904843931e-12
C24_196 V24 V196 -2.414878452419957e-19

R24_197 V24 V197 2770.5627507880945
L24_197 V24 V197 2.8964747169980223e-12
C24_197 V24 V197 -2.3841300949854175e-20

R24_198 V24 V198 8097.702468617337
L24_198 V24 V198 1.6887283263685167e-11
C24_198 V24 V198 4.9912561555860405e-20

R24_199 V24 V199 1966.8828295546996
L24_199 V24 V199 5.204126891532492e-12
C24_199 V24 V199 3.4337027336513196e-20

R24_200 V24 V200 -1062.342567166599
L24_200 V24 V200 4.520829431985535e-12
C24_200 V24 V200 -1.22165986585054e-20

R25_25 V25 0 73.37129882897668
L25_25 V25 0 1.4712201158317021e-13
C25_25 V25 0 9.780899529079811e-19

R25_26 V25 V26 -1666.3298570922213
L25_26 V25 V26 -1.2341103444377822e-12
C25_26 V25 V26 -2.5888228874412926e-19

R25_27 V25 V27 -3262.331035461593
L25_27 V25 V27 -1.2869177969426242e-12
C25_27 V25 V27 -2.4583050612351916e-19

R25_28 V25 V28 -1930.4276123894585
L25_28 V25 V28 -8.541200279686715e-13
C25_28 V25 V28 -3.9417088122598807e-19

R25_29 V25 V29 -311.60977030799285
L25_29 V25 V29 -1.1223107396658728e-12
C25_29 V25 V29 2.19019043064864e-19

R25_30 V25 V30 -2902.9787251241346
L25_30 V25 V30 -7.745880296101128e-12
C25_30 V25 V30 1.2568979295316408e-19

R25_31 V25 V31 -2896.5526543478136
L25_31 V25 V31 -3.191500008150205e-11
C25_31 V25 V31 1.3948953735434807e-19

R25_32 V25 V32 -1913.5323806014096
L25_32 V25 V32 -3.78768791245257e-11
C25_32 V25 V32 2.0642778621636536e-19

R25_33 V25 V33 -712.4052565211299
L25_33 V25 V33 9.68574528735533e-12
C25_33 V25 V33 2.613772899868087e-19

R25_34 V25 V34 10006.613326736993
L25_34 V25 V34 1.474583980985701e-11
C25_34 V25 V34 1.2387455713486992e-19

R25_35 V25 V35 2947.0615081034166
L25_35 V25 V35 7.881367562010846e-12
C25_35 V25 V35 5.3389742794822415e-20

R25_36 V25 V36 1821.614660339154
L25_36 V25 V36 3.3980298391360596e-12
C25_36 V25 V36 9.349121796714641e-20

R25_37 V25 V37 721.0809337505814
L25_37 V25 V37 8.786162657670496e-13
C25_37 V25 V37 1.5695913757002185e-20

R25_38 V25 V38 3685.752311099669
L25_38 V25 V38 3.1278220959008446e-12
C25_38 V25 V38 -2.7914647090911045e-20

R25_39 V25 V39 2798.2834514258416
L25_39 V25 V39 3.651886001818104e-12
C25_39 V25 V39 -3.207835448462776e-20

R25_40 V25 V40 1815.0512243611474
L25_40 V25 V40 2.5117303589197947e-12
C25_40 V25 V40 -5.379078290831388e-20

R25_41 V25 V41 3591.778145054259
L25_41 V25 V41 3.1136313229960337e-12
C25_41 V25 V41 -1.2696332150152404e-20

R25_42 V25 V42 3642.1081419815428
L25_42 V25 V42 1.481754206617615e-11
C25_42 V25 V42 8.175452687263841e-22

R25_43 V25 V43 2539.1151628295447
L25_43 V25 V43 4.146098860200034e-12
C25_43 V25 V43 5.1814532919884666e-20

R25_44 V25 V44 2055.444188474917
L25_44 V25 V44 3.68940673550495e-12
C25_44 V25 V44 6.852608502896135e-20

R25_45 V25 V45 -595.0848703842378
L25_45 V25 V45 -6.794046222970294e-13
C25_45 V25 V45 -2.8132194393341223e-19

R25_46 V25 V46 -15972.76948851052
L25_46 V25 V46 1.297921849857095e-11
C25_46 V25 V46 2.2866341314892795e-20

R25_47 V25 V47 -13996.898274725445
L25_47 V25 V47 -7.371645201809796e-12
C25_47 V25 V47 -6.089859435714609e-20

R25_48 V25 V48 -3415.4745556988164
L25_48 V25 V48 -2.7379082267875795e-12
C25_48 V25 V48 -1.1472772551247215e-19

R25_49 V25 V49 -553.0443463622914
L25_49 V25 V49 -2.4274080293617372e-12
C25_49 V25 V49 -1.3659966202660217e-19

R25_50 V25 V50 10185.064287753725
L25_50 V25 V50 -2.8689779178527683e-12
C25_50 V25 V50 -1.5720683940414356e-19

R25_51 V25 V51 55478.47616662476
L25_51 V25 V51 -3.133634911030504e-12
C25_51 V25 V51 -5.885066874824875e-20

R25_52 V25 V52 4534.884501595927
L25_52 V25 V52 -4.1545595708598594e-12
C25_52 V25 V52 -5.99072928400861e-20

R25_53 V25 V53 -914.8799928118765
L25_53 V25 V53 -2.394600278575385e-12
C25_53 V25 V53 2.5164107303944223e-19

R25_54 V25 V54 -3946.760392488288
L25_54 V25 V54 -7.050573295938234e-12
C25_54 V25 V54 1.0469740304711158e-19

R25_55 V25 V55 -3285.213005360598
L25_55 V25 V55 -4.487642785976297e-12
C25_55 V25 V55 2.974991686492758e-20

R25_56 V25 V56 -7492.122532991979
L25_56 V25 V56 -1.694502874352813e-11
C25_56 V25 V56 9.007747810049397e-20

R25_57 V25 V57 5780.0552525835765
L25_57 V25 V57 6.885060725234674e-13
C25_57 V25 V57 2.8601010109039867e-19

R25_58 V25 V58 2899.1262556037004
L25_58 V25 V58 2.0376253391759295e-12
C25_58 V25 V58 1.34730883697916e-19

R25_59 V25 V59 1647.0357872771606
L25_59 V25 V59 1.92184242514497e-12
C25_59 V25 V59 2.5416092650413377e-20

R25_60 V25 V60 1135.694433485058
L25_60 V25 V60 1.2321914006102273e-12
C25_60 V25 V60 7.770199888457322e-20

R25_61 V25 V61 3965.252373354443
L25_61 V25 V61 -1.14924808366422e-12
C25_61 V25 V61 -3.5854988315216763e-19

R25_62 V25 V62 13491.21747226875
L25_62 V25 V62 7.095491951521781e-11
C25_62 V25 V62 -1.1132540410077045e-19

R25_63 V25 V63 12365.717568123842
L25_63 V25 V63 3.174335093617669e-12
C25_63 V25 V63 9.160279918303386e-20

R25_64 V25 V64 -18479.775105328546
L25_64 V25 V64 6.997557772640172e-12
C25_64 V25 V64 3.318916093881735e-20

R25_65 V25 V65 -784.163323757667
L25_65 V25 V65 -3.0694799249062712e-12
C25_65 V25 V65 -5.227226986287503e-20

R25_66 V25 V66 6308.458333622977
L25_66 V25 V66 -4.7422424119600325e-11
C25_66 V25 V66 5.218614214747545e-21

R25_67 V25 V67 7655.45137596589
L25_67 V25 V67 -5.002423708875089e-12
C25_67 V25 V67 -3.3764773134827674e-21

R25_68 V25 V68 43426.83979279399
L25_68 V25 V68 -1.9192885804936667e-12
C25_68 V25 V68 -9.326223356726969e-20

R25_69 V25 V69 -1166.9245115158192
L25_69 V25 V69 -1.4391284931167907e-12
C25_69 V25 V69 -1.9784026855093816e-19

R25_70 V25 V70 124350.71842473454
L25_70 V25 V70 -6.73736891925096e-12
C25_70 V25 V70 1.6455392522903086e-20

R25_71 V25 V71 -14002.99476880779
L25_71 V25 V71 -2.326050207284898e-12
C25_71 V25 V71 -1.663815662993775e-19

R25_72 V25 V72 -12127.917811481962
L25_72 V25 V72 -2.5326648193708427e-12
C25_72 V25 V72 -1.2776088059593858e-19

R25_73 V25 V73 -1766.7594108090202
L25_73 V25 V73 -3.632339545921139e-11
C25_73 V25 V73 2.2787230629840152e-19

R25_74 V25 V74 -6168.7054956352185
L25_74 V25 V74 -2.387850906286188e-11
C25_74 V25 V74 -3.5602096115912327e-20

R25_75 V25 V75 -11408.19218987211
L25_75 V25 V75 3.74332849758282e-12
C25_75 V25 V75 6.241011798991987e-20

R25_76 V25 V76 4727.687639899749
L25_76 V25 V76 1.763772119423655e-12
C25_76 V25 V76 1.4823871966917855e-19

R25_77 V25 V77 3802.1470179016796
L25_77 V25 V77 9.004509794713494e-13
C25_77 V25 V77 3.2826947532905435e-19

R25_78 V25 V78 -11877.915780637957
L25_78 V25 V78 5.688909621833247e-12
C25_78 V25 V78 9.468186043074503e-20

R25_79 V25 V79 6081.038738595351
L25_79 V25 V79 3.056490677675842e-12
C25_79 V25 V79 1.104282776798324e-19

R25_80 V25 V80 8098.060525755183
L25_80 V25 V80 3.513194993278002e-12
C25_80 V25 V80 7.217632585228274e-20

R25_81 V25 V81 -444.1367262705525
L25_81 V25 V81 -8.967360550789168e-13
C25_81 V25 V81 -5.016356787906311e-19

R25_82 V25 V82 2733.2938875306336
L25_82 V25 V82 1.4062301380201004e-11
C25_82 V25 V82 -1.4689632078095e-20

R25_83 V25 V83 1687.6538157279042
L25_83 V25 V83 3.0682949275049774e-11
C25_83 V25 V83 4.318828709824983e-21

R25_84 V25 V84 1699.7827643108803
L25_84 V25 V84 -9.914783263332643e-11
C25_84 V25 V84 -5.589633801325854e-20

R25_85 V25 V85 22979.81583550496
L25_85 V25 V85 -9.974331675072719e-12
C25_85 V25 V85 6.872691614307387e-20

R25_86 V25 V86 1488.3584506408752
L25_86 V25 V86 -3.693178449482434e-12
C25_86 V25 V86 -1.1701961173497843e-19

R25_87 V25 V87 7944.882794188884
L25_87 V25 V87 -7.858650684644322e-12
C25_87 V25 V87 -6.798531888441158e-20

R25_88 V25 V88 7957.831259840374
L25_88 V25 V88 -3.669788696191606e-12
C25_88 V25 V88 -7.304421491784538e-20

R25_89 V25 V89 -1295.4145831668254
L25_89 V25 V89 -1.095758749475509e-12
C25_89 V25 V89 -1.5481319193669495e-19

R25_90 V25 V90 -2421.335585862252
L25_90 V25 V90 2.022049607431285e-11
C25_90 V25 V90 4.784678420040828e-20

R25_91 V25 V91 -3880.6553534077284
L25_91 V25 V91 -2.350896268146673e-12
C25_91 V25 V91 -1.5035880885428339e-19

R25_92 V25 V92 115304.82841055747
L25_92 V25 V92 -4.934795658499925e-12
C25_92 V25 V92 -6.07413719272256e-20

R25_93 V25 V93 -1088.7233989558476
L25_93 V25 V93 1.4891609428676287e-12
C25_93 V25 V93 1.5203942333101185e-19

R25_94 V25 V94 -2361.148196371436
L25_94 V25 V94 4.502827405914206e-12
C25_94 V25 V94 7.297246999547941e-20

R25_95 V25 V95 37921.98997646172
L25_95 V25 V95 2.678737562947514e-12
C25_95 V25 V95 1.4492929169624994e-19

R25_96 V25 V96 -1267648.3477222784
L25_96 V25 V96 1.911617782994996e-12
C25_96 V25 V96 1.6231518607614646e-19

R25_97 V25 V97 -864.1117359066807
L25_97 V25 V97 1.4483162441322825e-12
C25_97 V25 V97 3.5995187445392424e-19

R25_98 V25 V98 842.8917319346024
L25_98 V25 V98 -5.60718780054857e-12
C25_98 V25 V98 -5.85535622803778e-20

R25_99 V25 V99 930.2628420983461
L25_99 V25 V99 2.7769819433301104e-12
C25_99 V25 V99 7.775803322220416e-20

R25_100 V25 V100 932.8550166083514
L25_100 V25 V100 2.949725140213335e-12
C25_100 V25 V100 4.900227083856899e-20

R25_101 V25 V101 4299.5498562332605
L25_101 V25 V101 -9.42489101807825e-13
C25_101 V25 V101 -4.3123311293984684e-19

R25_102 V25 V102 6184.244766568755
L25_102 V25 V102 1.1494972007031495e-11
C25_102 V25 V102 7.268420301706178e-20

R25_103 V25 V103 -42729.31788695715
L25_103 V25 V103 -6.443327568497179e-12
C25_103 V25 V103 -1.7815364135215664e-20

R25_104 V25 V104 5798.776755542875
L25_104 V25 V104 -5.3402021297941876e-12
C25_104 V25 V104 -6.848057754038723e-20

R25_105 V25 V105 -390.18844791927194
L25_105 V25 V105 -1.7663140655413394e-12
C25_105 V25 V105 -7.573445677170538e-20

R25_106 V25 V106 -34468.989460062265
L25_106 V25 V106 5.764695273752945e-12
C25_106 V25 V106 -8.571437259691067e-20

R25_107 V25 V107 -17108.731378185068
L25_107 V25 V107 -5.6897989369885706e-12
C25_107 V25 V107 -1.3204972882959137e-19

R25_108 V25 V108 -4969.26613880965
L25_108 V25 V108 -2.534585345217843e-12
C25_108 V25 V108 -1.1747443447079597e-19

R25_109 V25 V109 4232.708218675642
L25_109 V25 V109 -9.952411837492977e-12
C25_109 V25 V109 7.789192256195098e-20

R25_110 V25 V110 6524.629298428552
L25_110 V25 V110 -5.594385853619874e-12
C25_110 V25 V110 7.279919462107826e-21

R25_111 V25 V111 -18996.58467274285
L25_111 V25 V111 -4.7813611279208426e-12
C25_111 V25 V111 -7.555485451754368e-20

R25_112 V25 V112 10543.322864720758
L25_112 V25 V112 9.381679217799792e-12
C25_112 V25 V112 3.480105790313644e-21

R25_113 V25 V113 -1451.714368176284
L25_113 V25 V113 2.949805104944903e-12
C25_113 V25 V113 1.0310692602384777e-19

R25_114 V25 V114 3189.3497451357275
L25_114 V25 V114 1.1441974021346477e-11
C25_114 V25 V114 8.359527808924707e-20

R25_115 V25 V115 2096.007219801414
L25_115 V25 V115 2.847362333096292e-12
C25_115 V25 V115 2.2079143109839024e-19

R25_116 V25 V116 3303.672589612322
L25_116 V25 V116 2.30782228176369e-12
C25_116 V25 V116 2.0678858303430417e-19

R25_117 V25 V117 -1512.9275831742777
L25_117 V25 V117 1.370954820565765e-12
C25_117 V25 V117 2.0406923373277113e-19

R25_118 V25 V118 -4431.108966524236
L25_118 V25 V118 2.4562744493885324e-11
C25_118 V25 V118 -4.2683693674187357e-20

R25_119 V25 V119 8494.230482218456
L25_119 V25 V119 -8.835075938150437e-12
C25_119 V25 V119 -6.143562944410075e-20

R25_120 V25 V120 3337.9386609383355
L25_120 V25 V120 -4.057154321183252e-12
C25_120 V25 V120 -6.99054389302745e-20

R25_121 V25 V121 -3539.546950848929
L25_121 V25 V121 -9.02055456636238e-13
C25_121 V25 V121 -3.7066763357957464e-19

R25_122 V25 V122 4246.938445035002
L25_122 V25 V122 -4.2634694700638207e-10
C25_122 V25 V122 -5.383824021070052e-21

R25_123 V25 V123 -3651.776358493705
L25_123 V25 V123 7.237952188019482e-12
C25_123 V25 V123 -2.638516398491135e-20

R25_124 V25 V124 -3085.2109218599417
L25_124 V25 V124 2.8762035288259863e-11
C25_124 V25 V124 -1.156019596330355e-19

R25_125 V25 V125 -466.44060460514714
L25_125 V25 V125 -9.077903107300975e-13
C25_125 V25 V125 -1.9145379573360284e-19

R25_126 V25 V126 4621.590648106576
L25_126 V25 V126 -3.0722478161444462e-12
C25_126 V25 V126 -1.2172609812227535e-19

R25_127 V25 V127 3247.6305722277543
L25_127 V25 V127 -1.0378595204262503e-11
C25_127 V25 V127 -3.5235879875177524e-20

R25_128 V25 V128 432085.550504722
L25_128 V25 V128 -5.052083768914512e-12
C25_128 V25 V128 -3.80734554996891e-20

R25_129 V25 V129 1927.7297686930317
L25_129 V25 V129 1.233460344874933e-12
C25_129 V25 V129 2.964945994877124e-19

R25_130 V25 V130 -15225.86106272457
L25_130 V25 V130 3.261056065405782e-12
C25_130 V25 V130 1.4588190521068994e-19

R25_131 V25 V131 -4876.941340846033
L25_131 V25 V131 -2.898744037751784e-11
C25_131 V25 V131 6.43900782465738e-20

R25_132 V25 V132 3875.3463305519067
L25_132 V25 V132 5.724568732752199e-12
C25_132 V25 V132 1.7961470478400702e-19

R25_133 V25 V133 841.8649091276387
L25_133 V25 V133 2.2666996719142664e-12
C25_133 V25 V133 -3.338287790921728e-20

R25_134 V25 V134 2092.7145534142683
L25_134 V25 V134 3.748461942106667e-12
C25_134 V25 V134 -1.373629041203148e-21

R25_135 V25 V135 -5022.01773982238
L25_135 V25 V135 7.281642201903389e-12
C25_135 V25 V135 -7.146619397859827e-21

R25_136 V25 V136 -2000.1077772988717
L25_136 V25 V136 5.1300060313747696e-12
C25_136 V25 V136 -3.2504880595822344e-20

R25_137 V25 V137 -577.5110397406612
L25_137 V25 V137 5.22239354692712e-12
C25_137 V25 V137 1.4686471040151174e-19

R25_138 V25 V138 -1363.833344237626
L25_138 V25 V138 -2.49280630225651e-12
C25_138 V25 V138 -6.889145670647197e-20

R25_139 V25 V139 1716.9894830734872
L25_139 V25 V139 -2.605799697592763e-12
C25_139 V25 V139 -4.8228429324750715e-20

R25_140 V25 V140 1657.7158096015805
L25_140 V25 V140 -4.399606028801732e-12
C25_140 V25 V140 4.151917252642644e-20

R25_141 V25 V141 1909.4215468483249
L25_141 V25 V141 -1.432668808058309e-12
C25_141 V25 V141 -2.3004908049646694e-19

R25_142 V25 V142 984.3850418768079
L25_142 V25 V142 -6.657414780730083e-11
C25_142 V25 V142 -3.2025591659916213e-21

R25_143 V25 V143 3718.745787729565
L25_143 V25 V143 1.930471090421615e-12
C25_143 V25 V143 6.822955472064504e-20

R25_144 V25 V144 1214.317972024009
L25_144 V25 V144 6.959817389697489e-12
C25_144 V25 V144 -7.452036543943151e-20

R25_145 V25 V145 -609.1582466926604
L25_145 V25 V145 -1.4108203918940057e-12
C25_145 V25 V145 -2.1857526050560126e-19

R25_146 V25 V146 9259.583647950583
L25_146 V25 V146 1.8980940135031685e-12
C25_146 V25 V146 8.852337882104125e-20

R25_147 V25 V147 -11224.637283567998
L25_147 V25 V147 -7.88996367085057e-12
C25_147 V25 V147 -9.593718074833649e-20

R25_148 V25 V148 -732.0175585864
L25_148 V25 V148 -3.802976018668389e-12
C25_148 V25 V148 -1.0446130987454781e-19

R25_149 V25 V149 310.29911521504977
L25_149 V25 V149 3.060136214802653e-12
C25_149 V25 V149 1.489064207285086e-19

R25_150 V25 V150 -752.1319074234098
L25_150 V25 V150 -1.7874792281061926e-12
C25_150 V25 V150 -1.3295599682673244e-19

R25_151 V25 V151 -755.2739854921903
L25_151 V25 V151 -1.39334020957649e-12
C25_151 V25 V151 -8.033252342574515e-20

R25_152 V25 V152 1972.907513792975
L25_152 V25 V152 -1.0714921583336781e-11
C25_152 V25 V152 5.3023399893616237e-20

R25_153 V25 V153 -408.1235928785012
L25_153 V25 V153 1.4313538995460895e-12
C25_153 V25 V153 2.866464464809929e-19

R25_154 V25 V154 2052.3484535200996
L25_154 V25 V154 2.2046767012832262e-11
C25_154 V25 V154 6.609777444278729e-20

R25_155 V25 V155 483.95388877576715
L25_155 V25 V155 8.199504529042056e-12
C25_155 V25 V155 2.496522208528085e-20

R25_156 V25 V156 -4402.663348926652
L25_156 V25 V156 3.1188433049265796e-11
C25_156 V25 V156 9.843556659711973e-20

R25_157 V25 V157 -425.1730207060037
L25_157 V25 V157 -1.2807868545135707e-10
C25_157 V25 V157 9.537312217794652e-21

R25_158 V25 V158 1919.7957469549506
L25_158 V25 V158 3.3647183767995166e-12
C25_158 V25 V158 6.691725333791119e-21

R25_159 V25 V159 -3570.2103599981237
L25_159 V25 V159 1.3051388164917377e-12
C25_159 V25 V159 1.471721897652903e-19

R25_160 V25 V160 1077.9508089034316
L25_160 V25 V160 1.3815931843475545e-12
C25_160 V25 V160 4.749362389085085e-20

R25_161 V25 V161 -17618.496054328378
L25_161 V25 V161 -1.4357415208820107e-12
C25_161 V25 V161 -2.9845782268327415e-19

R25_162 V25 V162 28998.023497017028
L25_162 V25 V162 5.596001139370399e-12
C25_162 V25 V162 1.2579260178633192e-19

R25_163 V25 V163 1194.58776402327
L25_163 V25 V163 2.2105699849221263e-12
C25_163 V25 V163 1.0167420803910372e-19

R25_164 V25 V164 -5929.363810618131
L25_164 V25 V164 -2.212198255905805e-11
C25_164 V25 V164 9.34085060651766e-21

R25_165 V25 V165 -488.6584664893251
L25_165 V25 V165 -6.949881954754815e-13
C25_165 V25 V165 -1.7811583310431095e-19

R25_166 V25 V166 3880.8456551214367
L25_166 V25 V166 -1.1419978171369204e-12
C25_166 V25 V166 -1.6575223773192984e-19

R25_167 V25 V167 -2378.718501543236
L25_167 V25 V167 -1.2064267818296574e-12
C25_167 V25 V167 -1.8935217226801855e-19

R25_168 V25 V168 777.7653262300621
L25_168 V25 V168 -1.2378425253587447e-12
C25_168 V25 V168 -2.4250590922086477e-19

R25_169 V25 V169 -2656.0026889415262
L25_169 V25 V169 9.362268211636301e-13
C25_169 V25 V169 2.663735781885662e-19

R25_170 V25 V170 -821.9461185282254
L25_170 V25 V170 -8.452693013286925e-11
C25_170 V25 V170 -5.462567547969862e-20

R25_171 V25 V171 -1011.8957047273966
L25_171 V25 V171 -1.8879743849742838e-12
C25_171 V25 V171 -9.252245569728555e-20

R25_172 V25 V172 -1080.4894880811016
L25_172 V25 V172 -2.1088720943873614e-11
C25_172 V25 V172 5.513524511543316e-20

R25_173 V25 V173 -1117.6899725390135
L25_173 V25 V173 1.4445784240612942e-12
C25_173 V25 V173 1.9190540365790473e-19

R25_174 V25 V174 630.7195999464095
L25_174 V25 V174 6.777286216060315e-13
C25_174 V25 V174 2.892688352280502e-19

R25_175 V25 V175 825.203629054643
L25_175 V25 V175 7.862416973865436e-13
C25_175 V25 V175 2.5002532807453197e-19

R25_176 V25 V176 1050.9227560459285
L25_176 V25 V176 6.698477259316165e-13
C25_176 V25 V176 3.1490201423216497e-19

R25_177 V25 V177 2076.364505809685
L25_177 V25 V177 -2.0944233498376438e-12
C25_177 V25 V177 -1.4925103812153703e-19

R25_178 V25 V178 -1574.6830462915232
L25_178 V25 V178 -3.588726742138302e-12
C25_178 V25 V178 -3.060596643239449e-20

R25_179 V25 V179 4803.221846279077
L25_179 V25 V179 -8.77511155951722e-12
C25_179 V25 V179 -1.5944981756721874e-20

R25_180 V25 V180 -2283.3531028041875
L25_180 V25 V180 -2.2261005082486534e-12
C25_180 V25 V180 -1.0705041225071328e-19

R25_181 V25 V181 635.1702748353641
L25_181 V25 V181 -1.8362322806772263e-12
C25_181 V25 V181 -4.472996772973798e-19

R25_182 V25 V182 -1994.763171706149
L25_182 V25 V182 -1.398432308356244e-12
C25_182 V25 V182 -7.577643527904981e-20

R25_183 V25 V183 -1874.36378232601
L25_183 V25 V183 -6.540475811344216e-12
C25_183 V25 V183 -1.710605764280407e-20

R25_184 V25 V184 -2033.1242493647367
L25_184 V25 V184 -1.8128207549956737e-12
C25_184 V25 V184 -6.193472986002167e-20

R25_185 V25 V185 -267.6900073049596
L25_185 V25 V185 -2.4528286752290384e-12
C25_185 V25 V185 3.4362551003153017e-19

R25_186 V25 V186 807.6746076371629
L25_186 V25 V186 -1.377565304148731e-12
C25_186 V25 V186 -1.7917069351637176e-19

R25_187 V25 V187 77298.91245175025
L25_187 V25 V187 -2.5051995239527514e-12
C25_187 V25 V187 -4.6996332132717955e-20

R25_188 V25 V188 3179.701354138082
L25_188 V25 V188 -2.352655950108454e-12
C25_188 V25 V188 -1.0024993688946159e-19

R25_189 V25 V189 346.42025617029026
L25_189 V25 V189 8.856425030059046e-13
C25_189 V25 V189 1.050862291349897e-19

R25_190 V25 V190 -3215.0443023775224
L25_190 V25 V190 1.7267819785611993e-12
C25_190 V25 V190 4.293968323696912e-20

R25_191 V25 V191 -883.0792472504988
L25_191 V25 V191 -1.489549056141136e-11
C25_191 V25 V191 -1.8151408027993572e-20

R25_192 V25 V192 -1188.3313342977058
L25_192 V25 V192 1.5805403877768146e-12
C25_192 V25 V192 1.602452177934705e-19

R25_193 V25 V193 1043.4312311485464
L25_193 V25 V193 4.079878210781984e-12
C25_193 V25 V193 4.8423116334611565e-20

R25_194 V25 V194 -1067.4397686394716
L25_194 V25 V194 8.810376119115496e-13
C25_194 V25 V194 2.27177820145652e-19

R25_195 V25 V195 4456.291083994769
L25_195 V25 V195 3.1067993230531634e-12
C25_195 V25 V195 2.5923133917530797e-20

R25_196 V25 V196 14399.174126415739
L25_196 V25 V196 1.4301438891922656e-12
C25_196 V25 V196 9.339145949868236e-20

R25_197 V25 V197 -585.8667220521403
L25_197 V25 V197 -1.6329284827401783e-12
C25_197 V25 V197 -1.8701181049406424e-19

R25_198 V25 V198 1297.5981320929664
L25_198 V25 V198 -1.5930947599689828e-12
C25_198 V25 V198 -5.0431935262083304e-20

R25_199 V25 V199 707.6084838287017
L25_199 V25 V199 -2.0799746788869498e-11
C25_199 V25 V199 1.1006529844578643e-19

R25_200 V25 V200 633.5001957767812
L25_200 V25 V200 -1.2092510861964998e-12
C25_200 V25 V200 -1.274796500790589e-19

R26_26 V26 0 179.6711015584109
L26_26 V26 0 2.8185945445541526e-13
C26_26 V26 0 2.0698440398784045e-18

R26_27 V26 V27 -4579.7976252045155
L26_27 V26 V27 -1.340001079056442e-12
C26_27 V26 V27 -4.197464333679253e-19

R26_28 V26 V28 -3498.866374274132
L26_28 V26 V28 -9.946521912568339e-13
C26_28 V26 V28 -5.984993950467607e-19

R26_29 V26 V29 -2103.603091895309
L26_29 V26 V29 -1.6438350320109237e-11
C26_29 V26 V29 1.11995284225604e-19

R26_30 V26 V30 -1517.397776590797
L26_30 V26 V30 2.368792106417356e-12
C26_30 V26 V30 6.028294803067849e-19

R26_31 V26 V31 -2188.155189669383
L26_31 V26 V31 3.944330128746659e-12
C26_31 V26 V31 2.3502356463346267e-19

R26_32 V26 V32 -2025.53323211788
L26_32 V26 V32 2.7188627058363008e-12
C26_32 V26 V32 3.6659068604373326e-19

R26_33 V26 V33 -9021.004215190724
L26_33 V26 V33 2.2668724284996296e-11
C26_33 V26 V33 9.552410514755454e-20

R26_34 V26 V34 3447.13243718402
L26_34 V26 V34 7.680288732191193e-13
C26_34 V26 V34 8.001721839760683e-19

R26_35 V26 V35 3421.925320140036
L26_35 V26 V35 3.975602356812243e-12
C26_35 V26 V35 1.4955069319753944e-19

R26_36 V26 V36 2189.8204509716998
L26_36 V26 V36 2.230938309404709e-12
C26_36 V26 V36 2.7404998612761905e-19

R26_37 V26 V37 4260.386033938001
L26_37 V26 V37 3.686428605313997e-12
C26_37 V26 V37 1.319275747693257e-20

R26_38 V26 V38 3593.726851960858
L26_38 V26 V38 -1.6672595381815522e-12
C26_38 V26 V38 -5.88915260962765e-19

R26_39 V26 V39 2500.379763344932
L26_39 V26 V39 -4.753896343101835e-12
C26_39 V26 V39 -1.9645220989084229e-19

R26_40 V26 V40 1889.1415897411052
L26_40 V26 V40 -3.975147843917452e-12
C26_40 V26 V40 -2.6613162426869834e-19

R26_41 V26 V41 -10905.221642992696
L26_41 V26 V41 4.690252465991097e-12
C26_41 V26 V41 5.364579292310535e-20

R26_42 V26 V42 4888.28179046849
L26_42 V26 V42 -2.981859342595999e-11
C26_42 V26 V42 3.764810781577191e-20

R26_43 V26 V43 17695.052328914167
L26_43 V26 V43 4.944764100670551e-12
C26_43 V26 V43 1.5192273176582237e-19

R26_44 V26 V44 42983.990188657306
L26_44 V26 V44 3.763147740071521e-12
C26_44 V26 V44 2.2853919402320307e-19

R26_45 V26 V45 -2624.6033852455853
L26_45 V26 V45 -1.5039659200424085e-12
C26_45 V26 V45 -3.157184342644671e-19

R26_46 V26 V46 -2171.821303854505
L26_46 V26 V46 -2.3449722029729557e-12
C26_46 V26 V46 -2.928908014994907e-19

R26_47 V26 V47 -3168.630629088219
L26_47 V26 V47 -1.6892501921034734e-11
C26_47 V26 V47 -9.36259480828065e-20

R26_48 V26 V48 -2124.2153697194053
L26_48 V26 V48 -5.047574527797822e-12
C26_48 V26 V48 -1.5922365136169106e-19

R26_49 V26 V49 -6178.831513718131
L26_49 V26 V49 -1.511250122117114e-11
C26_49 V26 V49 -1.0580591150075875e-20

R26_50 V26 V50 -5592.92157819528
L26_50 V26 V50 -3.3008475326189698e-12
C26_50 V26 V50 -1.1225605094403435e-19

R26_51 V26 V51 -11017.02692917204
L26_51 V26 V51 -4.212536386077846e-12
C26_51 V26 V51 -9.180825140023122e-20

R26_52 V26 V52 12643.196553465224
L26_52 V26 V52 -4.747577097578486e-12
C26_52 V26 V52 -8.494914971744902e-20

R26_53 V26 V53 -5637.697535231659
L26_53 V26 V53 5.942683731613021e-12
C26_53 V26 V53 3.1391634105309944e-19

R26_54 V26 V54 8316.809729289902
L26_54 V26 V54 1.3646466374300084e-12
C26_54 V26 V54 5.878786216922574e-19

R26_55 V26 V55 8886.081862452866
L26_55 V26 V55 5.1508467724013335e-12
C26_55 V26 V55 1.9532371424164978e-19

R26_56 V26 V56 2739.643109486319
L26_56 V26 V56 2.487683127015831e-12
C26_56 V26 V56 3.4437864823115094e-19

R26_57 V26 V57 56502.05812014839
L26_57 V26 V57 5.792177646995682e-12
C26_57 V26 V57 -1.3643104690327209e-19

R26_58 V26 V58 -16977.902612782033
L26_58 V26 V58 -6.2562726777070114e-12
C26_58 V26 V58 -2.670217744854873e-19

R26_59 V26 V59 5388.958652734293
L26_59 V26 V59 6.973536795267241e-11
C26_59 V26 V59 -9.261695748631167e-20

R26_60 V26 V60 3952.476830684339
L26_60 V26 V60 7.0988456544164305e-12
C26_60 V26 V60 -4.202467026909667e-20

R26_61 V26 V61 155671.47135239554
L26_61 V26 V61 -3.3567234022389705e-12
C26_61 V26 V61 -1.5637449782753667e-19

R26_62 V26 V62 5222.487783162802
L26_62 V26 V62 -3.137091228807773e-12
C26_62 V26 V62 -2.059102739989751e-19

R26_63 V26 V63 -37270.881231143074
L26_63 V26 V63 -1.3484759137317802e-11
C26_63 V26 V63 -1.069059293262503e-19

R26_64 V26 V64 -5910.97963137666
L26_64 V26 V64 -3.4647717373173888e-12
C26_64 V26 V64 -2.4638161977027245e-19

R26_65 V26 V65 -4065.4638164859784
L26_65 V26 V65 4.933052333589249e-11
C26_65 V26 V65 1.718595581156364e-20

R26_66 V26 V66 -3613.418635266416
L26_66 V26 V66 6.2041661000160456e-12
C26_66 V26 V66 5.083384822905333e-20

R26_67 V26 V67 -23415.980712782904
L26_67 V26 V67 4.699548030580794e-12
C26_67 V26 V67 1.672973081885091e-19

R26_68 V26 V68 -5833.413607184161
L26_68 V26 V68 1.1725792151929714e-11
C26_68 V26 V68 9.427790862413197e-20

R26_69 V26 V69 -23460.30858199208
L26_69 V26 V69 -1.2768144174129136e-11
C26_69 V26 V69 1.4228176146819262e-19

R26_70 V26 V70 -11601.091143933838
L26_70 V26 V70 -2.5182973571271784e-12
C26_70 V26 V70 -1.575958672846875e-19

R26_71 V26 V71 -6952.656124962193
L26_71 V26 V71 -1.1210419458440707e-11
C26_71 V26 V71 -7.986820275702588e-21

R26_72 V26 V72 -8777.865882098196
L26_72 V26 V72 6.973616579515936e-12
C26_72 V26 V72 1.6825586459248727e-19

R26_73 V26 V73 -4487.46166730278
L26_73 V26 V73 -6.6867950469079315e-12
C26_73 V26 V73 -7.974592951333102e-20

R26_74 V26 V74 3143.2248857856857
L26_74 V26 V74 1.9090409543912202e-12
C26_74 V26 V74 3.5480643696440627e-19

R26_75 V26 V75 27451.62998927685
L26_75 V26 V75 -3.8874321018232035e-12
C26_75 V26 V75 -1.991966295123922e-19

R26_76 V26 V76 2443.107508761203
L26_76 V26 V76 -1.0779029101829815e-11
C26_76 V26 V76 -7.018770498733456e-20

R26_77 V26 V77 7410.0645402776745
L26_77 V26 V77 2.749659195146887e-12
C26_77 V26 V77 -5.8051265029208146e-21

R26_78 V26 V78 -1991.0149436448073
L26_78 V26 V78 -5.454750714806343e-12
C26_78 V26 V78 -7.566794444494823e-20

R26_79 V26 V79 5162.304490858482
L26_79 V26 V79 6.231152024963803e-12
C26_79 V26 V79 7.482900940125894e-20

R26_80 V26 V80 -41409.477598557416
L26_80 V26 V80 6.40242052249708e-10
C26_80 V26 V80 -8.936254661286734e-20

R26_81 V26 V81 -1782.710134484113
L26_81 V26 V81 -2.0797514364188353e-12
C26_81 V26 V81 -1.7989547004003032e-19

R26_82 V26 V82 5226.508949618842
L26_82 V26 V82 -2.689574437848157e-12
C26_82 V26 V82 -4.455147440189092e-19

R26_83 V26 V83 10390.566157311041
L26_83 V26 V83 3.4762895167171417e-12
C26_83 V26 V83 1.3789670319693377e-19

R26_84 V26 V84 -80550.62723255625
L26_84 V26 V84 4.9900197915425505e-12
C26_84 V26 V84 4.935608342027415e-20

R26_85 V26 V85 7907.075772983911
L26_85 V26 V85 -3.749592667911619e-11
C26_85 V26 V85 -1.6016360992747244e-20

R26_86 V26 V86 8473.251618610768
L26_86 V26 V86 2.9288504300550274e-12
C26_86 V26 V86 2.2962897094589263e-19

R26_87 V26 V87 -5288.780028965905
L26_87 V26 V87 -4.800631180830093e-12
C26_87 V26 V87 -9.751498481353087e-20

R26_88 V26 V88 -8182.264615140092
L26_88 V26 V88 -6.369398144125637e-12
C26_88 V26 V88 1.3420209888659692e-20

R26_89 V26 V89 -100087.39201966263
L26_89 V26 V89 1.1412455603780905e-11
C26_89 V26 V89 2.1046004191636163e-19

R26_90 V26 V90 -4067.2565785176953
L26_90 V26 V90 3.36198434448189e-12
C26_90 V26 V90 4.466041556197533e-19

R26_91 V26 V91 -6911.363756459943
L26_91 V26 V91 -4.761693339687315e-12
C26_91 V26 V91 -7.656230944123846e-20

R26_92 V26 V92 6242.727982994222
L26_92 V26 V92 3.626581018504146e-11
C26_92 V26 V92 2.9613192578701937e-20

R26_93 V26 V93 -2226.75704883084
L26_93 V26 V93 -1.4725841416337154e-11
C26_93 V26 V93 -7.64917969364663e-20

R26_94 V26 V94 3176.7628717686907
L26_94 V26 V94 -3.5634564510510212e-12
C26_94 V26 V94 -4.97881356848632e-19

R26_95 V26 V95 2360.4382219443214
L26_95 V26 V95 6.382430725819127e-12
C26_95 V26 V95 1.9052019227849203e-20

R26_96 V26 V96 2111.6369171787846
L26_96 V26 V96 7.117834926181972e-12
C26_96 V26 V96 -3.5602310218314706e-20

R26_97 V26 V97 9022.818216828373
L26_97 V26 V97 -1.2526581411353367e-11
C26_97 V26 V97 -2.902766996806469e-19

R26_98 V26 V98 -4946.314533539059
L26_98 V26 V98 -2.265433151955383e-12
C26_98 V26 V98 -1.8194431069843516e-19

R26_99 V26 V99 11790.615703984527
L26_99 V26 V99 4.317119395933581e-12
C26_99 V26 V99 1.0931136965705898e-19

R26_100 V26 V100 -4016.1489517027153
L26_100 V26 V100 6.149923327061661e-11
C26_100 V26 V100 1.0860570884425122e-20

R26_101 V26 V101 -35098.73489332405
L26_101 V26 V101 5.225867689377792e-11
C26_101 V26 V101 1.594545363063255e-19

R26_102 V26 V102 -14374.846368960574
L26_102 V26 V102 2.178674629442272e-12
C26_102 V26 V102 6.146819724723935e-19

R26_103 V26 V103 -6986.762260352864
L26_103 V26 V103 -1.896171061312228e-10
C26_103 V26 V103 1.152414708537673e-19

R26_104 V26 V104 -11414.627877087256
L26_104 V26 V104 -2.0416103335677294e-11
C26_104 V26 V104 5.0555762259246244e-20

R26_105 V26 V105 -1680.8522767075015
L26_105 V26 V105 -9.929194143579944e-12
C26_105 V26 V105 1.3493690253988433e-19

R26_106 V26 V106 -4791.352196566359
L26_106 V26 V106 2.983006724711337e-12
C26_106 V26 V106 -1.9218268641347377e-19

R26_107 V26 V107 -9281.476774630339
L26_107 V26 V107 -3.5813972062549755e-12
C26_107 V26 V107 -2.298750612593599e-19

R26_108 V26 V108 4860.974542439012
L26_108 V26 V108 3.0980632372687345e-10
C26_108 V26 V108 2.7091389145838827e-20

R26_109 V26 V109 10834.801944980734
L26_109 V26 V109 -2.456420651489175e-12
C26_109 V26 V109 -2.4673812065860014e-19

R26_110 V26 V110 2515.308383072148
L26_110 V26 V110 -1.1192497017071228e-12
C26_110 V26 V110 -5.169288048358752e-19

R26_111 V26 V111 -3045.6520101804626
L26_111 V26 V111 1.3884749825480696e-11
C26_111 V26 V111 -4.3634336555751175e-20

R26_112 V26 V112 -3139.924559689589
L26_112 V26 V112 1.408670925410633e-11
C26_112 V26 V112 -7.475834221951324e-20

R26_113 V26 V113 -4041.711749847061
L26_113 V26 V113 2.986182553351204e-11
C26_113 V26 V113 -1.2986440276659906e-19

R26_114 V26 V114 4254.709578786486
L26_114 V26 V114 7.725204488627938e-12
C26_114 V26 V114 4.017820492270367e-19

R26_115 V26 V115 1317.2236916959407
L26_115 V26 V115 7.321420390501037e-12
C26_115 V26 V115 2.4063524599986327e-19

R26_116 V26 V116 2510.4868177093163
L26_116 V26 V116 -8.521303066186817e-12
C26_116 V26 V116 1.719074209914733e-20

R26_117 V26 V117 2301.9364519267765
L26_117 V26 V117 1.9787992299479238e-12
C26_117 V26 V117 1.8623998792380508e-19

R26_118 V26 V118 -2416.6844698401146
L26_118 V26 V118 9.252139256813053e-13
C26_118 V26 V118 3.2953202828003376e-19

R26_119 V26 V119 -3262.6516057716062
L26_119 V26 V119 -1.8380202064390562e-11
C26_119 V26 V119 -2.803318739550186e-20

R26_120 V26 V120 -4508.7670743690205
L26_120 V26 V120 -8.352677038874898e-11
C26_120 V26 V120 8.896343874463165e-20

R26_121 V26 V121 -3138.8669837526813
L26_121 V26 V121 -2.6042100992783608e-12
C26_121 V26 V121 1.228833145164272e-19

R26_122 V26 V122 -4657.391604247618
L26_122 V26 V122 -1.1095857663784272e-12
C26_122 V26 V122 -5.713006079173983e-19

R26_123 V26 V123 -2270.690277049141
L26_123 V26 V123 3.7773771443901945e-12
C26_123 V26 V123 1.5145180026709573e-20

R26_124 V26 V124 -2814.163555974611
L26_124 V26 V124 3.6114855148305715e-12
C26_124 V26 V124 -4.39055598031669e-20

R26_125 V26 V125 -896.60918073601
L26_125 V26 V125 -2.4239089649570654e-12
C26_125 V26 V125 -1.4527810628538154e-19

R26_126 V26 V126 -5456.7430543060145
L26_126 V26 V126 -1.230168197394038e-12
C26_126 V26 V126 4.019657534216262e-20

R26_127 V26 V127 2053.7418821869387
L26_127 V26 V127 -2.2578252502398004e-12
C26_127 V26 V127 -1.233318855335288e-19

R26_128 V26 V128 2258.6397291739454
L26_128 V26 V128 -2.452057979847344e-12
C26_128 V26 V128 -9.485572719124965e-20

R26_129 V26 V129 1129.2593119463331
L26_129 V26 V129 -6.967789166491674e-11
C26_129 V26 V129 -3.7120011081360204e-19

R26_130 V26 V130 1102.3667674985445
L26_130 V26 V130 9.048099751563496e-13
C26_130 V26 V130 4.2934653206910736e-19

R26_131 V26 V131 -4225.494415976249
L26_131 V26 V131 5.153932573866943e-12
C26_131 V26 V131 4.8782701226558614e-20

R26_132 V26 V132 -5667.768839933291
L26_132 V26 V132 4.137926300465494e-12
C26_132 V26 V132 9.998640588201759e-20

R26_133 V26 V133 1463.429034778701
L26_133 V26 V133 2.4038715897970996e-12
C26_133 V26 V133 4.484486674534638e-19

R26_134 V26 V134 -1398.5974738264588
L26_134 V26 V134 -1.2825715537435569e-11
C26_134 V26 V134 -4.784794984274038e-19

R26_135 V26 V135 -4383.683160540273
L26_135 V26 V135 1.9100665417829718e-12
C26_135 V26 V135 1.9449013869168436e-19

R26_136 V26 V136 -2320.347209359875
L26_136 V26 V136 2.133251567134446e-12
C26_136 V26 V136 -2.290063184566614e-20

R26_137 V26 V137 -697.2369141848757
L26_137 V26 V137 2.3876852519234324e-12
C26_137 V26 V137 2.701123395219892e-19

R26_138 V26 V138 -5926.13112947457
L26_138 V26 V138 -1.900941650568238e-12
C26_138 V26 V138 2.0423841824469422e-19

R26_139 V26 V139 2273.586034804177
L26_139 V26 V139 -1.3200536230859302e-12
C26_139 V26 V139 -9.336385471182789e-20

R26_140 V26 V140 8643.930611989908
L26_140 V26 V140 -1.1306106029124635e-12
C26_140 V26 V140 7.776164858612801e-20

R26_141 V26 V141 -5545.772004868788
L26_141 V26 V141 -1.3338261886990092e-12
C26_141 V26 V141 -6.579424436491132e-19

R26_142 V26 V142 707.5894276883215
L26_142 V26 V142 -4.022233386493904e-12
C26_142 V26 V142 8.164426237669409e-20

R26_143 V26 V143 -5253.431180942807
L26_143 V26 V143 9.071866157003133e-12
C26_143 V26 V143 -1.8597785411196544e-19

R26_144 V26 V144 1126.3038304050672
L26_144 V26 V144 4.082551896900975e-12
C26_144 V26 V144 -1.1158171920400663e-19

R26_145 V26 V145 885.61681522077
L26_145 V26 V145 -1.783461789143877e-12
C26_145 V26 V145 -1.8677868489485173e-19

R26_146 V26 V146 -2086.2185389686315
L26_146 V26 V146 1.100394148656082e-12
C26_146 V26 V146 1.2125232905743313e-20

R26_147 V26 V147 1104.5967083533567
L26_147 V26 V147 2.8400937067635945e-12
C26_147 V26 V147 9.293036232196672e-20

R26_148 V26 V148 -741.5281953473919
L26_148 V26 V148 3.634350171440465e-11
C26_148 V26 V148 -5.389258399171178e-20

R26_149 V26 V149 2375.5949867473373
L26_149 V26 V149 7.268391665612326e-13
C26_149 V26 V149 8.043673229401815e-19

R26_150 V26 V150 -563.8137457877147
L26_150 V26 V150 4.9698576124123534e-12
C26_150 V26 V150 -5.271776991143111e-19

R26_151 V26 V151 -674.7524697622478
L26_151 V26 V151 -1.9583365495597504e-12
C26_151 V26 V151 5.0413516621035836e-20

R26_152 V26 V152 1283.4317880081937
L26_152 V26 V152 -2.6678300294052804e-12
C26_152 V26 V152 -3.9316780613176684e-21

R26_153 V26 V153 -675.0296358666125
L26_153 V26 V153 6.467300904694248e-12
C26_153 V26 V153 1.287124411128357e-19

R26_154 V26 V154 14198.620179207446
L26_154 V26 V154 -1.347435222646236e-12
C26_154 V26 V154 4.0153675829809956e-19

R26_155 V26 V155 349.8383493478167
L26_155 V26 V155 1.8984826368998566e-11
C26_155 V26 V155 1.3057973118690115e-19

R26_156 V26 V156 -761.5795533134853
L26_156 V26 V156 1.5598178041745606e-10
C26_156 V26 V156 1.0775335601663374e-19

R26_157 V26 V157 -1638.0932081720532
L26_157 V26 V157 -7.514968614781448e-13
C26_157 V26 V157 -7.586885337234924e-19

R26_158 V26 V158 878.8690558509497
L26_158 V26 V158 -5.054843223450028e-12
C26_158 V26 V158 -1.010238327417925e-19

R26_159 V26 V159 -609.394405752925
L26_159 V26 V159 1.3936443757853555e-12
C26_159 V26 V159 8.077697302446955e-20

R26_160 V26 V160 1226.5284993762166
L26_160 V26 V160 1.0517697268949275e-12
C26_160 V26 V160 1.374406912942004e-19

R26_161 V26 V161 1833.7178860680622
L26_161 V26 V161 -3.0551079262711802e-12
C26_161 V26 V161 -1.1517927813182137e-19

R26_162 V26 V162 4549.564762905942
L26_162 V26 V162 8.471462660648108e-13
C26_162 V26 V162 1.4239133419033956e-19

R26_163 V26 V163 -9628.272403957995
L26_163 V26 V163 -3.706345208357745e-12
C26_163 V26 V163 -2.0792515917258944e-19

R26_164 V26 V164 -915.2530238360999
L26_164 V26 V164 -1.9532303886694564e-12
C26_164 V26 V164 -7.145521444745359e-20

R26_165 V26 V165 -1649.0972927400092
L26_165 V26 V165 1.5718685648353664e-12
C26_165 V26 V165 3.853800555128823e-19

R26_166 V26 V166 -413.3661372721955
L26_166 V26 V166 -6.642841913685104e-12
C26_166 V26 V166 -9.074014509785153e-20

R26_167 V26 V167 -5655.387827727208
L26_167 V26 V167 -1.90837578860917e-12
C26_167 V26 V167 -9.662734203881035e-20

R26_168 V26 V168 511.38328461135393
L26_168 V26 V168 -2.4902715071631463e-12
C26_168 V26 V168 -1.9983594320027736e-19

R26_169 V26 V169 -1709.853878114337
L26_169 V26 V169 2.3092328566083106e-12
C26_169 V26 V169 2.702969813214793e-20

R26_170 V26 V170 781.0940315292194
L26_170 V26 V170 -1.1924769157146499e-12
C26_170 V26 V170 1.3635743258618434e-19

R26_171 V26 V171 1153.6788297624998
L26_171 V26 V171 1.5662424223382059e-12
C26_171 V26 V171 3.776796134011392e-19

R26_172 V26 V172 -4807.725686160505
L26_172 V26 V172 1.636001320035921e-12
C26_172 V26 V172 2.8061272605235865e-19

R26_173 V26 V173 6094.485826647092
L26_173 V26 V173 -1.6778717859322367e-12
C26_173 V26 V173 -1.1467894859822805e-19

R26_174 V26 V174 445.0387240282316
L26_174 V26 V174 1.06465991420102e-12
C26_174 V26 V174 -9.536365336827165e-20

R26_175 V26 V175 -1688.6003919413552
L26_175 V26 V175 2.11192967298078e-12
C26_175 V26 V175 6.673504114985335e-20

R26_176 V26 V176 -1146.9908407664473
L26_176 V26 V176 2.957696168334619e-12
C26_176 V26 V176 1.2447146357046275e-19

R26_177 V26 V177 -2535.962305966909
L26_177 V26 V177 -8.206142572186378e-12
C26_177 V26 V177 5.115247254672687e-20

R26_178 V26 V178 -463.22992417746826
L26_178 V26 V178 1.1220272061104819e-11
C26_178 V26 V178 -1.8298332336772422e-19

R26_179 V26 V179 1906.9858088549583
L26_179 V26 V179 -1.4426034555982577e-12
C26_179 V26 V179 -3.5934831036808375e-19

R26_180 V26 V180 7288.791041793714
L26_180 V26 V180 -1.3511823605841441e-12
C26_180 V26 V180 -3.090533890271207e-19

R26_181 V26 V181 2141.008313930644
L26_181 V26 V181 3.4831763469678863e-12
C26_181 V26 V181 -1.9242195542987922e-19

R26_182 V26 V182 4148.476969503081
L26_182 V26 V182 -1.5516345258232984e-11
C26_182 V26 V182 2.660201627567954e-19

R26_183 V26 V183 -1374.2115658533116
L26_183 V26 V183 -1.0035860978764175e-11
C26_183 V26 V183 -8.634031038141838e-20

R26_184 V26 V184 -7980.997277885081
L26_184 V26 V184 3.0830817006809693e-10
C26_184 V26 V184 -3.992564824954934e-21

R26_185 V26 V185 -2127.4979102116454
L26_185 V26 V185 -2.171612139670161e-12
C26_185 V26 V185 5.700779203974233e-20

R26_186 V26 V186 957.7266314924321
L26_186 V26 V186 7.980781312983291e-12
C26_186 V26 V186 1.2154049132384784e-21

R26_187 V26 V187 3593.0523171558534
L26_187 V26 V187 2.614333469902361e-12
C26_187 V26 V187 2.451490426698337e-19

R26_188 V26 V188 1069.3963754424844
L26_188 V26 V188 5.2588076216756634e-12
C26_188 V26 V188 1.6525877214441266e-19

R26_189 V26 V189 71624.05773615946
L26_189 V26 V189 2.234730834441488e-12
C26_189 V26 V189 3.1376355840249294e-19

R26_190 V26 V190 -1533.9072536121337
L26_190 V26 V190 3.336889143033043e-11
C26_190 V26 V190 -3.214505966173918e-19

R26_191 V26 V191 4327.848817238928
L26_191 V26 V191 3.702360409978186e-12
C26_191 V26 V191 2.6756722541215615e-19

R26_192 V26 V192 -2973.849391978991
L26_192 V26 V192 3.090873033970288e-12
C26_192 V26 V192 2.5378442614887705e-19

R26_193 V26 V193 1747.5214119104623
L26_193 V26 V193 3.1843099615115787e-12
C26_193 V26 V193 -1.3302727486172348e-19

R26_194 V26 V194 -65040.49314192007
L26_194 V26 V194 9.181657141248933e-12
C26_194 V26 V194 7.160610955676721e-20

R26_195 V26 V195 -1618.63003380711
L26_195 V26 V195 -2.030927290490716e-12
C26_195 V26 V195 -4.987311759938884e-19

R26_196 V26 V196 -972.8918810691309
L26_196 V26 V196 -3.092726326289841e-12
C26_196 V26 V196 -4.221284909944505e-19

R26_197 V26 V197 -4884.5746928828685
L26_197 V26 V197 -1.3083519473340141e-12
C26_197 V26 V197 -2.812599907777188e-19

R26_198 V26 V198 149199.19169672285
L26_198 V26 V198 -7.475052615527504e-11
C26_198 V26 V198 1.2047108956839969e-20

R26_199 V26 V199 -3812.7259513311
L26_199 V26 V199 -3.806619280144022e-12
C26_199 V26 V199 -2.43227357542903e-19

R26_200 V26 V200 970.3849422440401
L26_200 V26 V200 -2.8060589735871586e-12
C26_200 V26 V200 -1.0487012973581616e-19

R27_27 V27 0 377.139239786758
L27_27 V27 0 2.541918289614486e-13
C27_27 V27 0 1.853134903574287e-18

R27_28 V27 V28 -3388.5990000448646
L27_28 V27 V28 -8.075260542376684e-13
C27_28 V27 V28 -6.56843355008615e-19

R27_29 V27 V29 -4155.368365140829
L27_29 V27 V29 -2.910268256695352e-12
C27_29 V27 V29 -2.469584046468838e-21

R27_30 V27 V30 -6808.390301546525
L27_30 V27 V30 1.9389495896822244e-11
C27_30 V27 V30 1.15725862938011e-19

R27_31 V27 V31 -2519.3985889678743
L27_31 V27 V31 -2.1478502849860762e-11
C27_31 V27 V31 2.9765821105195006e-19

R27_32 V27 V32 -3133.103305521706
L27_32 V27 V32 1.330560597371138e-11
C27_32 V27 V32 2.6806518985636315e-19

R27_33 V27 V33 -77595.22131112024
L27_33 V27 V33 4.5630619746342465e-12
C27_33 V27 V33 1.3860619787959927e-19

R27_34 V27 V34 9431.023847742865
L27_34 V27 V34 2.3647804806450535e-12
C27_34 V27 V34 2.3828893237927326e-19

R27_35 V27 V35 3382.062221282587
L27_35 V27 V35 6.518106782769693e-13
C27_35 V27 V35 9.034827916308847e-19

R27_36 V27 V36 3074.5121933833857
L27_36 V27 V36 1.4339516301689407e-12
C27_36 V27 V36 3.917684823511852e-19

R27_37 V27 V37 6371.566454337069
L27_37 V27 V37 2.0544273343907887e-12
C27_37 V27 V37 1.3568317044984163e-19

R27_38 V27 V38 10253.002105653559
L27_38 V27 V38 1.032716817410046e-11
C27_38 V27 V38 -5.458304192624395e-21

R27_39 V27 V39 4217.3235952181
L27_39 V27 V39 -2.0463021213801804e-12
C27_39 V27 V39 -6.073539670469932e-19

R27_40 V27 V40 3064.186272959506
L27_40 V27 V40 -6.97159043694033e-12
C27_40 V27 V40 -3.02717652447302e-19

R27_41 V27 V41 -16355.893432969298
L27_41 V27 V41 1.6345186716203923e-11
C27_41 V27 V41 -4.7872207695715076e-20

R27_42 V27 V42 -42028.04027891436
L27_42 V27 V42 -7.917628347510353e-11
C27_42 V27 V42 -4.470485192983336e-20

R27_43 V27 V43 5924.213147088467
L27_43 V27 V43 4.722772527945067e-12
C27_43 V27 V43 9.117489475528758e-20

R27_44 V27 V44 15689.921431257788
L27_44 V27 V44 4.1242420224381414e-12
C27_44 V27 V44 2.0895098606187893e-19

R27_45 V27 V45 -4317.686534893283
L27_45 V27 V45 -1.393667642179463e-12
C27_45 V27 V45 -3.109020720026011e-19

R27_46 V27 V46 -5054.674009277199
L27_46 V27 V46 -2.398659213290887e-12
C27_46 V27 V46 -2.5568321465892904e-19

R27_47 V27 V47 -4190.970099226691
L27_47 V27 V47 -1.6764311761627488e-12
C27_47 V27 V47 -2.2806113585738434e-19

R27_48 V27 V48 -2839.489844245487
L27_48 V27 V48 -1.938519233011079e-12
C27_48 V27 V48 -2.5227519991898396e-19

R27_49 V27 V49 -14883.059336793822
L27_49 V27 V49 -2.3702949567676967e-11
C27_49 V27 V49 -2.499531157607646e-20

R27_50 V27 V50 -29668.674923385315
L27_50 V27 V50 -2.442166904828414e-11
C27_50 V27 V50 -2.6101753367124688e-20

R27_51 V27 V51 -4916.721889367382
L27_51 V27 V51 -6.42864061178193e-12
C27_51 V27 V51 -4.592623802534273e-20

R27_52 V27 V52 -169980.02623071522
L27_52 V27 V52 6.071046135755867e-11
C27_52 V27 V52 4.04104773425928e-20

R27_53 V27 V53 -16149.988028582195
L27_53 V27 V53 7.344245304514755e-12
C27_53 V27 V53 2.46380149160264e-19

R27_54 V27 V54 11518.171312723101
L27_54 V27 V54 2.4592460349926918e-12
C27_54 V27 V54 3.072445651032344e-19

R27_55 V27 V55 -33716.54363021078
L27_55 V27 V55 1.6149551846945272e-12
C27_55 V27 V55 4.751425844029949e-19

R27_56 V27 V56 3970.626375023896
L27_56 V27 V56 2.074790159171349e-12
C27_56 V27 V56 3.391698558722561e-19

R27_57 V27 V57 61426.33690102527
L27_57 V27 V57 3.3607061628682334e-12
C27_57 V27 V57 -2.8238601711505675e-20

R27_58 V27 V58 -8684.37702078925
L27_58 V27 V58 -1.611778586241498e-11
C27_58 V27 V58 -8.381672300361539e-20

R27_59 V27 V59 3625.554656533713
L27_59 V27 V59 -3.827817833590813e-12
C27_59 V27 V59 -3.93999545412323e-19

R27_60 V27 V60 5422.236765600067
L27_60 V27 V60 -1.9903944060592698e-11
C27_60 V27 V60 -1.6097994404367278e-19

R27_61 V27 V61 -73221.87368422838
L27_61 V27 V61 -3.255298861918948e-12
C27_61 V27 V61 -1.6519618190926277e-19

R27_62 V27 V62 16338.576463900377
L27_62 V27 V62 -3.929407198922561e-12
C27_62 V27 V62 -2.5267469962006515e-19

R27_63 V27 V63 -13883.015505091465
L27_63 V27 V63 1.993195205405785e-11
C27_63 V27 V63 6.528844437089042e-20

R27_64 V27 V64 -8508.27442237646
L27_64 V27 V64 -2.0093866249287755e-11
C27_64 V27 V64 -4.023015495308373e-20

R27_65 V27 V65 -8161.920902952337
L27_65 V27 V65 -5.309713619748401e-12
C27_65 V27 V65 -1.2128023218143766e-19

R27_66 V27 V66 -12209.625947085826
L27_66 V27 V66 7.688686871029305e-11
C27_66 V27 V66 2.481118718117866e-20

R27_67 V27 V67 -44546.34496542588
L27_67 V27 V67 3.5735703962116315e-12
C27_67 V27 V67 1.8338496195299927e-19

R27_68 V27 V68 -7946.678744275981
L27_68 V27 V68 -2.217072099198477e-11
C27_68 V27 V68 2.4005226608668272e-20

R27_69 V27 V69 -19253.24227598701
L27_69 V27 V69 -5.66824075627774e-11
C27_69 V27 V69 1.512426118895794e-19

R27_70 V27 V70 35586.46887167148
L27_70 V27 V70 5.4177772109256725e-12
C27_70 V27 V70 1.7115532016715442e-19

R27_71 V27 V71 -5115.372908879933
L27_71 V27 V71 -1.0255925938705846e-12
C27_71 V27 V71 -4.6412413042446765e-19

R27_72 V27 V72 -7931.3184587321875
L27_72 V27 V72 -4.79599144359841e-12
C27_72 V27 V72 -1.795742055356865e-20

R27_73 V27 V73 -12017.030782436657
L27_73 V27 V73 -7.118776839230839e-12
C27_73 V27 V73 -6.036549682848153e-20

R27_74 V27 V74 13685.557411053951
L27_74 V27 V74 -1.0714320135484921e-11
C27_74 V27 V74 -1.309737542792796e-19

R27_75 V27 V75 7609.1308410646925
L27_75 V27 V75 1.3093089649586383e-12
C27_75 V27 V75 3.637283870748006e-19

R27_76 V27 V76 3085.7743690042184
L27_76 V27 V76 3.167261250604981e-12
C27_76 V27 V76 1.3508470174104012e-19

R27_77 V27 V77 8167.4469417407045
L27_77 V27 V77 2.5784846609621432e-12
C27_77 V27 V77 3.3296668650222117e-20

R27_78 V27 V78 -8309.574390563426
L27_78 V27 V78 5.183265293431945e-12
C27_78 V27 V78 2.222914531450818e-19

R27_79 V27 V79 80905.20310840209
L27_79 V27 V79 1.8642967275939507e-11
C27_79 V27 V79 1.1797431353930213e-20

R27_80 V27 V80 230410.45932062573
L27_80 V27 V80 1.1802218296683877e-11
C27_80 V27 V80 -9.792975554838833e-21

R27_81 V27 V81 -3211.0361846140536
L27_81 V27 V81 -2.446663913560946e-12
C27_81 V27 V81 -1.4713280143272142e-19

R27_82 V27 V82 13875.558629387995
L27_82 V27 V82 -3.783010154108883e-12
C27_82 V27 V82 -2.519019135282926e-19

R27_83 V27 V83 20227.74889237551
L27_83 V27 V83 -2.5553288080175413e-12
C27_83 V27 V83 -2.8340221742117844e-19

R27_84 V27 V84 -33971.933549361805
L27_84 V27 V84 -5.7834882240045e-12
C27_84 V27 V84 -1.2326326600528722e-19

R27_85 V27 V85 49578.69961648077
L27_85 V27 V85 -2.7491799588305846e-12
C27_85 V27 V85 -2.0226746503867432e-19

R27_86 V27 V86 -9224.354152945982
L27_86 V27 V86 -2.0769329126427773e-12
C27_86 V27 V86 -3.057828143871317e-19

R27_87 V27 V87 3170.9041289922125
L27_87 V27 V87 1.1249477944537216e-12
C27_87 V27 V87 5.76058733317942e-19

R27_88 V27 V88 -14990.665839232852
L27_88 V27 V88 1.8340793676830303e-11
C27_88 V27 V88 1.3878610763972371e-19

R27_89 V27 V89 11155.54624038178
L27_89 V27 V89 3.339688344203886e-12
C27_89 V27 V89 2.7261442341856415e-19

R27_90 V27 V90 10012.450885730455
L27_90 V27 V90 9.57746131772369e-13
C27_90 V27 V90 7.025952515112226e-19

R27_91 V27 V91 -993.4986908402304
L27_91 V27 V91 -6.031232338418871e-13
C27_91 V27 V91 -8.308326608152852e-19

R27_92 V27 V92 -34092.853845517544
L27_92 V27 V92 -3.5669646089673243e-12
C27_92 V27 V92 -1.569653394654341e-19

R27_93 V27 V93 -4047.3397170290464
L27_93 V27 V93 4.605432829111378e-12
C27_93 V27 V93 1.3487398655197228e-19

R27_94 V27 V94 11291.98854943411
L27_94 V27 V94 -1.8000984706394215e-11
C27_94 V27 V94 -1.194083324357558e-19

R27_95 V27 V95 3673.7152716421074
L27_95 V27 V95 -5.8962622676400024e-12
C27_95 V27 V95 -2.9675031449600175e-19

R27_96 V27 V96 2688.602166288301
L27_96 V27 V96 5.53390230025042e-12
C27_96 V27 V96 -2.5955727765430864e-20

R27_97 V27 V97 -21894.55997257079
L27_97 V27 V97 -2.0912223214598933e-12
C27_97 V27 V97 -5.082713830713791e-19

R27_98 V27 V98 -6302.517898865719
L27_98 V27 V98 -1.1284805318702513e-12
C27_98 V27 V98 -5.413476630519401e-19

R27_99 V27 V99 1093.5189720935875
L27_99 V27 V99 5.309133879993702e-13
C27_99 V27 V99 1.1073235256414073e-18

R27_100 V27 V100 -7362.013708611622
L27_100 V27 V100 2.84083455091468e-12
C27_100 V27 V100 3.091544142727231e-19

R27_101 V27 V101 11725.446876967373
L27_101 V27 V101 6.204943483517078e-12
C27_101 V27 V101 1.9614616181708444e-19

R27_102 V27 V102 77192.06309250041
L27_102 V27 V102 3.309223336830052e-12
C27_102 V27 V102 2.7105488332019847e-19

R27_103 V27 V103 -1284.4847817894017
L27_103 V27 V103 -2.3332729281197927e-12
C27_103 V27 V103 -1.273520111915968e-19

R27_104 V27 V104 -5021.444482159814
L27_104 V27 V104 -2.4797927491448744e-12
C27_104 V27 V104 -2.3605685776834103e-19

R27_105 V27 V105 -3145.238496097137
L27_105 V27 V105 -3.332804397606246e-11
C27_105 V27 V105 1.5047006531908857e-19

R27_106 V27 V106 12146.867896059277
L27_106 V27 V106 1.1486500958075809e-12
C27_106 V27 V106 4.687012534595118e-19

R27_107 V27 V107 -3753.1375125480913
L27_107 V27 V107 -9.069808656421918e-13
C27_107 V27 V107 -7.384675130949944e-19

R27_108 V27 V108 5495.718541320431
L27_108 V27 V108 1.0896931347618802e-11
C27_108 V27 V108 6.207649392726946e-20

R27_109 V27 V109 -24021.975590374357
L27_109 V27 V109 -2.0939982443141943e-12
C27_109 V27 V109 -3.9372733612509256e-19

R27_110 V27 V110 5139.502173745949
L27_110 V27 V110 -1.782890831726726e-12
C27_110 V27 V110 -3.5793694446911845e-19

R27_111 V27 V111 1956.7480607739537
L27_111 V27 V111 -4.345872311510999e-12
C27_111 V27 V111 -1.7126062428070666e-19

R27_112 V27 V112 -17787.964698842192
L27_112 V27 V112 5.56806917227754e-12
C27_112 V27 V112 6.180637871911855e-20

R27_113 V27 V113 -8486.483745487134
L27_113 V27 V113 7.473374820393021e-12
C27_113 V27 V113 4.869671635134579e-20

R27_114 V27 V114 -10715.451885992252
L27_114 V27 V114 -1.5543810767259926e-12
C27_114 V27 V114 -3.8999759518859318e-19

R27_115 V27 V115 2968.145371064409
L27_115 V27 V115 7.19080488069995e-13
C27_115 V27 V115 7.820813668398725e-19

R27_116 V27 V116 8425.724596199248
L27_116 V27 V116 -1.156027753599041e-11
C27_116 V27 V116 -9.582251116585604e-20

R27_117 V27 V117 2280.3604144893943
L27_117 V27 V117 2.0347414756845714e-12
C27_117 V27 V117 2.3025516422341244e-19

R27_118 V27 V118 -8785.932347114172
L27_118 V27 V118 1.319416187466181e-12
C27_118 V27 V118 4.794876619015012e-19

R27_119 V27 V119 -1138.2742130196482
L27_119 V27 V119 -2.8988679129755937e-11
C27_119 V27 V119 4.5883689984962704e-20

R27_120 V27 V120 -3244.741019718547
L27_120 V27 V120 9.725742902838992e-12
C27_120 V27 V120 2.3778354758551327e-19

R27_121 V27 V121 -2372.188034328256
L27_121 V27 V121 -2.1494958456163956e-12
C27_121 V27 V121 -1.8933887645269484e-19

R27_122 V27 V122 22744.23845422009
L27_122 V27 V122 -1.8349226330885957e-11
C27_122 V27 V122 -8.529620928615237e-21

R27_123 V27 V123 3367.2482033765223
L27_123 V27 V123 -6.934219007812649e-13
C27_123 V27 V123 -9.430860165450368e-19

R27_124 V27 V124 13482.309490688438
L27_124 V27 V124 -2.0772972995668272e-11
C27_124 V27 V124 -2.0747929698385763e-19

R27_125 V27 V125 -1319.585208764804
L27_125 V27 V125 -3.3323732774630843e-12
C27_125 V27 V125 -4.9073559396303344e-21

R27_126 V27 V126 56273.00024211312
L27_126 V27 V126 -1.3649354309695995e-12
C27_126 V27 V126 -3.5367844766380175e-19

R27_127 V27 V127 1713.0362126749262
L27_127 V27 V127 4.4350100569964e-12
C27_127 V27 V127 3.7179696412621983e-19

R27_128 V27 V128 2364.884459234133
L27_128 V27 V128 -3.348657358597207e-12
C27_128 V27 V128 -1.4963453043580936e-19

R27_129 V27 V129 1065.5684771533067
L27_129 V27 V129 -2.7514876439906005e-11
C27_129 V27 V129 -2.0466839572420239e-19

R27_130 V27 V130 4289.826902639361
L27_130 V27 V130 1.89862302720893e-12
C27_130 V27 V130 2.462913938956117e-19

R27_131 V27 V131 -2331.0409455111626
L27_131 V27 V131 1.2697062491528702e-12
C27_131 V27 V131 3.764678548350541e-19

R27_132 V27 V132 -1872.4296440036583
L27_132 V27 V132 1.6520235033994692e-12
C27_132 V27 V132 4.621838951304788e-19

R27_133 V27 V133 4495.719496010614
L27_133 V27 V133 2.839193626072999e-12
C27_133 V27 V133 2.477318332773392e-19

R27_134 V27 V134 -2429.094243491309
L27_134 V27 V134 7.200721204132415e-12
C27_134 V27 V134 4.892591639976562e-20

R27_135 V27 V135 -160596.51640270997
L27_135 V27 V135 -1.7694382202555937e-12
C27_135 V27 V135 -8.520002118455362e-19

R27_136 V27 V136 -3736.629537395886
L27_136 V27 V136 2.86724712655963e-12
C27_136 V27 V136 -1.3323048912271093e-19

R27_137 V27 V137 -985.7653103424351
L27_137 V27 V137 1.9274106343387065e-12
C27_137 V27 V137 1.4774589153424077e-19

R27_138 V27 V138 5842.119221884008
L27_138 V27 V138 -1.9147070431450605e-12
C27_138 V27 V138 -2.3275706700433394e-19

R27_139 V27 V139 -5263.166887842906
L27_139 V27 V139 1.586335351816964e-12
C27_139 V27 V139 9.832830344066146e-19

R27_140 V27 V140 4271.2085850952535
L27_140 V27 V140 -1.382458502434762e-12
C27_140 V27 V140 8.273259930044713e-20

R27_141 V27 V141 -12304.55008187582
L27_141 V27 V141 -1.088119877156394e-12
C27_141 V27 V141 -4.77984277990666e-19

R27_142 V27 V142 1202.9256185832032
L27_142 V27 V142 -6.503994708145039e-12
C27_142 V27 V142 9.460767109094126e-21

R27_143 V27 V143 5994.959001289301
L27_143 V27 V143 -1.5382797712741855e-12
C27_143 V27 V143 -1.8937198921562617e-19

R27_144 V27 V144 1978.8969079129906
L27_144 V27 V144 1.7294602103648112e-11
C27_144 V27 V144 -2.186549357720683e-20

R27_145 V27 V145 971.4891167027233
L27_145 V27 V145 -1.3233819256794617e-12
C27_145 V27 V145 -1.694809491805151e-19

R27_146 V27 V146 -3617.414015660754
L27_146 V27 V146 1.6096687035835451e-12
C27_146 V27 V146 1.9674793216602965e-19

R27_147 V27 V147 802.4400691708545
L27_147 V27 V147 6.286747577655808e-12
C27_147 V27 V147 -6.725779949438032e-19

R27_148 V27 V148 -1724.2094949119676
L27_148 V27 V148 7.133149367791158e-11
C27_148 V27 V148 -1.5091612987330804e-19

R27_149 V27 V149 14607.605961241337
L27_149 V27 V149 5.973092946781183e-13
C27_149 V27 V149 6.338681846509524e-19

R27_150 V27 V150 -853.4800806861932
L27_150 V27 V150 -8.889054345030268e-12
C27_150 V27 V150 -2.6824895811679963e-19

R27_151 V27 V151 -554.4475708796497
L27_151 V27 V151 4.052215131778299e-12
C27_151 V27 V151 2.2999880977050037e-19

R27_152 V27 V152 5797.24317022459
L27_152 V27 V152 -4.927982264605744e-12
C27_152 V27 V152 -3.920941798512831e-21

R27_153 V27 V153 -930.1497756059966
L27_153 V27 V153 3.6221703746499e-12
C27_153 V27 V153 1.1061990043649627e-20

R27_154 V27 V154 -10580.593839786372
L27_154 V27 V154 -3.4438678130651206e-12
C27_154 V27 V154 4.387513790332256e-20

R27_155 V27 V155 611.1185060133122
L27_155 V27 V155 2.0529503033397383e-12
C27_155 V27 V155 5.190366014797927e-19

R27_156 V27 V156 -1692.5297821621687
L27_156 V27 V156 -2.4652087078457105e-09
C27_156 V27 V156 1.0427721154932532e-19

R27_157 V27 V157 -1768.7969008254008
L27_157 V27 V157 -7.321616724687351e-13
C27_157 V27 V157 -4.38399131161822e-19

R27_158 V27 V158 1716.750253865053
L27_158 V27 V158 3.607607965591413e-12
C27_158 V27 V158 9.250785387740875e-20

R27_159 V27 V159 -9629.701021215227
L27_159 V27 V159 -1.070126028562601e-12
C27_159 V27 V159 -3.8791045446940204e-19

R27_160 V27 V160 2008.1663299658596
L27_160 V27 V160 1.6372306609320788e-12
C27_160 V27 V160 7.788492637374077e-20

R27_161 V27 V161 1631.0233036225893
L27_161 V27 V161 -5.879242029873811e-11
C27_161 V27 V161 1.7385005963274176e-20

R27_162 V27 V162 8661.278832577167
L27_162 V27 V162 1.4397652892132473e-12
C27_162 V27 V162 1.9647140015602596e-19

R27_163 V27 V163 2142.426661404224
L27_163 V27 V163 9.180556087209043e-13
C27_163 V27 V163 2.7136279107758253e-19

R27_164 V27 V164 -1816.9594851941508
L27_164 V27 V164 -7.264103436231029e-12
C27_164 V27 V164 5.948619933616111e-20

R27_165 V27 V165 -5791.873165047811
L27_165 V27 V165 4.6349781393237194e-12
C27_165 V27 V165 -1.593912999560603e-20

R27_166 V27 V166 -1301.8297604806835
L27_166 V27 V166 -1.901666756370337e-12
C27_166 V27 V166 -2.1178813864918266e-19

R27_167 V27 V167 -540.1147502385815
L27_167 V27 V167 -3.1357137573240905e-12
C27_167 V27 V167 -9.309730488048378e-20

R27_168 V27 V168 869.2412823684693
L27_168 V27 V168 -6.6472234096624534e-12
C27_168 V27 V168 -5.676108223720938e-20

R27_169 V27 V169 -1912.2167208149378
L27_169 V27 V169 -1.8055314018773434e-10
C27_169 V27 V169 -1.4869576234152046e-19

R27_170 V27 V170 2268.1000822321125
L27_170 V27 V170 2.97094294239726e-10
C27_170 V27 V170 1.1441194150332223e-19

R27_171 V27 V171 851.9939736498736
L27_171 V27 V171 -1.4269393442237015e-12
C27_171 V27 V171 -8.926207905440136e-20

R27_172 V27 V172 -30214.89740285318
L27_172 V27 V172 1.5792322069133127e-10
C27_172 V27 V172 -2.2258477795617122e-22

R27_173 V27 V173 4231.887860328603
L27_173 V27 V173 5.936462774399615e-12
C27_173 V27 V173 2.5548690463924387e-19

R27_174 V27 V174 1793.2873224150312
L27_174 V27 V174 1.4867667265849181e-12
C27_174 V27 V174 -3.9960502416595317e-20

R27_175 V27 V175 1829.95647703448
L27_175 V27 V175 6.802063266528993e-13
C27_175 V27 V175 4.99126145968221e-19

R27_176 V27 V176 -2863.4001091352493
L27_176 V27 V176 1.851194127248531e-12
C27_176 V27 V176 1.7281381531087523e-19

R27_177 V27 V177 -3551.8173513281045
L27_177 V27 V177 -3.692607243850818e-12
C27_177 V27 V177 -1.2095209938187474e-19

R27_178 V27 V178 -1446.3909022149137
L27_178 V27 V178 -2.1503018390345223e-12
C27_178 V27 V178 -5.911828340751141e-20

R27_179 V27 V179 -2938.1370139593228
L27_179 V27 V179 -3.82132465433284e-12
C27_179 V27 V179 -4.285136575466774e-19

R27_180 V27 V180 -7702.827727874866
L27_180 V27 V180 -1.8630862116753148e-12
C27_180 V27 V180 -1.900046265692621e-19

R27_181 V27 V181 3543.074106887827
L27_181 V27 V181 6.0819081067768036e-12
C27_181 V27 V181 -1.7934759042460356e-19

R27_182 V27 V182 2581.4326375470073
L27_182 V27 V182 3.748788966245535e-12
C27_182 V27 V182 1.0869176615063946e-19

R27_183 V27 V183 -1553.4853694589851
L27_183 V27 V183 -9.33739158941863e-13
C27_183 V27 V183 2.3704411506433336e-22

R27_184 V27 V184 -7918.2770961268425
L27_184 V27 V184 -2.215933532936876e-12
C27_184 V27 V184 -6.325589915683089e-20

R27_185 V27 V185 -3730.373535497999
L27_185 V27 V185 -3.497622494968399e-12
C27_185 V27 V185 1.806529136566953e-19

R27_186 V27 V186 9182.094980913103
L27_186 V27 V186 -2.9662095579624716e-12
C27_186 V27 V186 -2.1012120291340907e-19

R27_187 V27 V187 1440.319289768826
L27_187 V27 V187 8.969503242760966e-13
C27_187 V27 V187 4.595101793475983e-19

R27_188 V27 V188 1386.2701308324422
L27_188 V27 V188 1.8672716827949597e-12
C27_188 V27 V188 1.7236975117158833e-19

R27_189 V27 V189 -13774.384760393781
L27_189 V27 V189 4.528262971019361e-12
C27_189 V27 V189 9.646717583811498e-21

R27_190 V27 V190 -2989.073215833528
L27_190 V27 V190 1.6446664756884664e-11
C27_190 V27 V190 -4.8258096340193454e-20

R27_191 V27 V191 14441.295750208043
L27_191 V27 V191 2.750032762498808e-12
C27_191 V27 V191 -3.273127570233011e-19

R27_192 V27 V192 -4934.032813387569
L27_192 V27 V192 2.3801185989352475e-12
C27_192 V27 V192 1.4999387081016529e-21

R27_193 V27 V193 2528.9647933750703
L27_193 V27 V193 2.7287593766758524e-12
C27_193 V27 V193 -1.2948963106159296e-20

R27_194 V27 V194 -28863.432379997463
L27_194 V27 V194 7.019885092379152e-12
C27_194 V27 V194 -1.284925593581552e-19

R27_195 V27 V195 -2300.85744194905
L27_195 V27 V195 -1.681712727595847e-12
C27_195 V27 V195 2.9726315650134626e-19

R27_196 V27 V196 -1320.5720689017726
L27_196 V27 V196 -1.4357448961854759e-12
C27_196 V27 V196 -2.0547262285109717e-19

R27_197 V27 V197 -7532.4513630843585
L27_197 V27 V197 -2.030295316775961e-12
C27_197 V27 V197 -8.998043259841168e-20

R27_198 V27 V198 -12187.196097206644
L27_198 V27 V198 -1.452999210264512e-10
C27_198 V27 V198 6.0872811913516224e-21

R27_199 V27 V199 -14689.582593022848
L27_199 V27 V199 2.4379959098948356e-11
C27_199 V27 V199 5.47419313148079e-20

R27_200 V27 V200 1355.5195370009485
L27_200 V27 V200 -1.5886903269459592e-11
C27_200 V27 V200 1.3875930320856448e-19

R28_28 V28 0 201.7893807364711
L28_28 V28 0 1.1245152341083728e-13
C28_28 V28 0 3.947621448535314e-18

R28_29 V28 V29 -2268.2378760332444
L28_29 V28 V29 -1.6560242682772769e-12
C28_29 V28 V29 -1.0667249880173017e-20

R28_30 V28 V30 -5338.061406047357
L28_30 V28 V30 3.316895651848304e-11
C28_30 V28 V30 1.6315049476832207e-19

R28_31 V28 V31 -2906.9713368211656
L28_31 V28 V31 5.732698654219096e-11
C28_31 V28 V31 1.7099978638637392e-19

R28_32 V28 V32 -2104.1150428514798
L28_32 V28 V32 1.3288592802718452e-11
C28_32 V28 V32 6.245906960446697e-19

R28_33 V28 V33 -17374.75656288837
L28_33 V28 V33 2.6069199616037077e-12
C28_33 V28 V33 1.9069046247655958e-19

R28_34 V28 V34 6470.742737301738
L28_34 V28 V34 1.6636397762873108e-12
C28_34 V28 V34 2.92978752771067e-19

R28_35 V28 V35 4704.84748990494
L28_35 V28 V35 1.2951871390540161e-12
C28_35 V28 V35 3.483280827500159e-19

R28_36 V28 V36 1572.9969683607267
L28_36 V28 V36 4.374601583212102e-13
C28_36 V28 V36 1.3316520929010494e-18

R28_37 V28 V37 3546.8334655149833
L28_37 V28 V37 1.2463167946151712e-12
C28_37 V28 V37 2.38259333622496e-19

R28_38 V28 V38 6400.545016659394
L28_38 V28 V38 3.8802409509447766e-12
C28_38 V28 V38 3.253390427090994e-20

R28_39 V28 V39 3806.134693654282
L28_39 V28 V39 -7.990130876134945e-12
C28_39 V28 V39 -2.4017159588990744e-19

R28_40 V28 V40 2417.6101879447606
L28_40 V28 V40 -1.6373400555142743e-12
C28_40 V28 V40 -7.541412335176771e-19

R28_41 V28 V41 -12515.593099042691
L28_41 V28 V41 -2.7469656505902807e-10
C28_41 V28 V41 -9.989650307205041e-20

R28_42 V28 V42 -41420.221877622724
L28_42 V28 V42 -1.6357568361267143e-11
C28_42 V28 V42 -8.297880995477365e-20

R28_43 V28 V43 26444.558158037453
L28_43 V28 V43 2.901194368086836e-12
C28_43 V28 V43 1.5017704120356954e-19

R28_44 V28 V44 4387.692200053524
L28_44 V28 V44 2.685706123109823e-12
C28_44 V28 V44 2.0234316877686894e-19

R28_45 V28 V45 -2672.292804772082
L28_45 V28 V45 -8.833442047219349e-13
C28_45 V28 V45 -4.683945178719232e-19

R28_46 V28 V46 -3562.5628823819216
L28_46 V28 V46 -1.3822132760273303e-12
C28_46 V28 V46 -3.7870176065937577e-19

R28_47 V28 V47 -3586.922136153953
L28_47 V28 V47 -1.7818567510503465e-12
C28_47 V28 V47 -2.6989471195511427e-19

R28_48 V28 V48 -1907.4551957986143
L28_48 V28 V48 -7.340230416532414e-13
C28_48 V28 V48 -5.346589825962177e-19

R28_49 V28 V49 -6417.2102066143825
L28_49 V28 V49 -1.753730286053898e-11
C28_49 V28 V49 -6.304216026604932e-20

R28_50 V28 V50 -42381.398875583014
L28_50 V28 V50 -1.0078732966046532e-10
C28_50 V28 V50 -7.925732747810446e-20

R28_51 V28 V51 -6739.934136718356
L28_51 V28 V51 -5.39505166632664e-12
C28_51 V28 V51 -7.680702474972247e-20

R28_52 V28 V52 -64383.547537193605
L28_52 V28 V52 4.869780624684412e-12
C28_52 V28 V52 1.8396208228366883e-19

R28_53 V28 V53 -11659.41065900817
L28_53 V28 V53 3.710078286483297e-12
C28_53 V28 V53 3.607757587014803e-19

R28_54 V28 V54 6704.848943166559
L28_54 V28 V54 1.4517330232116673e-12
C28_54 V28 V54 4.562731000688458e-19

R28_55 V28 V55 14787.061271323379
L28_55 V28 V55 2.701657601799203e-12
C28_55 V28 V55 2.728642785658471e-19

R28_56 V28 V56 3597.933339176742
L28_56 V28 V56 7.699041053437559e-13
C28_56 V28 V56 9.127189348496728e-19

R28_57 V28 V57 30263.788778725
L28_57 V28 V57 2.3659582953089456e-12
C28_57 V28 V57 -1.6187795217697532e-20

R28_58 V28 V58 -7616.08726365919
L28_58 V28 V58 -7.147048841722706e-12
C28_58 V28 V58 -1.2328978422868962e-19

R28_59 V28 V59 9024.689800119379
L28_59 V28 V59 -4.5782739386795445e-12
C28_59 V28 V59 -3.2506302062756666e-19

R28_60 V28 V60 2133.0352529089155
L28_60 V28 V60 -8.356055725118656e-12
C28_60 V28 V60 -4.482192410897571e-19

R28_61 V28 V61 -34178.14145848689
L28_61 V28 V61 -1.8546968776352027e-12
C28_61 V28 V61 -2.7304912309438593e-19

R28_62 V28 V62 18253.353796568288
L28_62 V28 V62 -2.1668765936785575e-12
C28_62 V28 V62 -3.842505419979138e-19

R28_63 V28 V63 -70342.13780602386
L28_63 V28 V63 4.41789958979881e-12
C28_63 V28 V63 9.433869392961708e-20

R28_64 V28 V64 -4387.955342948492
L28_64 V28 V64 -2.2533565393502173e-12
C28_64 V28 V64 -9.535183373621903e-20

R28_65 V28 V65 -4577.551604326964
L28_65 V28 V65 -3.0978832438450306e-12
C28_65 V28 V65 -2.0846631840300861e-19

R28_66 V28 V66 -10485.801240687571
L28_66 V28 V66 2.6193132561214397e-11
C28_66 V28 V66 -1.6489354551667778e-21

R28_67 V28 V67 -54617.70472522356
L28_67 V28 V67 3.5082966754786767e-12
C28_67 V28 V67 1.8603693778849413e-19

R28_68 V28 V68 -4959.04992060532
L28_68 V28 V68 -1.3279746526341664e-11
C28_68 V28 V68 1.1412871886247664e-19

R28_69 V28 V69 -17600.60039347679
L28_69 V28 V69 9.125861381079864e-12
C28_69 V28 V69 2.410205583100751e-19

R28_70 V28 V70 14192.769565364773
L28_70 V28 V70 2.6337329473558715e-12
C28_70 V28 V70 2.9173390823591965e-19

R28_71 V28 V71 -7553.497604270004
L28_71 V28 V71 -1.5418656454605066e-12
C28_71 V28 V71 -2.457179508632987e-19

R28_72 V28 V72 -11276.51195286924
L28_72 V28 V72 -1.2824766434943615e-12
C28_72 V28 V72 -3.750295835158511e-19

R28_73 V28 V73 -10883.581559742854
L28_73 V28 V73 -4.921062396160519e-12
C28_73 V28 V73 -8.026517021101419e-20

R28_74 V28 V74 9576.868371216813
L28_74 V28 V74 -7.79951753929763e-12
C28_74 V28 V74 -1.524832414092709e-19

R28_75 V28 V75 119941.1118473167
L28_75 V28 V75 -2.6719465957910925e-11
C28_75 V28 V75 -1.5143353967303446e-19

R28_76 V28 V76 2343.667329071293
L28_76 V28 V76 6.57438289367569e-13
C28_76 V28 V76 7.621719887961287e-19

R28_77 V28 V77 6706.191871586513
L28_77 V28 V77 2.0283789104906265e-12
C28_77 V28 V77 4.6902939481193207e-20

R28_78 V28 V78 -5297.896006945133
L28_78 V28 V78 5.9713865558326546e-12
C28_78 V28 V78 2.1665617585970513e-19

R28_79 V28 V79 7016.540915462009
L28_79 V28 V79 2.39647767664239e-12
C28_79 V28 V79 2.191528554444578e-19

R28_80 V28 V80 -11680.650334932898
L28_80 V28 V80 -3.896525991863718e-12
C28_80 V28 V80 -1.9599853445211637e-19

R28_81 V28 V81 -1873.0934293675236
L28_81 V28 V81 -1.3883882528477382e-12
C28_81 V28 V81 -3.1989692701921012e-19

R28_82 V28 V82 9325.747944855168
L28_82 V28 V82 -2.686492066064308e-12
C28_82 V28 V82 -3.4408699521229363e-19

R28_83 V28 V83 22063.278791098342
L28_83 V28 V83 1.455475902275198e-11
C28_83 V28 V83 -2.872718871808673e-20

R28_84 V28 V84 -60613.556276100535
L28_84 V28 V84 -9.977134127259776e-13
C28_84 V28 V84 -5.429017661062476e-19

R28_85 V28 V85 42678.86254023547
L28_85 V28 V85 -2.0120897493200608e-12
C28_85 V28 V85 -2.483331302569521e-19

R28_86 V28 V86 -9775.026214492704
L28_86 V28 V86 -1.614121901101976e-12
C28_86 V28 V86 -3.5315660361995973e-19

R28_87 V28 V87 -20988.231829312073
L28_87 V28 V87 8.11106977718703e-12
C28_87 V28 V87 7.005354066463788e-20

R28_88 V28 V88 2857.3955629943675
L28_88 V28 V88 7.346721735932204e-13
C28_88 V28 V88 7.925331628480643e-19

R28_89 V28 V89 8207.777128920878
L28_89 V28 V89 1.6718672467942236e-12
C28_89 V28 V89 4.260719039317359e-19

R28_90 V28 V90 11645.803808823684
L28_90 V28 V90 6.513185067481458e-13
C28_90 V28 V90 8.886367076038016e-19

R28_91 V28 V91 -2772.759331289884
L28_91 V28 V91 -9.87499565170968e-13
C28_91 V28 V91 -4.134899245693492e-19

R28_92 V28 V92 -1163.17062296449
L28_92 V28 V92 -6.113718139272535e-13
C28_92 V28 V92 -6.267009417577722e-19

R28_93 V28 V93 -3056.1808427453834
L28_93 V28 V93 3.343844856095135e-12
C28_93 V28 V93 1.3885317663010156e-19

R28_94 V28 V94 7735.396950464123
L28_94 V28 V94 -7.44879085409488e-12
C28_94 V28 V94 -2.0858035435429715e-19

R28_95 V28 V95 3261.138383508122
L28_95 V28 V95 5.8252521903991595e-12
C28_95 V28 V95 -1.3335960931539743e-20

R28_96 V28 V96 2757.585966004047
L28_96 V28 V96 -1.3746250577095504e-11
C28_96 V28 V96 -3.8458321889319676e-19

R28_97 V28 V97 -7927.173177135954
L28_97 V28 V97 -1.206361244876356e-12
C28_97 V28 V97 -6.875040290637218e-19

R28_98 V28 V98 -5384.024868828803
L28_98 V28 V98 -7.528166355657752e-13
C28_98 V28 V98 -7.010730750721891e-19

R28_99 V28 V99 3607.3520091105365
L28_99 V28 V99 7.984775704429021e-13
C28_99 V28 V99 5.202118481014673e-19

R28_100 V28 V100 1069.5050983954516
L28_100 V28 V100 5.844324381388174e-13
C28_100 V28 V100 1.0715130597712474e-18

R28_101 V28 V101 7605.539471665387
L28_101 V28 V101 4.95610264871332e-12
C28_101 V28 V101 1.7769155212046989e-19

R28_102 V28 V102 162025.2670731539
L28_102 V28 V102 1.8019903236906984e-12
C28_102 V28 V102 4.2402783487944945e-19

R28_103 V28 V103 -3116.593914279861
L28_103 V28 V103 -2.0145066067029047e-12
C28_103 V28 V103 -1.4333989101368258e-19

R28_104 V28 V104 -1270.9661306657165
L28_104 V28 V104 -1.3761431253401502e-12
C28_104 V28 V104 -2.4026305637662333e-19

R28_105 V28 V105 -2183.800469093797
L28_105 V28 V105 1.2800471983529113e-11
C28_105 V28 V105 2.095201477144118e-19

R28_106 V28 V106 5506.189101864126
L28_106 V28 V106 9.090674029126202e-13
C28_106 V28 V106 4.625687561128388e-19

R28_107 V28 V107 -17543.041165110415
L28_107 V28 V107 -1.437482859778296e-12
C28_107 V28 V107 -4.052156220066687e-19

R28_108 V28 V108 -5828.317514982216
L28_108 V28 V108 -2.6895301732676393e-12
C28_108 V28 V108 -3.5506703586075824e-19

R28_109 V28 V109 -7024.930562826704
L28_109 V28 V109 -1.3769234055569261e-12
C28_109 V28 V109 -5.219407479503599e-19

R28_110 V28 V110 7057.487397575923
L28_110 V28 V110 -1.5328580102175507e-12
C28_110 V28 V110 -3.3384535629884397e-19

R28_111 V28 V111 12365.226514882044
L28_111 V28 V111 6.631214714702839e-12
C28_111 V28 V111 1.0149327103828242e-19

R28_112 V28 V112 2460.7806366757018
L28_112 V28 V112 -1.3944410111038908e-12
C28_112 V28 V112 -5.332809611943278e-19

R28_113 V28 V113 -9390.956405652858
L28_113 V28 V113 9.758378467046344e-12
C28_113 V28 V113 5.778358765411795e-20

R28_114 V28 V114 -10213.153972789356
L28_114 V28 V114 -1.1216358626170665e-12
C28_114 V28 V114 -4.161751028154095e-19

R28_115 V28 V115 3036.2985066672563
L28_115 V28 V115 1.788904700401914e-12
C28_115 V28 V115 2.465896388406002e-19

R28_116 V28 V116 2519.3837575029947
L28_116 V28 V116 7.472860007695417e-13
C28_116 V28 V116 6.89187974512501e-19

R28_117 V28 V117 1758.8995427455957
L28_117 V28 V117 1.234822922916134e-12
C28_117 V28 V117 3.5247538337353475e-19

R28_118 V28 V118 -26598.187481532947
L28_118 V28 V118 9.766679200551003e-13
C28_118 V28 V118 5.365130009024223e-19

R28_119 V28 V119 -3335.5668335808878
L28_119 V28 V119 8.134671217812658e-12
C28_119 V28 V119 1.9955536914474034e-19

R28_120 V28 V120 -1017.7643672526344
L28_120 V28 V120 2.289739577982698e-12
C28_120 V28 V120 5.715119680267843e-19

R28_121 V28 V121 -1549.1563578131725
L28_121 V28 V121 -1.4880706196109047e-12
C28_121 V28 V121 -3.0288851867148013e-19

R28_122 V28 V122 -28508.35629098413
L28_122 V28 V122 -2.169186031029884e-11
C28_122 V28 V122 6.80042356226757e-21

R28_123 V28 V123 -18254.74011115568
L28_123 V28 V123 -2.912358248048618e-12
C28_123 V28 V123 -1.8723218265290867e-19

R28_124 V28 V124 3318.8839399830445
L28_124 V28 V124 -4.3941873416316466e-13
C28_124 V28 V124 -1.6386184514381055e-18

R28_125 V28 V125 -951.2614054824556
L28_125 V28 V125 -1.7181055710034721e-12
C28_125 V28 V125 -7.86010746109519e-20

R28_126 V28 V126 -19193.151131181985
L28_126 V28 V126 -9.139572716013971e-13
C28_126 V28 V126 -3.9503828497944384e-19

R28_127 V28 V127 3413.371759928065
L28_127 V28 V127 -2.017986214417961e-12
C28_127 V28 V127 -3.2163860095678245e-19

R28_128 V28 V128 1368.2900348473772
L28_128 V28 V128 4.4682767852733915e-12
C28_128 V28 V128 2.894355958799748e-19

R28_129 V28 V129 833.8911236537011
L28_129 V28 V129 -2.0116764421420796e-11
C28_129 V28 V129 -2.65764326328694e-19

R28_130 V28 V130 2661.155618759165
L28_130 V28 V130 1.1686668843916392e-12
C28_130 V28 V130 3.8283278578786374e-19

R28_131 V28 V131 -3070.8756162036407
L28_131 V28 V131 1.836287715523021e-12
C28_131 V28 V131 4.085188752914362e-19

R28_132 V28 V132 -1560.1646284603742
L28_132 V28 V132 6.750064729835286e-13
C28_132 V28 V132 8.656261984822855e-19

R28_133 V28 V133 2464.7044281757167
L28_133 V28 V133 1.246749285629554e-12
C28_133 V28 V133 5.335982879788735e-19

R28_134 V28 V134 -2148.15663685284
L28_134 V28 V134 3.1873557405553457e-12
C28_134 V28 V134 1.5984254149417725e-19

R28_135 V28 V135 -58666.615143387295
L28_135 V28 V135 2.0187690084325426e-12
C28_135 V28 V135 1.478403015752655e-19

R28_136 V28 V136 -4381.839197568745
L28_136 V28 V136 -1.4523217521268227e-12
C28_136 V28 V136 -1.0908804270438143e-18

R28_137 V28 V137 -763.0339667495525
L28_137 V28 V137 1.895131533673409e-12
C28_137 V28 V137 1.2878052431070366e-19

R28_138 V28 V138 8883.224639126478
L28_138 V28 V138 -1.1463625249372391e-12
C28_138 V28 V138 -3.316362966565589e-19

R28_139 V28 V139 4309.9955542805865
L28_139 V28 V139 -1.5019419287487022e-12
C28_139 V28 V139 -1.684285675867074e-19

R28_140 V28 V140 -3903.4523930321775
L28_140 V28 V140 1.2255955502421776e-11
C28_140 V28 V140 1.0737163974465743e-18

R28_141 V28 V141 -8892.381832658837
L28_141 V28 V141 -6.938654572937932e-13
C28_141 V28 V141 -7.628040668048979e-19

R28_142 V28 V142 960.5407691749792
L28_142 V28 V142 -6.363198347301364e-12
C28_142 V28 V142 3.460283926444792e-21

R28_143 V28 V143 29841.35557036406
L28_143 V28 V143 -5.955378244580702e-12
C28_143 V28 V143 -7.020131932617869e-20

R28_144 V28 V144 821.0346465869673
L28_144 V28 V144 -5.906752488586967e-12
C28_144 V28 V144 -2.082233766031874e-19

R28_145 V28 V145 903.5633845921918
L28_145 V28 V145 -1.1195616621895541e-12
C28_145 V28 V145 -1.6581333635991447e-19

R28_146 V28 V146 -5981.842665381214
L28_146 V28 V146 1.0232130164626961e-12
C28_146 V28 V146 2.5135350379967113e-19

R28_147 V28 V147 1298.226654466236
L28_147 V28 V147 2.3630180350561135e-11
C28_147 V28 V147 -2.390768088356881e-19

R28_148 V28 V148 -1063.9358200726147
L28_148 V28 V148 -1.210416223254575e-12
C28_148 V28 V148 -7.008181515270383e-19

R28_149 V28 V149 2273.8187509458608
L28_149 V28 V149 4.3930493948503014e-13
C28_149 V28 V149 7.534580536044497e-19

R28_150 V28 V150 -675.6980306228576
L28_150 V28 V150 -2.4733155339573765e-12
C28_150 V28 V150 -5.363349803868429e-19

R28_151 V28 V151 -801.2066098132218
L28_151 V28 V151 -5.82697459845107e-12
C28_151 V28 V151 6.939579869175345e-20

R28_152 V28 V152 5759.979920975385
L28_152 V28 V152 8.957341239213205e-13
C28_152 V28 V152 1.872110492311103e-19

R28_153 V28 V153 -680.2708011874175
L28_153 V28 V153 1.4701858663342292e-12
C28_153 V28 V153 2.365349366150123e-19

R28_154 V28 V154 -11136.106750140843
L28_154 V28 V154 -1.5349325682683955e-11
C28_154 V28 V154 1.9302352592733103e-19

R28_155 V28 V155 566.518720423171
L28_155 V28 V155 1.6702807589096555e-12
C28_155 V28 V155 1.747408789997705e-19

R28_156 V28 V156 -546.6206447558704
L28_156 V28 V156 -1.1016589006578703e-12
C28_156 V28 V156 5.99228516893025e-19

R28_157 V28 V157 -1008.0234883988041
L28_157 V28 V157 -4.2267949986171593e-13
C28_157 V28 V157 -8.232131282090545e-19

R28_158 V28 V158 1447.759582634378
L28_158 V28 V158 5.1371599203710454e-12
C28_158 V28 V158 7.120112749028328e-20

R28_159 V28 V159 -962.9698548960961
L28_159 V28 V159 3.3560544194113135e-12
C28_159 V28 V159 8.147044555234516e-20

R28_160 V28 V160 536.9906579610273
L28_160 V28 V160 -2.083865851721046e-11
C28_160 V28 V160 -2.1222274958684472e-19

R28_161 V28 V161 1494.1055492135026
L28_161 V28 V161 1.257812201974842e-11
C28_161 V28 V161 -6.862209400760985e-20

R28_162 V28 V162 7470.036336914956
L28_162 V28 V162 1.1384638609827825e-12
C28_162 V28 V162 2.087529037447225e-19

R28_163 V28 V163 -32337.792717275093
L28_163 V28 V163 -3.127206368014327e-11
C28_163 V28 V163 -7.626298481825239e-20

R28_164 V28 V164 -3268.926889313238
L28_164 V28 V164 1.65760996211672e-12
C28_164 V28 V164 2.415623517289327e-19

R28_165 V28 V165 -3417.423764124518
L28_165 V28 V165 6.216277623398334e-12
C28_165 V28 V165 6.691908741325378e-20

R28_166 V28 V166 -966.474419440193
L28_166 V28 V166 -1.1393766821298845e-12
C28_166 V28 V166 -3.7059806689989727e-19

R28_167 V28 V167 -5726.338475730675
L28_167 V28 V167 -2.3329822295673364e-12
C28_167 V28 V167 -4.69156553436768e-20

R28_168 V28 V168 -2653.8393384661335
L28_168 V28 V168 -6.184892883051538e-11
C28_168 V28 V168 -2.316118475122985e-19

R28_169 V28 V169 -1543.9729111567103
L28_169 V28 V169 2.1983655951442655e-11
C28_169 V28 V169 -1.7841429550055694e-19

R28_170 V28 V170 2218.5964683800166
L28_170 V28 V170 6.65241788302659e-12
C28_170 V28 V170 1.6189912275264499e-19

R28_171 V28 V171 1687.8578381060659
L28_171 V28 V171 2.4025835446399606e-12
C28_171 V28 V171 6.854767856793805e-20

R28_172 V28 V172 2270.8162227023518
L28_172 V28 V172 -1.0537096071074686e-12
C28_172 V28 V172 5.2875415863142785e-20

R28_173 V28 V173 5258.261764798916
L28_173 V28 V173 3.77163062915379e-12
C28_173 V28 V173 3.25023830160346e-19

R28_174 V28 V174 1198.6636239782572
L28_174 V28 V174 9.9642437379213e-13
C28_174 V28 V174 1.4765081137539163e-20

R28_175 V28 V175 -2954.304987370668
L28_175 V28 V175 1.4810730868546721e-12
C28_175 V28 V175 2.5008924918706913e-19

R28_176 V28 V176 2018.1195352401226
L28_176 V28 V176 5.965634285072719e-13
C28_176 V28 V176 7.193093641940098e-19

R28_177 V28 V177 -4314.292698606439
L28_177 V28 V177 -2.456367842388697e-12
C28_177 V28 V177 -1.7340480677434132e-19

R28_178 V28 V178 -1234.2299937921919
L28_178 V28 V178 -1.3212268602477312e-12
C28_178 V28 V178 -1.1285113491506252e-19

R28_179 V28 V179 3279.8218946951415
L28_179 V28 V179 -1.0419256265735727e-12
C28_179 V28 V179 -3.3164687647934114e-19

R28_180 V28 V180 -1236.4876897300267
L28_180 V28 V180 -2.1324908077930947e-12
C28_180 V28 V180 -6.543652252265653e-19

R28_181 V28 V181 2809.7197840480753
L28_181 V28 V181 8.82501530746162e-12
C28_181 V28 V181 -3.047152178906295e-19

R28_182 V28 V182 2586.7169953005787
L28_182 V28 V182 3.388468034284525e-12
C28_182 V28 V182 9.51746598214313e-20

R28_183 V28 V183 -2114.4012281152272
L28_183 V28 V183 -2.073240244228395e-12
C28_183 V28 V183 -1.512993367391875e-19

R28_184 V28 V184 -3364.7414074661524
L28_184 V28 V184 -6.487059020248858e-13
C28_184 V28 V184 4.495069229887909e-20

R28_185 V28 V185 -1905.700297055491
L28_185 V28 V185 -2.2810348732712337e-12
C28_185 V28 V185 2.7072652556515394e-19

R28_186 V28 V186 6578.42491188554
L28_186 V28 V186 -1.4697346064198892e-12
C28_186 V28 V186 -1.7813399820656426e-19

R28_187 V28 V187 12378.660835307495
L28_187 V28 V187 2.4290514973028937e-12
C28_187 V28 V187 2.9900600056914895e-19

R28_188 V28 V188 712.8730775045971
L28_188 V28 V188 4.855269486659051e-13
C28_188 V28 V188 3.7078549034084386e-19

R28_189 V28 V189 12706.8104619309
L28_189 V28 V189 3.0820828867902328e-12
C28_189 V28 V189 7.223242748963692e-20

R28_190 V28 V190 -2262.2035448506367
L28_190 V28 V190 1.3069720953054538e-11
C28_190 V28 V190 -1.4422861641840087e-19

R28_191 V28 V191 8064.6140243001655
L28_191 V28 V191 1.066473964071743e-12
C28_191 V28 V191 1.5658857129518125e-19

R28_192 V28 V192 -2714.266663276548
L28_192 V28 V192 -4.993536825135162e-12
C28_192 V28 V192 -3.088586432237768e-19

R28_193 V28 V193 1720.9633480375562
L28_193 V28 V193 2.02307616167897e-12
C28_193 V28 V193 -6.331784048273882e-20

R28_194 V28 V194 -13862.152712193109
L28_194 V28 V194 1.9965356848329906e-11
C28_194 V28 V194 -2.338743170313892e-19

R28_195 V28 V195 -2283.534169567849
L28_195 V28 V195 -7.330354342241251e-13
C28_195 V28 V195 -5.953120703111094e-19

R28_196 V28 V196 -1064.7591717313817
L28_196 V28 V196 -7.003263555574066e-12
C28_196 V28 V196 6.0870312435557585e-19

R28_197 V28 V197 -4576.971751078098
L28_197 V28 V197 -1.4627853228217029e-12
C28_197 V28 V197 -1.4328362938102122e-19

R28_198 V28 V198 -8559.470155730467
L28_198 V28 V198 -6.5377563545946035e-12
C28_198 V28 V198 -9.869495153802302e-20

R28_199 V28 V199 -3658.8591822636395
L28_199 V28 V199 -5.019394147450189e-12
C28_199 V28 V199 -1.2633527023426569e-20

R28_200 V28 V200 874.2518652900089
L28_200 V28 V200 -6.609162098075789e-12
C28_200 V28 V200 -9.064833116701218e-20

R29_29 V29 0 86.29456917316487
L29_29 V29 0 1.8723277658857307e-13
C29_29 V29 0 7.603801656469119e-19

R29_30 V29 V30 -3526.706211873612
L29_30 V29 V30 -3.871557060594076e-12
C29_30 V29 V30 -6.786953152040003e-20

R29_31 V29 V31 -4115.202920249547
L29_31 V29 V31 -3.811276232026477e-12
C29_31 V29 V31 -3.870955144081322e-20

R29_32 V29 V32 -2287.6978481878464
L29_32 V29 V32 -2.612983616676409e-12
C29_32 V29 V32 -4.030426044530115e-20

R29_33 V29 V33 -987.0737485521158
L29_33 V29 V33 5.4897942291070844e-12
C29_33 V29 V33 1.764612122014989e-19

R29_34 V29 V34 6984.641476897509
L29_34 V29 V34 -8.007115982419006e-12
C29_34 V29 V34 -1.0672429417265808e-19

R29_35 V29 V35 2915.956043475356
L29_35 V29 V35 6.633267481457177e-12
C29_35 V29 V35 3.7054362055210764e-20

R29_36 V29 V36 1909.5830117309065
L29_36 V29 V36 4.136918332579933e-12
C29_36 V29 V36 8.813242937258673e-20

R29_37 V29 V37 689.777280150927
L29_37 V29 V37 8.319686999307339e-13
C29_37 V29 V37 2.8255023604462887e-19

R29_38 V29 V38 4239.956368445838
L29_38 V29 V38 1.905219186091817e-12
C29_38 V29 V38 1.5549020316328357e-19

R29_39 V29 V39 4167.6020322176055
L29_39 V29 V39 3.701835405011268e-12
C29_39 V29 V39 -1.7499727275500617e-20

R29_40 V29 V40 2542.228117900413
L29_40 V29 V40 2.7190843865533644e-12
C29_40 V29 V40 -2.2134132478592914e-20

R29_41 V29 V41 2010.876496698658
L29_41 V29 V41 -6.443295383034984e-12
C29_41 V29 V41 -2.0227532102024651e-19

R29_42 V29 V42 3650.945977711819
L29_42 V29 V42 1.5854639059691442e-11
C29_42 V29 V42 -1.989684855896556e-20

R29_43 V29 V43 2612.136429671306
L29_43 V29 V43 5.1710337812678995e-12
C29_43 V29 V43 2.820879688011829e-20

R29_44 V29 V44 2131.6941443282244
L29_44 V29 V44 6.1717571724482184e-12
C29_44 V29 V44 2.741318827248611e-20

R29_45 V29 V45 -496.65143757528193
L29_45 V29 V45 -9.751912401217412e-13
C29_45 V29 V45 -1.4155780683322303e-19

R29_46 V29 V46 -16961.444176831785
L29_46 V29 V46 -3.096286345772949e-12
C29_46 V29 V46 -1.4983892860902114e-19

R29_47 V29 V47 37384.9510526088
L29_47 V29 V47 -4.2711446294667625e-12
C29_47 V29 V47 -2.5572622991091067e-20

R29_48 V29 V48 -5354.121936947378
L29_48 V29 V48 -2.2008400047474494e-12
C29_48 V29 V48 -6.530971572743206e-20

R29_49 V29 V49 -495.44416876367944
L29_49 V29 V49 5.2755425528028226e-11
C29_49 V29 V49 1.0390999063000214e-19

R29_50 V29 V50 5398.053744261737
L29_50 V29 V50 7.757863866265896e-12
C29_50 V29 V50 1.1236622621545314e-19

R29_51 V29 V51 11789.19383946419
L29_51 V29 V51 -5.439923034134348e-12
C29_51 V29 V51 -1.6024543611110027e-20

R29_52 V29 V52 4215.1522187676
L29_52 V29 V52 -7.20587224529946e-12
C29_52 V29 V52 1.6334524959874174e-20

R29_53 V29 V53 -1168.8978615185517
L29_53 V29 V53 -4.15371057555366e-12
C29_53 V29 V53 -1.2061892401841817e-20

R29_54 V29 V54 -4157.128414023378
L29_54 V29 V54 -1.9125722851408625e-11
C29_54 V29 V54 8.861400469312868e-21

R29_55 V29 V55 -3173.691048068711
L29_55 V29 V55 -2.7412011924763436e-11
C29_55 V29 V55 3.4556358070891245e-20

R29_56 V29 V56 -5472.790777900039
L29_56 V29 V56 8.238407026569192e-12
C29_56 V29 V56 8.017017541514763e-20

R29_57 V29 V57 4275.009998203228
L29_57 V29 V57 1.4209300601389548e-12
C29_57 V29 V57 -2.01080682811145e-20

R29_58 V29 V58 2561.347793701203
L29_58 V29 V58 3.873063550643042e-12
C29_58 V29 V58 -1.1597597625555984e-20

R29_59 V29 V59 1794.6469518199947
L29_59 V29 V59 2.9371522918901512e-12
C29_59 V29 V59 -1.9434317724667217e-20

R29_60 V29 V60 1239.7716733867712
L29_60 V29 V60 2.1113306614531246e-12
C29_60 V29 V60 -1.8041271852068514e-20

R29_61 V29 V61 3119.8971437724745
L29_61 V29 V61 -2.4870252114983584e-12
C29_61 V29 V61 1.0122962294056708e-20

R29_62 V29 V62 -407815.5848570324
L29_62 V29 V62 1.2086680677624805e-11
C29_62 V29 V62 9.497933580728782e-21

R29_63 V29 V63 15524.103932103593
L29_63 V29 V63 5.651891779785151e-12
C29_63 V29 V63 2.798784940365666e-20

R29_64 V29 V64 -15713.0539981992
L29_64 V29 V64 5.021973616079367e-11
C29_64 V29 V64 2.1080021470241036e-20

R29_65 V29 V65 -643.790577747718
L29_65 V29 V65 -2.0575215778614233e-12
C29_65 V29 V65 -1.6718449995057972e-19

R29_66 V29 V66 4989.894751768425
L29_66 V29 V66 -6.8921475976541575e-12
C29_66 V29 V66 -1.0040648258121145e-19

R29_67 V29 V67 6138.345036821022
L29_67 V29 V67 -4.20164399426693e-12
C29_67 V29 V67 -5.378744128707181e-20

R29_68 V29 V68 17443.638089632354
L29_68 V29 V68 -1.7554828050692238e-12
C29_68 V29 V68 -1.16815331034256e-19

R29_69 V29 V69 -1350.0112143849572
L29_69 V29 V69 6.34063996059419e-12
C29_69 V29 V69 3.0361384338362885e-19

R29_70 V29 V70 7666.588637705699
L29_70 V29 V70 5.933519912966276e-11
C29_70 V29 V70 8.243179248694578e-20

R29_71 V29 V71 33072.09301560285
L29_71 V29 V71 -4.317302730735559e-12
C29_71 V29 V71 -1.629578973112358e-20

R29_72 V29 V72 13132.459041994849
L29_72 V29 V72 -7.451710238297975e-12
C29_72 V29 V72 2.3182513372744616e-20

R29_73 V29 V73 -2599.687856761795
L29_73 V29 V73 -4.4734980148975295e-10
C29_73 V29 V73 -1.1972612056177288e-19

R29_74 V29 V74 -4272.345314164853
L29_74 V29 V74 2.7415652016619412e-12
C29_74 V29 V74 1.2282988582328687e-19

R29_75 V29 V75 -4696.624830083305
L29_75 V29 V75 2.8904668343500987e-12
C29_75 V29 V75 8.17143982635621e-20

R29_76 V29 V76 137087.43450449262
L29_76 V29 V76 1.357692087503479e-12
C29_76 V29 V76 1.9365742678218696e-19

R29_77 V29 V77 3016.6512732184588
L29_77 V29 V77 3.4166740185401614e-12
C29_77 V29 V77 -1.6960952144353996e-19

R29_78 V29 V78 -9454.78839199803
L29_78 V29 V78 -5.629999348263966e-12
C29_78 V29 V78 -7.388086150021694e-20

R29_79 V29 V79 8110.623682863841
L29_79 V29 V79 -1.1827635866590152e-10
C29_79 V29 V79 -5.847463335082394e-20

R29_80 V29 V80 9916.841763056413
L29_80 V29 V80 -3.5562823702051567e-12
C29_80 V29 V80 -1.560053051091032e-19

R29_81 V29 V81 -373.5091317727974
L29_81 V29 V81 -1.3122754247542582e-12
C29_81 V29 V81 9.351087571843275e-21

R29_82 V29 V82 2566.933838236218
L29_82 V29 V82 -4.47411266313867e-12
C29_82 V29 V82 -1.6148856382097919e-19

R29_83 V29 V83 1390.3437478570202
L29_83 V29 V83 4.590308217390325e-11
C29_83 V29 V83 -2.6298685611506454e-20

R29_84 V29 V84 1559.9435725998278
L29_84 V29 V84 -4.249652820722512e-12
C29_84 V29 V84 -1.0276145516762159e-19

R29_85 V29 V85 -23656.393585960195
L29_85 V29 V85 -1.7613924755999215e-11
C29_85 V29 V85 8.172262388001075e-21

R29_86 V29 V86 1029.506428833086
L29_86 V29 V86 5.509863338533135e-12
C29_86 V29 V86 6.603491264097308e-20

R29_87 V29 V87 3931.719837175872
L29_87 V29 V87 5.874982283408992e-12
C29_87 V29 V87 1.354551743128096e-19

R29_88 V29 V88 3189.5073700531093
L29_88 V29 V88 3.896941036484056e-12
C29_88 V29 V88 2.0160232410894745e-19

R29_89 V29 V89 -3648.1744689511
L29_89 V29 V89 1.190593747215378e-11
C29_89 V29 V89 1.6370586138357814e-19

R29_90 V29 V90 -1674.5606434048618
L29_90 V29 V90 2.3520969357316267e-12
C29_90 V29 V90 2.594760097077382e-19

R29_91 V29 V91 -2207.436765602059
L29_91 V29 V91 -1.5779058898444655e-12
C29_91 V29 V91 -1.797168087293268e-19

R29_92 V29 V92 -5406.990600298239
L29_92 V29 V92 -2.1923645429687693e-12
C29_92 V29 V92 -1.2594366782225933e-19

R29_93 V29 V93 -757.1855811146938
L29_93 V29 V93 8.826366450156595e-12
C29_93 V29 V93 -3.908701094218811e-20

R29_94 V29 V94 -1782.3146165102403
L29_94 V29 V94 -3.583650739314684e-12
C29_94 V29 V94 -1.5164858512390857e-19

R29_95 V29 V95 -4038.7690199846106
L29_95 V29 V95 6.910108393643643e-12
C29_95 V29 V95 -7.656285590294621e-20

R29_96 V29 V96 -2618.3808424715457
L29_96 V29 V96 4.465038509215242e-12
C29_96 V29 V96 -1.0074419095722723e-19

R29_97 V29 V97 -862.9774572671131
L29_97 V29 V97 -2.3870753437857345e-11
C29_97 V29 V97 -3.3312541690939165e-19

R29_98 V29 V98 706.5374840257726
L29_98 V29 V98 -7.337382820625927e-12
C29_98 V29 V98 -1.5465668471308143e-19

R29_99 V29 V99 630.3235650956645
L29_99 V29 V99 1.5783188708786045e-12
C29_99 V29 V99 2.57933491213926e-19

R29_100 V29 V100 619.8643106317778
L29_100 V29 V100 3.5160212411307066e-12
C29_100 V29 V100 1.796171428470711e-19

R29_101 V29 V101 1913.8747035789577
L29_101 V29 V101 -6.4990853140249156e-12
C29_101 V29 V101 1.571945796773928e-19

R29_102 V29 V102 10035.54468217227
L29_102 V29 V102 2.769184583115911e-12
C29_102 V29 V102 1.276801660879406e-19

R29_103 V29 V103 -21974.958723242107
L29_103 V29 V103 -9.591502544665232e-12
C29_103 V29 V103 -3.5479861183680976e-20

R29_104 V29 V104 7069.686252465758
L29_104 V29 V104 -8.845276279023623e-12
C29_104 V29 V104 -4.245710323755116e-20

R29_105 V29 V105 -305.83857382369354
L29_105 V29 V105 -2.3951689488837117e-12
C29_105 V29 V105 1.2894471355130357e-19

R29_106 V29 V106 2214.660542439011
L29_106 V29 V106 -1.8083176550537237e-10
C29_106 V29 V106 1.4233731883444757e-19

R29_107 V29 V107 -6457.867894032875
L29_107 V29 V107 -3.2734449643240026e-12
C29_107 V29 V107 -1.363689587980188e-19

R29_108 V29 V108 -3242.1564218504104
L29_108 V29 V108 -1.604080334781792e-11
C29_108 V29 V108 1.275734186554002e-20

R29_109 V29 V109 1338.168520591121
L29_109 V29 V109 -4.627826925708755e-12
C29_109 V29 V109 -1.5956143322381523e-19

R29_110 V29 V110 -3648.1999612192412
L29_110 V29 V110 -1.578228851118685e-11
C29_110 V29 V110 -8.09677096537736e-20

R29_111 V29 V111 6452.406420970619
L29_111 V29 V111 -3.159436152100237e-12
C29_111 V29 V111 6.198325210768186e-21

R29_112 V29 V112 3367.491016763316
L29_112 V29 V112 -3.9708593017861135e-12
C29_112 V29 V112 -6.097861531722713e-20

R29_113 V29 V113 -1785.219110402355
L29_113 V29 V113 2.151594778923464e-12
C29_113 V29 V113 -3.796100938428171e-20

R29_114 V29 V114 10318.63649399788
L29_114 V29 V114 -2.3151236040349715e-10
C29_114 V29 V114 -1.658850746990697e-19

R29_115 V29 V115 4802.44824869444
L29_115 V29 V115 1.6639728556088472e-12
C29_115 V29 V115 1.0429002216058217e-19

R29_116 V29 V116 15360.306699319248
L29_116 V29 V116 2.373749443410957e-12
C29_116 V29 V116 3.6536655455614595e-21

R29_117 V29 V117 -674.5397333756518
L29_117 V29 V117 4.234294377661134e-12
C29_117 V29 V117 4.26791009042012e-20

R29_118 V29 V118 7137.211442887818
L29_118 V29 V118 -1.92003648328338e-11
C29_118 V29 V118 1.7567559527996316e-19

R29_119 V29 V119 2616.937561704952
L29_119 V29 V119 -2.3186959969885966e-11
C29_119 V29 V119 4.065789535988347e-20

R29_120 V29 V120 1535.8398493278157
L29_120 V29 V120 1.0506949723946229e-11
C29_120 V29 V120 1.5284230594629191e-19

R29_121 V29 V121 3571.2471965531545
L29_121 V29 V121 -1.6740129552094954e-12
C29_121 V29 V121 -1.0004929645924055e-20

R29_122 V29 V122 2408.5582388237194
L29_122 V29 V122 -3.5249914274925383e-11
C29_122 V29 V122 -2.768316021982649e-20

R29_123 V29 V123 -6231.518470327141
L29_123 V29 V123 -2.891254520810362e-12
C29_123 V29 V123 -1.2611247026758034e-19

R29_124 V29 V124 -3109.884198943803
L29_124 V29 V124 -1.862345065668824e-12
C29_124 V29 V124 -2.0272782389427544e-19

R29_125 V29 V125 -451.0921160216522
L29_125 V29 V125 -1.6314945391308936e-12
C29_125 V29 V125 -2.752618961255708e-20

R29_126 V29 V126 -16897.895749689153
L29_126 V29 V126 -4.6306383836781065e-12
C29_126 V29 V126 -1.098863451499951e-19

R29_127 V29 V127 -6735.570035123649
L29_127 V29 V127 7.880393273442551e-12
C29_127 V29 V127 -1.0435524318975037e-20

R29_128 V29 V128 -2055.552963860647
L29_128 V29 V128 9.173593168955946e-12
C29_128 V29 V128 -9.589428757913298e-21

R29_129 V29 V129 5368.072817883426
L29_129 V29 V129 5.023364245276433e-12
C29_129 V29 V129 -1.2286434526818e-19

R29_130 V29 V130 -4534.650519055787
L29_130 V29 V130 2.7381212184722314e-12
C29_130 V29 V130 1.3700486521235053e-19

R29_131 V29 V131 5372.189965619541
L29_131 V29 V131 2.7571175830669843e-11
C29_131 V29 V131 9.801612124347471e-20

R29_132 V29 V132 1138.701033925651
L29_132 V29 V132 3.5625418904365964e-12
C29_132 V29 V132 1.8969967505449994e-19

R29_133 V29 V133 647.0857184961015
L29_133 V29 V133 1.6610100972380297e-12
C29_133 V29 V133 2.421920708937693e-19

R29_134 V29 V134 919.7612593864097
L29_134 V29 V134 -7.294514923942452e-12
C29_134 V29 V134 -7.176430200427254e-20

R29_135 V29 V135 -27203.49496042499
L29_135 V29 V135 -5.750591935816413e-12
C29_135 V29 V135 -6.35114577482333e-20

R29_136 V29 V136 -3852.3489850727187
L29_136 V29 V136 -2.9199989478451063e-12
C29_136 V29 V136 -1.5569504197571693e-19

R29_137 V29 V137 -491.55394908432606
L29_137 V29 V137 3.533979823955957e-12
C29_137 V29 V137 2.89388056983269e-20

R29_138 V29 V138 -687.7897693807273
L29_138 V29 V138 -6.084548593627447e-12
C29_138 V29 V138 -3.91945628836395e-20

R29_139 V29 V139 3401.649176025594
L29_139 V29 V139 3.272428072817061e-12
C29_139 V29 V139 1.0739639733018403e-19

R29_140 V29 V140 5243.615409256992
L29_140 V29 V140 2.1547992354413046e-12
C29_140 V29 V140 1.2189037852853114e-19

R29_141 V29 V141 956.4994022306454
L29_141 V29 V141 -8.529016032913507e-13
C29_141 V29 V141 -3.8275377176535155e-19

R29_142 V29 V142 1324.9150231051913
L29_142 V29 V142 2.9453163040005404e-12
C29_142 V29 V142 3.580037505431345e-20

R29_143 V29 V143 2758.0101980891613
L29_143 V29 V143 -2.8494868822683327e-11
C29_143 V29 V143 -8.554518299288664e-20

R29_144 V29 V144 1514.9776922175572
L29_144 V29 V144 -1.645930945733011e-11
C29_144 V29 V144 -2.806508020647998e-20

R29_145 V29 V145 -403.68357791085197
L29_145 V29 V145 -1.9626703237362707e-12
C29_145 V29 V145 -1.6206742794719476e-20

R29_146 V29 V146 1088.900004417815
L29_146 V29 V146 -5.005943396275939e-12
C29_146 V29 V146 3.0081856308146554e-20

R29_147 V29 V147 -1817.8228054612214
L29_147 V29 V147 -1.985755064149365e-12
C29_147 V29 V147 -1.2373502013141936e-19

R29_148 V29 V148 -967.4757112665615
L29_148 V29 V148 -1.489440089436576e-12
C29_148 V29 V148 -1.12839332707104e-19

R29_149 V29 V149 241.91000259924857
L29_149 V29 V149 9.10918552947873e-13
C29_149 V29 V149 4.343210842934858e-19

R29_150 V29 V150 -976.7624673949795
L29_150 V29 V150 -2.4971752448217817e-12
C29_150 V29 V150 -1.481026498366164e-19

R29_151 V29 V151 -1883.3797268379988
L29_151 V29 V151 -8.883688029489303e-12
C29_151 V29 V151 1.1947636360296775e-19

R29_152 V29 V152 1694.143860441496
L29_152 V29 V152 5.4159656019649626e-12
C29_152 V29 V152 2.9509550404073364e-20

R29_153 V29 V153 -375.0696145415432
L29_153 V29 V153 1.5574620525452784e-12
C29_153 V29 V153 2.912405100684126e-20

R29_154 V29 V154 3537.289805006523
L29_154 V29 V154 2.035794605608034e-12
C29_154 V29 V154 1.0836597178761365e-19

R29_155 V29 V155 883.8689458624307
L29_155 V29 V155 1.495627827845716e-12
C29_155 V29 V155 8.62682767649892e-20

R29_156 V29 V156 14345.859810618525
L29_156 V29 V156 2.777261861013888e-12
C29_156 V29 V156 1.0856459191473672e-19

R29_157 V29 V157 -416.28601537801063
L29_157 V29 V157 -1.503984973926159e-12
C29_157 V29 V157 -3.448231645366288e-19

R29_158 V29 V158 2990.354269720999
L29_158 V29 V158 5.056236458082453e-12
C29_158 V29 V158 4.967840561018993e-21

R29_159 V29 V159 -21389.52326139703
L29_159 V29 V159 1.044678243052111e-11
C29_159 V29 V159 -5.132988909247347e-20

R29_160 V29 V160 2899.78715675046
L29_160 V29 V160 5.340881277588372e-12
C29_160 V29 V160 -5.251055113324086e-20

R29_161 V29 V161 -954.6117268949831
L29_161 V29 V161 -2.954700790870548e-12
C29_161 V29 V161 -5.334868602525178e-20

R29_162 V29 V162 3556.0400676263794
L29_162 V29 V162 7.614621796422267e-12
C29_162 V29 V162 6.917317746468646e-20

R29_163 V29 V163 884.5649404389509
L29_163 V29 V163 1.7113762341343678e-10
C29_163 V29 V163 -2.2416485758197616e-20

R29_164 V29 V164 2030.862437012753
L29_164 V29 V164 -4.342863507042044e-12
C29_164 V29 V164 5.718879863291007e-20

R29_165 V29 V165 -724.5505291934044
L29_165 V29 V165 -1.0026293734962472e-12
C29_165 V29 V165 7.986887251962791e-20

R29_166 V29 V166 793.10766238935
L29_166 V29 V166 -1.681734161094139e-12
C29_166 V29 V166 -6.216779398863304e-20

R29_167 V29 V167 -12359.616130443246
L29_167 V29 V167 -3.8892144500489025e-12
C29_167 V29 V167 7.839196578317356e-21

R29_168 V29 V168 986.1990770999896
L29_168 V29 V168 -5.117704478159954e-12
C29_168 V29 V168 -4.565555388161619e-20

R29_169 V29 V169 10735.864891108824
L29_169 V29 V169 1.5579186020210925e-12
C29_169 V29 V169 -3.724906623026793e-20

R29_170 V29 V170 -451.22895012234164
L29_170 V29 V170 6.375055574540118e-12
C29_170 V29 V170 1.0389543212185183e-19

R29_171 V29 V171 -584.7416658984486
L29_171 V29 V171 3.226616626442153e-11
C29_171 V29 V171 1.0658130412803352e-19

R29_172 V29 V172 -770.505772520065
L29_172 V29 V172 4.430353060459558e-11
C29_172 V29 V172 5.3993723718041925e-20

R29_173 V29 V173 -450.5519134532665
L29_173 V29 V173 1.63781545741022e-12
C29_173 V29 V173 3.3788339969740005e-20

R29_174 V29 V174 740.3806124791171
L29_174 V29 V174 1.1397142583849316e-12
C29_174 V29 V174 -8.083891708694908e-20

R29_175 V29 V175 549.8911018562085
L29_175 V29 V175 1.3624606009446138e-12
C29_175 V29 V175 8.585975779625403e-20

R29_176 V29 V176 701.1635912868506
L29_176 V29 V176 1.0763523430783347e-12
C29_176 V29 V176 1.1306160704154524e-19

R29_177 V29 V177 712.4214789720272
L29_177 V29 V177 -1.8245655083765543e-12
C29_177 V29 V177 3.2373607961212344e-20

R29_178 V29 V178 -7409.262127568944
L29_178 V29 V178 -2.8058399349021755e-12
C29_178 V29 V178 -5.0000047056216875e-20

R29_179 V29 V179 -5869.394397203703
L29_179 V29 V179 -2.8782162868876453e-12
C29_179 V29 V179 -2.0273902345811683e-19

R29_180 V29 V180 -1778.231820581018
L29_180 V29 V180 -1.862308596938691e-12
C29_180 V29 V180 -1.9480322750619435e-19

R29_181 V29 V181 792.959319911328
L29_181 V29 V181 -5.7862577355735896e-12
C29_181 V29 V181 -7.630050362806713e-20

R29_182 V29 V182 -1241.5202611350837
L29_182 V29 V182 -1.8013446189957653e-11
C29_182 V29 V182 8.775835407144587e-20

R29_183 V29 V183 -2024.8580587401598
L29_183 V29 V183 -3.1921826927981017e-12
C29_183 V29 V183 -4.2805006705534003e-20

R29_184 V29 V184 -1950.578959228624
L29_184 V29 V184 -2.128604472129594e-12
C29_184 V29 V184 8.781593118470164e-22

R29_185 V29 V185 -214.90141526881703
L29_185 V29 V185 1.6689226594864398e-10
C29_185 V29 V185 -2.6673011846333864e-21

R29_186 V29 V186 549.297864155543
L29_186 V29 V186 -1.782646103696814e-12
C29_186 V29 V186 -5.386410064512051e-20

R29_187 V29 V187 2268.518525987994
L29_187 V29 V187 1.005042518175047e-09
C29_187 V29 V187 1.4798220451213597e-19

R29_188 V29 V188 3097.6795706706157
L29_188 V29 V188 5.00804995082792e-12
C29_188 V29 V188 1.2586512206922975e-19

R29_189 V29 V189 223.48586679377578
L29_189 V29 V189 2.306690173569635e-12
C29_189 V29 V189 2.548682501346257e-20

R29_190 V29 V190 -3490.669666337121
L29_190 V29 V190 4.411457420906438e-12
C29_190 V29 V190 -5.670721878996003e-20

R29_191 V29 V191 -689.9596933400449
L29_191 V29 V191 2.21426091597034e-12
C29_191 V29 V191 8.14499253938219e-20

R29_192 V29 V192 -992.3239018284481
L29_192 V29 V192 1.920050673720563e-12
C29_192 V29 V192 2.6828547760091357e-20

R29_193 V29 V193 1528.331029977389
L29_193 V29 V193 -1.6099400785690998e-11
C29_193 V29 V193 1.639684277973826e-20

R29_194 V29 V194 -574.4144818388147
L29_194 V29 V194 1.2461393344304893e-12
C29_194 V29 V194 -5.132542926037081e-20

R29_195 V29 V195 7172.062360009146
L29_195 V29 V195 -3.0380873983732497e-12
C29_195 V29 V195 -1.656878067363527e-19

R29_196 V29 V196 5668.60486065036
L29_196 V29 V196 2.0034218632880487e-11
C29_196 V29 V196 -6.595305367380109e-20

R29_197 V29 V197 -365.9801217005953
L29_197 V29 V197 -4.058372706368119e-12
C29_197 V29 V197 -3.694785453113627e-20

R29_198 V29 V198 675.1150169989719
L29_198 V29 V198 -3.0949974728568193e-12
C29_198 V29 V198 3.428714977156195e-20

R29_199 V29 V199 447.5201296295659
L29_199 V29 V199 -4.1195669408815275e-12
C29_199 V29 V199 -1.840216211403477e-20

R29_200 V29 V200 599.5503737406185
L29_200 V29 V200 -1.6021186094028868e-12
C29_200 V29 V200 -2.666728044337039e-20

R30_30 V30 0 194.44537653932466
L30_30 V30 0 5.279043889881512e-13
C30_30 V30 0 -2.217921104568986e-19

R30_31 V30 V31 -3372.1731410901198
L30_31 V30 V31 -3.929293743543098e-12
C30_31 V30 V31 -1.361692318129793e-19

R30_32 V30 V32 -2834.2996121560127
L30_32 V30 V32 -3.254559391975547e-12
C30_32 V30 V32 -1.4375946435355567e-19

R30_33 V30 V33 -89975.7688158915
L30_33 V30 V33 -3.855570485621083e-12
C30_33 V30 V33 -1.206402938941052e-19

R30_34 V30 V34 1565.1606091127667
L30_34 V30 V34 3.6263764088520847e-12
C30_34 V30 V34 2.2839153601897224e-19

R30_35 V30 V35 4106.430086321542
L30_35 V30 V35 -1.749979642425427e-11
C30_35 V30 V35 -5.861001619107505e-20

R30_36 V30 V36 2663.571528442381
L30_36 V30 V36 -1.0823331854554625e-11
C30_36 V30 V36 -7.27773868959095e-20

R30_37 V30 V37 9650.662130054596
L30_37 V30 V37 3.4487785188167087e-12
C30_37 V30 V37 1.1522334641431315e-19

R30_38 V30 V38 1881.6136817974193
L30_38 V30 V38 9.111796452313892e-13
C30_38 V30 V38 7.049015735435365e-19

R30_39 V30 V39 4354.027437813662
L30_39 V30 V39 5.2654823184360985e-12
C30_39 V30 V39 1.322826640838408e-19

R30_40 V30 V40 3037.988144589801
L30_40 V30 V40 4.74455552162164e-12
C30_40 V30 V40 1.5260194432366792e-19

R30_41 V30 V41 -9007.972633879817
L30_41 V30 V41 2.8664115478311636e-11
C30_41 V30 V41 -7.377818491391985e-20

R30_42 V30 V42 1906.9223553399715
L30_42 V30 V42 -1.2056778359263276e-12
C30_42 V30 V42 -5.974619231099622e-19

R30_43 V30 V43 35829.80635174549
L30_43 V30 V43 -2.271506756024136e-11
C30_43 V30 V43 -1.4509582825229582e-19

R30_44 V30 V44 -52018.710933209746
L30_44 V30 V44 -1.8291185720029237e-11
C30_44 V30 V44 -1.7384932829495724e-19

R30_45 V30 V45 -4114.686520262453
L30_45 V30 V45 -1.308594017705758e-10
C30_45 V30 V45 1.1097947442545604e-19

R30_46 V30 V46 -1211.3224048225786
L30_46 V30 V46 -1.9425395259669047e-12
C30_46 V30 V46 -1.9738187501781947e-19

R30_47 V30 V47 -9643.154189471788
L30_47 V30 V47 5.815855347048731e-10
C30_47 V30 V47 2.2925359682658758e-20

R30_48 V30 V48 -4201.688501162733
L30_48 V30 V48 -2.1213835629139315e-11
C30_48 V30 V48 1.1729237888994286e-20

R30_49 V30 V49 -24771.09161596599
L30_49 V30 V49 -1.537527667573781e-11
C30_49 V30 V49 3.768398901982543e-20

R30_50 V30 V50 -1520.520658303751
L30_50 V30 V50 1.7885739176326793e-12
C30_50 V30 V50 4.439156385853348e-19

R30_51 V30 V51 -23024.951805081073
L30_51 V30 V51 9.262275659845012e-12
C30_51 V30 V51 1.6004023503078453e-19

R30_52 V30 V52 17677.20806572264
L30_52 V30 V52 6.433102953264359e-12
C30_52 V30 V52 2.339402737029293e-19

R30_53 V30 V53 -7011.362444493635
L30_53 V30 V53 -1.862263351687807e-12
C30_53 V30 V53 -2.7492308060919127e-19

R30_54 V30 V54 2179.800314561399
L30_54 V30 V54 4.925563399683871e-12
C30_54 V30 V54 -3.523775027976215e-21

R30_55 V30 V55 11851.259394489123
L30_55 V30 V55 -3.6464683646101335e-12
C30_55 V30 V55 -1.9673887326527303e-19

R30_56 V30 V56 3400.432739246806
L30_56 V30 V56 -3.4671546932107585e-12
C30_56 V30 V56 -2.1430741854060193e-19

R30_57 V30 V57 48673.54686009687
L30_57 V30 V57 2.067239119925459e-12
C30_57 V30 V57 1.6097408703584468e-19

R30_58 V30 V58 -6368.73904298753
L30_58 V30 V58 -2.096038964110213e-12
C30_58 V30 V58 -1.7013907804244985e-19

R30_59 V30 V59 13197.511594032658
L30_59 V30 V59 1.2657665882035904e-11
C30_59 V30 V59 -6.486465780310826e-20

R30_60 V30 V60 8093.194105549665
L30_60 V30 V60 1.2180228667959579e-11
C30_60 V30 V60 -1.1124201381130219e-19

R30_61 V30 V61 -37691.230484511856
L30_61 V30 V61 1.4641692023992905e-11
C30_61 V30 V61 1.1487577487025336e-19

R30_62 V30 V62 1788.853394605614
L30_62 V30 V62 -7.616418667293654e-12
C30_62 V30 V62 -9.687997183066852e-20

R30_63 V30 V63 -277932.1971474435
L30_63 V30 V63 2.8199630723011554e-12
C30_63 V30 V63 2.302156025268933e-19

R30_64 V30 V64 -6988.418751425199
L30_64 V30 V64 2.2817608737437468e-12
C30_64 V30 V64 3.382948536255705e-19

R30_65 V30 V65 -6086.586609156729
L30_65 V30 V65 -3.5966953966537462e-12
C30_65 V30 V65 -1.7708289153948848e-19

R30_66 V30 V66 -1488.4923740213271
L30_66 V30 V66 2.1471116129732308e-12
C30_66 V30 V66 1.2545762172203296e-19

R30_67 V30 V67 808171.0842089677
L30_67 V30 V67 -7.102757203034432e-12
C30_67 V30 V67 -9.74834855469753e-20

R30_68 V30 V68 -9530.120139326944
L30_68 V30 V68 -4.07928733249631e-12
C30_68 V30 V68 -1.2187404833037998e-19

R30_69 V30 V69 10526.450748068595
L30_69 V30 V69 -7.875176880723166e-12
C30_69 V30 V69 -1.0929130805113132e-20

R30_70 V30 V70 -1944.0875069206286
L30_70 V30 V70 -1.7746360468410382e-11
C30_70 V30 V70 1.8358546830082142e-19

R30_71 V30 V71 -10759.43180476891
L30_71 V30 V71 -4.796067062390033e-12
C30_71 V30 V71 -1.020458679308858e-19

R30_72 V30 V72 -14808.153207064834
L30_72 V30 V72 -3.098511054417968e-12
C30_72 V30 V72 -2.037285247433731e-19

R30_73 V30 V73 -2589.5880818782975
L30_73 V30 V73 1.0465787872940879e-11
C30_73 V30 V73 1.0323870464770734e-19

R30_74 V30 V74 1243.576416883698
L30_74 V30 V74 -2.041311604349637e-12
C30_74 V30 V74 -2.966474490822483e-19

R30_75 V30 V75 -11523.284861956368
L30_75 V30 V75 3.520612859546252e-12
C30_75 V30 V75 1.4691250988993422e-19

R30_76 V30 V76 4512.553677923453
L30_76 V30 V76 2.090999561573382e-12
C30_76 V30 V76 2.4506194376158006e-19

R30_77 V30 V77 5983.34617981275
L30_77 V30 V77 6.539898596548088e-12
C30_77 V30 V77 -4.0537642494567534e-20

R30_78 V30 V78 -2936.488155407331
L30_78 V30 V78 1.832983625263735e-12
C30_78 V30 V78 1.6160290378516674e-19

R30_79 V30 V79 4251.047533174294
L30_79 V30 V79 8.234306708731136e-11
C30_79 V30 V79 -2.5693163913413093e-20

R30_80 V30 V80 14190.261731755954
L30_80 V30 V80 -4.65155615978439e-11
C30_80 V30 V80 -2.5214638887554653e-20

R30_81 V30 V81 -2500.5448889641343
L30_81 V30 V81 -9.177377129742024e-12
C30_81 V30 V81 -2.4939871934524223e-21

R30_82 V30 V82 -37984.62297604624
L30_82 V30 V82 1.775052545170551e-11
C30_82 V30 V82 6.199258720057353e-20

R30_83 V30 V83 22886.72522008846
L30_83 V30 V83 -9.799291594817899e-12
C30_83 V30 V83 -7.743765739665709e-20

R30_84 V30 V84 -11563.956296868279
L30_84 V30 V84 -6.6882243831063426e-12
C30_84 V30 V84 -1.0734152351124298e-19

R30_85 V30 V85 5977.04884065982
L30_85 V30 V85 -2.0495971398447193e-11
C30_85 V30 V85 5.7344144938826985e-21

R30_86 V30 V86 -1160.0873313467741
L30_86 V30 V86 -1.8551477874393256e-12
C30_86 V30 V86 -1.8496363587663642e-19

R30_87 V30 V87 -438909.5966430493
L30_87 V30 V87 5.03620280507091e-12
C30_87 V30 V87 1.1274332002367463e-19

R30_88 V30 V88 17767.017400334626
L30_88 V30 V88 4.307828859862804e-12
C30_88 V30 V88 1.3219775481156164e-19

R30_89 V30 V89 50352.223824705274
L30_89 V30 V89 -8.466806196676048e-12
C30_89 V30 V89 -8.988090478022712e-21

R30_90 V30 V90 1389.628798327117
L30_90 V30 V90 1.803650410743219e-12
C30_90 V30 V90 1.422169075239705e-19

R30_91 V30 V91 -11333.16728752582
L30_91 V30 V91 -3.07438889978861e-12
C30_91 V30 V91 -1.4256313597842238e-19

R30_92 V30 V92 21259.705415559114
L30_92 V30 V92 -1.92405443022601e-12
C30_92 V30 V92 -1.8530278645437465e-19

R30_93 V30 V93 -2922.894494220393
L30_93 V30 V93 4.626019734925328e-12
C30_93 V30 V93 4.6953159797118e-20

R30_94 V30 V94 1192.850384058323
L30_94 V30 V94 1.365010350921582e-11
C30_94 V30 V94 -1.3165267516925065e-21

R30_95 V30 V95 -80350.62913116765
L30_95 V30 V95 1.3370993779214276e-11
C30_95 V30 V95 -7.389584092632673e-21

R30_96 V30 V96 15097.509604214983
L30_96 V30 V96 4.775460545531247e-12
C30_96 V30 V96 1.603204285224168e-20

R30_97 V30 V97 2722.01715806371
L30_97 V30 V97 1.4152046482060638e-11
C30_97 V30 V97 -2.9820286415061934e-20

R30_98 V30 V98 -890.9569849005562
L30_98 V30 V98 -2.055528852859259e-12
C30_98 V30 V98 -8.82932400563298e-20

R30_99 V30 V99 1416.2448835119353
L30_99 V30 V99 2.670857005184024e-12
C30_99 V30 V99 1.5401875501495075e-19

R30_100 V30 V100 2072.723564055718
L30_100 V30 V100 2.197794593495577e-12
C30_100 V30 V100 2.1265888516643883e-19

R30_101 V30 V101 -4158.4772778226425
L30_101 V30 V101 -5.381372067432043e-12
C30_101 V30 V101 -1.8650645758427822e-20

R30_102 V30 V102 3662.2331223337665
L30_102 V30 V102 2.6836886196773063e-12
C30_102 V30 V102 9.959639488316412e-20

R30_103 V30 V103 -2129.6217353653697
L30_103 V30 V103 -2.2914194057790452e-12
C30_103 V30 V103 -1.75218262895127e-19

R30_104 V30 V104 -1882.6654928888754
L30_104 V30 V104 -1.7581573770132834e-12
C30_104 V30 V104 -2.1982785803928017e-19

R30_105 V30 V105 -2107.2290737382173
L30_105 V30 V105 -3.8205261575464005e-12
C30_105 V30 V105 -1.436858776547139e-20

R30_106 V30 V106 -869.8126185701407
L30_106 V30 V106 -5.9281133342881564e-12
C30_106 V30 V106 -2.311372676297886e-21

R30_107 V30 V107 -5382.377529358984
L30_107 V30 V107 5.085508234678585e-12
C30_107 V30 V107 6.332853865406718e-20

R30_108 V30 V108 27196.169871633523
L30_108 V30 V108 8.596569482795693e-12
C30_108 V30 V108 4.99649357145987e-20

R30_109 V30 V109 1853.5078522239507
L30_109 V30 V109 6.786744868815921e-12
C30_109 V30 V109 1.707283841465766e-20

R30_110 V30 V110 771.7628436268974
L30_110 V30 V110 -9.294473637954391e-12
C30_110 V30 V110 -2.719598560987238e-20

R30_111 V30 V111 10858.423253320349
L30_111 V30 V111 2.3088049604306124e-11
C30_111 V30 V111 7.545740705687319e-20

R30_112 V30 V112 6184.386592278871
L30_112 V30 V112 1.077142200234292e-10
C30_112 V30 V112 4.9352310888191244e-20

R30_113 V30 V113 -3559.614916828256
L30_113 V30 V113 2.8893848871996942e-12
C30_113 V30 V113 8.75002601184502e-20

R30_114 V30 V114 1347.5425718726428
L30_114 V30 V114 6.873778353648052e-12
C30_114 V30 V114 -6.637417336963917e-20

R30_115 V30 V115 2442.6019361980666
L30_115 V30 V115 -1.1399181310934048e-11
C30_115 V30 V115 -8.0262912628191e-20

R30_116 V30 V116 5415.465856393552
L30_116 V30 V116 1.2412599410984492e-11
C30_116 V30 V116 -4.0694238534640563e-20

R30_117 V30 V117 16292.322039925313
L30_117 V30 V117 -4.337728489493857e-12
C30_117 V30 V117 -3.912623855697726e-20

R30_118 V30 V118 -551.8634307577258
L30_118 V30 V118 -2.0738515948253017e-12
C30_118 V30 V118 1.1309630658685369e-19

R30_119 V30 V119 -3068.673617383957
L30_119 V30 V119 -8.004467941984149e-11
C30_119 V30 V119 3.794693932373164e-20

R30_120 V30 V120 -5674.682360921823
L30_120 V30 V120 -2.4548955557223407e-10
C30_120 V30 V120 6.893419889978603e-20

R30_121 V30 V121 -5055.76906060635
L30_121 V30 V121 -3.0216177688426e-12
C30_121 V30 V121 -1.2508933204642965e-19

R30_122 V30 V122 -256390.85048639664
L30_122 V30 V122 3.888775656736078e-12
C30_122 V30 V122 6.565147112050851e-20

R30_123 V30 V123 -2359.1067311167108
L30_123 V30 V123 -4.824024521348472e-12
C30_123 V30 V123 -5.3621972644907527e-20

R30_124 V30 V124 -2012.468287763762
L30_124 V30 V124 -2.373839606665112e-12
C30_124 V30 V124 -1.33205281092268e-19

R30_125 V30 V125 -1415.7454695405063
L30_125 V30 V125 1.6577035500458313e-11
C30_125 V30 V125 6.008325799479666e-20

R30_126 V30 V126 1382.8853896350108
L30_126 V30 V126 5.68792353956355e-12
C30_126 V30 V126 -1.9860827024603739e-19

R30_127 V30 V127 1418.2156474932228
L30_127 V30 V127 3.5884278920849566e-12
C30_127 V30 V127 3.595452552340427e-20

R30_128 V30 V128 1511.8008455543354
L30_128 V30 V128 2.8097931143629954e-12
C30_128 V30 V128 4.965583175047357e-20

R30_129 V30 V129 1162.2490546520803
L30_129 V30 V129 3.1177503893641165e-12
C30_129 V30 V129 1.1167604371748812e-19

R30_130 V30 V130 3312.2753247176656
L30_130 V30 V130 -1.6944620483655792e-12
C30_130 V30 V130 2.1884962275150296e-20

R30_131 V30 V131 -1920.7981466281133
L30_131 V30 V131 -5.155623077628013e-12
C30_131 V30 V131 3.662737623622413e-20

R30_132 V30 V132 -1947.5365852499124
L30_132 V30 V132 -3.6226284699436495e-12
C30_132 V30 V132 6.902077615854799e-20

R30_133 V30 V133 2859.195286520645
L30_133 V30 V133 -2.8101468342718544e-12
C30_133 V30 V133 -9.619044186012663e-20

R30_134 V30 V134 -824.6167381434841
L30_134 V30 V134 1.853924071071212e-12
C30_134 V30 V134 2.48359930344236e-19

R30_135 V30 V135 -2161.952534451893
L30_135 V30 V135 -2.4833650257200604e-12
C30_135 V30 V135 -1.3478892691226547e-19

R30_136 V30 V136 -1331.5650402657084
L30_136 V30 V136 -2.024568282041588e-12
C30_136 V30 V136 -1.41928328043768e-19

R30_137 V30 V137 -607.2407201175107
L30_137 V30 V137 4.27172045051539e-11
C30_137 V30 V137 -6.912516165711451e-20

R30_138 V30 V138 3704.7446083458376
L30_138 V30 V138 -6.329135274573376e-12
C30_138 V30 V138 -2.6130915098077924e-19

R30_139 V30 V139 1112.6856287171129
L30_139 V30 V139 1.6706819293796768e-12
C30_139 V30 V139 1.2079460120502012e-19

R30_140 V30 V140 1232.7455497967953
L30_140 V30 V140 1.0863438401050417e-12
C30_140 V30 V140 1.4458687017930123e-19

R30_141 V30 V141 4104.455062914323
L30_141 V30 V141 1.2313119539796365e-11
C30_141 V30 V141 9.685221290511906e-20

R30_142 V30 V142 401.24178069167107
L30_142 V30 V142 -1.9337663502391857e-12
C30_142 V30 V142 -2.3321042026935182e-20

R30_143 V30 V143 -2592.623602412938
L30_143 V30 V143 -1.0025860528713266e-11
C30_143 V30 V143 4.86234400261493e-20

R30_144 V30 V144 1952.8229954699086
L30_144 V30 V144 -3.9016282371174605e-12
C30_144 V30 V144 3.0118648823977827e-21

R30_145 V30 V145 824.4544242310964
L30_145 V30 V145 -3.020108955421622e-12
C30_145 V30 V145 3.350520449272349e-20

R30_146 V30 V146 -340.4406765662495
L30_146 V30 V146 1.1341667750756188e-11
C30_146 V30 V146 1.1636256730384717e-19

R30_147 V30 V147 3268.871741138192
L30_147 V30 V147 -1.915865901052804e-12
C30_147 V30 V147 -1.7044767170900013e-19

R30_148 V30 V148 -587.2022521060107
L30_148 V30 V148 -1.940479231868306e-12
C30_148 V30 V148 -1.2578034663679727e-19

R30_149 V30 V149 -12304.695542058607
L30_149 V30 V149 -6.885022384028282e-12
C30_149 V30 V149 -1.641598587998696e-19

R30_150 V30 V150 -1040.0198420629008
L30_150 V30 V150 1.994487665103095e-12
C30_150 V30 V150 1.1546670889602646e-19

R30_151 V30 V151 28106.981286621434
L30_151 V30 V151 7.491049537589733e-11
C30_151 V30 V151 3.7666833394822546e-20

R30_152 V30 V152 402.02439372860584
L30_152 V30 V152 3.784189453741855e-12
C30_152 V30 V152 5.822803251109868e-20

R30_153 V30 V153 -650.7221953143872
L30_153 V30 V153 2.2124954660532067e-12
C30_153 V30 V153 1.0358989620052225e-20

R30_154 V30 V154 1336.1637514397967
L30_154 V30 V154 3.432527546843588e-12
C30_154 V30 V154 -1.7921110323982069e-19

R30_155 V30 V155 803.9268678501596
L30_155 V30 V155 2.859783328332309e-12
C30_155 V30 V155 7.17561524715218e-21

R30_156 V30 V156 -344.80286596063297
L30_156 V30 V156 4.779192182506061e-12
C30_156 V30 V156 6.462877160593343e-20

R30_157 V30 V157 10734.058824996488
L30_157 V30 V157 2.6285186393005846e-12
C30_157 V30 V157 1.764094458240774e-19

R30_158 V30 V158 948.7457320337608
L30_158 V30 V158 -1.2151446951672996e-12
C30_158 V30 V158 9.622118758288916e-20

R30_159 V30 V159 -387.8682676750158
L30_159 V30 V159 -2.0416292729790885e-11
C30_159 V30 V159 -4.6495721011931575e-20

R30_160 V30 V160 -1699.0251426155633
L30_160 V30 V160 -1.1098204893777875e-11
C30_160 V30 V160 -1.1239553936141728e-19

R30_161 V30 V161 926.0792994714143
L30_161 V30 V161 1.8087632226047293e-10
C30_161 V30 V161 2.8504686958948296e-20

R30_162 V30 V162 -3361.3340604585637
L30_162 V30 V162 -1.1252231595270117e-11
C30_162 V30 V162 -2.2901141238694338e-21

R30_163 V30 V163 754.1587390928495
L30_163 V30 V163 4.595093869801556e-12
C30_163 V30 V163 1.0170628200129269e-19

R30_164 V30 V164 1050.2504074196254
L30_164 V30 V164 1.7719982476436427e-11
C30_164 V30 V164 7.540050107883857e-20

R30_165 V30 V165 -866.4208205509748
L30_165 V30 V165 -1.1655417960108394e-12
C30_165 V30 V165 -2.0933216143973181e-19

R30_166 V30 V166 -407.001819162698
L30_166 V30 V166 1.0366078565327083e-12
C30_166 V30 V166 -3.103703749271807e-20

R30_167 V30 V167 7786.228020058252
L30_167 V30 V167 -5.4856985967605866e-12
C30_167 V30 V167 3.826417370884827e-20

R30_168 V30 V168 629.5678337638751
L30_168 V30 V168 -7.570184023459979e-12
C30_168 V30 V168 5.109355898431109e-20

R30_169 V30 V169 -1006.39179642033
L30_169 V30 V169 1.1923322010448507e-11
C30_169 V30 V169 -2.935933397456922e-20

R30_170 V30 V170 665.1357479605551
L30_170 V30 V170 -1.3026863674418372e-12
C30_170 V30 V170 -7.076351558512817e-20

R30_171 V30 V171 -1648.1779348259167
L30_171 V30 V171 -3.19081909028789e-12
C30_171 V30 V171 -1.7807015054290294e-19

R30_172 V30 V172 -697.5131158724162
L30_172 V30 V172 -4.077806865220438e-12
C30_172 V30 V172 -1.3221526280360461e-19

R30_173 V30 V173 2297.8861617468333
L30_173 V30 V173 1.5793113939113502e-12
C30_173 V30 V173 1.7131179692834214e-19

R30_174 V30 V174 378.34685122507534
L30_174 V30 V174 -2.084095018223695e-12
C30_174 V30 V174 8.821177864030097e-20

R30_175 V30 V175 27012.681854045946
L30_175 V30 V175 2.471306966201941e-12
C30_175 V30 V175 6.740219194369931e-20

R30_176 V30 V176 -4779.846660732252
L30_176 V30 V176 1.4208262975986293e-12
C30_176 V30 V176 9.618423280390436e-20

R30_177 V30 V177 -2059.2798426464365
L30_177 V30 V177 -4.857170175673057e-12
C30_177 V30 V177 -7.168181589312593e-20

R30_178 V30 V178 -402.39775946099985
L30_178 V30 V178 1.1946733862405213e-12
C30_178 V30 V178 3.434436224059108e-20

R30_179 V30 V179 2392.3783016826446
L30_179 V30 V179 6.30125219816278e-12
C30_179 V30 V179 6.46559177451668e-20

R30_180 V30 V180 8942.116316784817
L30_180 V30 V180 -9.765175753179707e-12
C30_180 V30 V180 1.0802215744301246e-20

R30_181 V30 V181 3392.9731744192545
L30_181 V30 V181 -1.5894112288502585e-11
C30_181 V30 V181 -1.9940141656980725e-20

R30_182 V30 V182 -7700.708111385104
L30_182 V30 V182 -2.5829267740597892e-12
C30_182 V30 V182 -6.931883064121661e-20

R30_183 V30 V183 -1075.7803486105029
L30_183 V30 V183 1.1181273266479539e-10
C30_183 V30 V183 5.271070818370465e-21

R30_184 V30 V184 -2246.3563012215463
L30_184 V30 V184 -7.013425644083521e-12
C30_184 V30 V184 -2.008283264334375e-20

R30_185 V30 V185 -5889.639786329254
L30_185 V30 V185 2.6499346929631125e-11
C30_185 V30 V185 4.7019589930044284e-20

R30_186 V30 V186 636.1647153092738
L30_186 V30 V186 -1.6455386704470189e-12
C30_186 V30 V186 -2.6980149737011454e-20

R30_187 V30 V187 1451.8583866822073
L30_187 V30 V187 -4.6238594147735185e-12
C30_187 V30 V187 -4.5017205357376664e-20

R30_188 V30 V188 664.7352577801865
L30_188 V30 V188 8.713690686605839e-12
C30_188 V30 V188 -3.2582589504093904e-20

R30_189 V30 V189 -1924.9305938092352
L30_189 V30 V189 -7.908460939813009e-11
C30_189 V30 V189 -1.1220305102753877e-19

R30_190 V30 V190 -1088.356766606034
L30_190 V30 V190 3.541577389799424e-12
C30_190 V30 V190 9.438774636018105e-20

R30_191 V30 V191 3903.5729132566935
L30_191 V30 V191 -2.1452684945641335e-11
C30_191 V30 V191 -1.0357103718339706e-19

R30_192 V30 V192 -1653.7913839151674
L30_192 V30 V192 -9.922460902606482e-12
C30_192 V30 V192 -1.0986423520134065e-19

R30_193 V30 V193 1453.7920341333556
L30_193 V30 V193 7.475656531542275e-12
C30_193 V30 V193 5.534812706675139e-20

R30_194 V30 V194 5361.683783029146
L30_194 V30 V194 -4.2318147339220874e-11
C30_194 V30 V194 -5.355279170887147e-20

R30_195 V30 V195 -1259.5318935025664
L30_195 V30 V195 2.495372161143862e-12
C30_195 V30 V195 1.6742318359523993e-19

R30_196 V30 V196 -1151.7029797421408
L30_196 V30 V196 1.34804048573013e-12
C30_196 V30 V196 2.647189572998139e-19

R30_197 V30 V197 4762.683695640929
L30_197 V30 V197 5.783718921291167e-12
C30_197 V30 V197 8.062541696752088e-20

R30_198 V30 V198 1327.0899532845028
L30_198 V30 V198 -6.794613401896129e-12
C30_198 V30 V198 -3.6162174590297935e-20

R30_199 V30 V199 12922.50199580937
L30_199 V30 V199 4.759605241062898e-12
C30_199 V30 V199 1.1538741174779728e-19

R30_200 V30 V200 1110.5539413558888
L30_200 V30 V200 -1.011505293889852e-11
C30_200 V30 V200 -6.158002878509321e-21

R31_31 V31 0 270.33477022754005
L31_31 V31 0 1.024181682207008e-12
C31_31 V31 0 -1.9127462894629667e-19

R31_32 V31 V32 -1441.944679068725
L31_32 V31 V32 -3.7856212371396636e-12
C31_32 V31 V32 -1.0855441251637942e-19

R31_33 V31 V33 11325.6828910429
L31_33 V31 V33 -1.0306564893986477e-11
C31_33 V31 V33 -1.100894742543166e-19

R31_34 V31 V34 4590.634534146386
L31_34 V31 V34 -5.225131941172629e-12
C31_34 V31 V34 -1.2897826631908247e-19

R31_35 V31 V35 1232.8692214027838
L31_35 V31 V35 1.5781960279740362e-12
C31_35 V31 V35 3.274485210156456e-19

R31_36 V31 V36 2072.3199758431488
L31_36 V31 V36 -8.013680626267747e-10
C31_36 V31 V36 -6.390862758468723e-20

R31_37 V31 V37 6350.940529527864
L31_37 V31 V37 3.687351309039893e-12
C31_37 V31 V37 6.237447684942645e-20

R31_38 V31 V38 7739.838310314136
L31_38 V31 V38 2.91286592142771e-12
C31_38 V31 V38 1.6748352229767485e-19

R31_39 V31 V39 681.967331993286
L31_39 V31 V39 2.788065535791061e-12
C31_39 V31 V39 2.8511421441763756e-19

R31_40 V31 V40 1124.8614477272324
L31_40 V31 V40 6.8530785257256895e-12
C31_40 V31 V40 1.0071505579195569e-19

R31_41 V31 V41 -5610.289102716408
L31_41 V31 V41 -9.798388165869332e-11
C31_41 V31 V41 -2.857283492329533e-20

R31_42 V31 V42 -9038.482930062119
L31_42 V31 V42 -1.145915758794973e-11
C31_42 V31 V42 -8.754155977262931e-20

R31_43 V31 V43 5224.656955728266
L31_43 V31 V43 -2.4303848021036103e-12
C31_43 V31 V43 -4.403860893685218e-19

R31_44 V31 V44 -4845.174983011092
L31_44 V31 V44 -1.473459446092029e-11
C31_44 V31 V44 -1.146472529396893e-19

R31_45 V31 V45 -4586.369999913784
L31_45 V31 V45 -8.669424813482222e-10
C31_45 V31 V45 1.3998051005194006e-19

R31_46 V31 V46 -3858.3929303762343
L31_46 V31 V46 -6.12671151093507e-12
C31_46 V31 V46 1.5929378935874363e-20

R31_47 V31 V47 -834.617509623804
L31_47 V31 V47 -6.683680168810448e-12
C31_47 V31 V47 1.0754566383384018e-19

R31_48 V31 V48 -1918.9667165716128
L31_48 V31 V48 -2.518579511396643e-11
C31_48 V31 V48 9.594519109358026e-20

R31_49 V31 V49 31794.85744877332
L31_49 V31 V49 -3.041704944667787e-11
C31_49 V31 V49 1.0320714108715888e-20

R31_50 V31 V50 -18294.181188669594
L31_50 V31 V50 4.008554434571082e-12
C31_50 V31 V50 1.5508170622553085e-19

R31_51 V31 V51 -1444.394063345812
L31_51 V31 V51 2.4722670564762374e-11
C31_51 V31 V51 1.1085182701736372e-20

R31_52 V31 V52 33757.32090453961
L31_52 V31 V52 1.682918819228599e-11
C31_52 V31 V52 3.416039757144168e-20

R31_53 V31 V53 -4957.425767926712
L31_53 V31 V53 -3.2188498925262278e-12
C31_53 V31 V53 -2.0970380648496371e-19

R31_54 V31 V54 153551.20749847067
L31_54 V31 V54 -6.1763322836663696e-12
C31_54 V31 V54 -1.7979871852290053e-19

R31_55 V31 V55 2110.912654647603
L31_55 V31 V55 2.9941404394460153e-12
C31_55 V31 V55 5.710888344371863e-20

R31_56 V31 V56 2925.2832710587436
L31_56 V31 V56 -6.8923402937147144e-12
C31_56 V31 V56 -1.6759587405328383e-19

R31_57 V31 V57 7478.46054584089
L31_57 V31 V57 2.8002614763083025e-12
C31_57 V31 V57 1.3280991929328564e-19

R31_58 V31 V58 -3144.7573035879614
L31_58 V31 V58 1.031744844142274e-08
C31_58 V31 V58 1.0138166356695766e-20

R31_59 V31 V59 1212.2156085683193
L31_59 V31 V59 -7.529743755040759e-12
C31_59 V31 V59 2.8464093735971224e-20

R31_60 V31 V60 2400.613734525112
L31_60 V31 V60 1.1981838013527392e-11
C31_60 V31 V60 8.807431410546462e-20

R31_61 V31 V61 -15935.660047832675
L31_61 V31 V61 -1.697415978617337e-11
C31_61 V31 V61 4.935083554975364e-20

R31_62 V31 V62 2842.8639106656356
L31_62 V31 V62 6.89575890105115e-12
C31_62 V31 V62 1.4056472440589766e-19

R31_63 V31 V63 -13973.024776955113
L31_63 V31 V63 -2.874802798757272e-12
C31_63 V31 V63 -2.6804798270933656e-19

R31_64 V31 V64 -4174.946848610642
L31_64 V31 V64 5.542522969443798e-12
C31_64 V31 V64 1.2744086125097294e-19

R31_65 V31 V65 -9309.913473349347
L31_65 V31 V65 -7.578475242374589e-12
C31_65 V31 V65 -3.915496023959849e-20

R31_66 V31 V66 -7606.899524467445
L31_66 V31 V66 -4.9757738430465687e-11
C31_66 V31 V66 -4.990499581832847e-20

R31_67 V31 V67 -1441.1008722308193
L31_67 V31 V67 4.084646240192542e-12
C31_67 V31 V67 1.1774042042296873e-19

R31_68 V31 V68 -2869.815258204477
L31_68 V31 V68 -6.498123809148333e-12
C31_68 V31 V68 -1.0079786128979721e-19

R31_69 V31 V69 -16755.375698746077
L31_69 V31 V69 9.384104809483439e-11
C31_69 V31 V69 4.760740543343398e-21

R31_70 V31 V70 -5708.47756870374
L31_70 V31 V70 -1.0880266096706232e-11
C31_70 V31 V70 -5.929619495173048e-20

R31_71 V31 V71 -1723.384670593351
L31_71 V31 V71 9.023741896479182e-12
C31_71 V31 V71 2.707352373422445e-19

R31_72 V31 V72 -4119.59483258373
L31_72 V31 V72 -5.491599453338932e-12
C31_72 V31 V72 -5.50496394364789e-20

R31_73 V31 V73 -3224.897893116806
L31_73 V31 V73 -2.6536558625762117e-11
C31_73 V31 V73 -2.80101880206941e-21

R31_74 V31 V74 4920.066762452878
L31_74 V31 V74 1.0455947693484937e-11
C31_74 V31 V74 6.538122782114824e-20

R31_75 V31 V75 1229.5643085944746
L31_75 V31 V75 -3.4617791550470612e-12
C31_75 V31 V75 -3.939052510294142e-19

R31_76 V31 V76 1823.5252760035994
L31_76 V31 V76 3.3428995672858707e-12
C31_76 V31 V76 1.2547154447537646e-19

R31_77 V31 V77 2664.2619762386826
L31_77 V31 V77 8.022546103504848e-12
C31_77 V31 V77 7.69016182083752e-21

R31_78 V31 V78 -5564.49674838064
L31_78 V31 V78 1.27537201103296e-11
C31_78 V31 V78 -2.8475971942985596e-20

R31_79 V31 V79 1437.7935772556257
L31_79 V31 V79 4.884265486637802e-12
C31_79 V31 V79 9.214413465033084e-20

R31_80 V31 V80 3007.2457502820976
L31_80 V31 V80 -3.313390415952686e-11
C31_80 V31 V80 -6.065292374913024e-20

R31_81 V31 V81 -3907.0395088785945
L31_81 V31 V81 -1.561821918637075e-11
C31_81 V31 V81 2.090240198851034e-21

R31_82 V31 V82 7212.852784574745
L31_82 V31 V82 -1.2146957993544361e-11
C31_82 V31 V82 1.6351408571331202e-20

R31_83 V31 V83 -2835.9301298017135
L31_83 V31 V83 4.09888159982343e-12
C31_83 V31 V83 2.125039788550644e-19

R31_84 V31 V84 -3513.940487871361
L31_84 V31 V84 -1.256924589006618e-11
C31_84 V31 V84 1.2137330133286157e-20

R31_85 V31 V85 18178.026222073466
L31_85 V31 V85 -3.198800083162053e-11
C31_85 V31 V85 5.191379740558221e-20

R31_86 V31 V86 -2383.8783875495055
L31_86 V31 V86 -2.1354459272361193e-11
C31_86 V31 V86 6.113598749800652e-20

R31_87 V31 V87 -941.0679287659384
L31_87 V31 V87 -2.4498394235096613e-12
C31_87 V31 V87 -3.428860194346248e-19

R31_88 V31 V88 -5208.058975472532
L31_88 V31 V88 9.727886088500005e-12
C31_88 V31 V88 4.9736257061836744e-20

R31_89 V31 V89 -5258.051540537139
L31_89 V31 V89 -1.6957971347819893e-11
C31_89 V31 V89 -4.682298936809468e-20

R31_90 V31 V90 -51935.27330555942
L31_90 V31 V90 7.271960269638993e-12
C31_90 V31 V90 -1.2905343336472893e-19

R31_91 V31 V91 6002.859639689608
L31_91 V31 V91 2.492438094958151e-12
C31_91 V31 V91 4.0558735428606275e-19

R31_92 V31 V92 -55676.737070275434
L31_92 V31 V92 -3.916051723957731e-12
C31_92 V31 V92 -1.0630840456658269e-19

R31_93 V31 V93 -3579.8850704035094
L31_93 V31 V93 1.1392455848529612e-11
C31_93 V31 V93 -4.4342052686206137e-20

R31_94 V31 V94 2697.7492751101786
L31_94 V31 V94 -1.2469555355784489e-11
C31_94 V31 V94 -5.4352428764486965e-21

R31_95 V31 V95 522.3581975502536
L31_95 V31 V95 4.7023471927453905e-11
C31_95 V31 V95 4.247388468898115e-20

R31_96 V31 V96 1416.3802698238233
L31_96 V31 V96 8.610504616620605e-12
C31_96 V31 V96 3.1060660312705216e-20

R31_97 V31 V97 1408.144015569054
L31_97 V31 V97 1.2976586263262643e-11
C31_97 V31 V97 1.1593990093863088e-19

R31_98 V31 V98 -3161.109668913087
L31_98 V31 V98 -1.658321171868164e-11
C31_98 V31 V98 1.1981255748567052e-19

R31_99 V31 V99 -615.5469120657432
L31_99 V31 V99 -2.2791388252224502e-12
C31_99 V31 V99 -4.7153259985932055e-19

R31_100 V31 V100 -6526.824075388467
L31_100 V31 V100 7.1134145544267115e-12
C31_100 V31 V100 9.774303503139902e-20

R31_101 V31 V101 -3811.482150237378
L31_101 V31 V101 -9.61636897873262e-12
C31_101 V31 V101 -5.0629102000432405e-20

R31_102 V31 V102 11329.498866872196
L31_102 V31 V102 9.300654118370936e-12
C31_102 V31 V102 -5.098813481796925e-20

R31_103 V31 V103 -4138.92710932825
L31_103 V31 V103 1.5697084627134808e-12
C31_103 V31 V103 3.4914239760202353e-19

R31_104 V31 V104 -2195.749801978618
L31_104 V31 V104 -7.31826334028758e-12
C31_104 V31 V104 -7.387921213644412e-20

R31_105 V31 V105 -1183.337346006147
L31_105 V31 V105 -7.301274081519293e-12
C31_105 V31 V105 -6.184269788767997e-20

R31_106 V31 V106 -1374.819035773552
L31_106 V31 V106 -5.128480205986591e-12
C31_106 V31 V106 -1.4198447508962014e-19

R31_107 V31 V107 1351.0235089365165
L31_107 V31 V107 -1.0809531252930423e-11
C31_107 V31 V107 1.9463878468842857e-20

R31_108 V31 V108 11284.43751238105
L31_108 V31 V108 2.808341959650646e-11
C31_108 V31 V108 4.37980306079613e-21

R31_109 V31 V109 2708.6639598210163
L31_109 V31 V109 2.7418323602753968e-11
C31_109 V31 V109 8.189480707657695e-20

R31_110 V31 V110 1456.4039423733534
L31_110 V31 V110 2.2764184467344673e-11
C31_110 V31 V110 1.1396461883069826e-19

R31_111 V31 V111 -556.1419485283818
L31_111 V31 V111 -1.714425972529449e-12
C31_111 V31 V111 -5.886071034869824e-20

R31_112 V31 V112 -2170.3878785012794
L31_112 V31 V112 -5.333749147331696e-12
C31_112 V31 V112 -6.197114643124498e-20

R31_113 V31 V113 2628.328830068431
L31_113 V31 V113 5.6086869573059026e-12
C31_113 V31 V113 2.847390609432391e-20

R31_114 V31 V114 1234.5954788256581
L31_114 V31 V114 5.589804787312341e-12
C31_114 V31 V114 1.0402849432258653e-19

R31_115 V31 V115 557.018052550662
L31_115 V31 V115 3.914760316370719e-12
C31_115 V31 V115 -7.961868713526278e-20

R31_116 V31 V116 1096.905634959202
L31_116 V31 V116 4.614228363767463e-12
C31_116 V31 V116 6.679181588834503e-20

R31_117 V31 V117 3055.1703591077376
L31_117 V31 V117 -8.87621733151808e-12
C31_117 V31 V117 -4.9794728333839944e-20

R31_118 V31 V118 -718.9025397100381
L31_118 V31 V118 -3.6306266438448315e-12
C31_118 V31 V118 -1.4433626040171654e-19

R31_119 V31 V119 -958.2911051243094
L31_119 V31 V119 4.711121105738217e-12
C31_119 V31 V119 -7.2714206287973e-21

R31_120 V31 V120 -1539.4624640450627
L31_120 V31 V120 1.9796544290879255e-11
C31_120 V31 V120 -6.80887010058849e-22

R31_121 V31 V121 -2170.0730641893665
L31_121 V31 V121 -3.6020857496828864e-11
C31_121 V31 V121 9.209896767097538e-21

R31_122 V31 V122 16973.3221109613
L31_122 V31 V122 -3.7640211848282576e-11
C31_122 V31 V122 5.972628156149833e-21

R31_123 V31 V123 -1002.6280363655167
L31_123 V31 V123 -3.610117891433665e-12
C31_123 V31 V123 3.0209623491575953e-19

R31_124 V31 V124 -1485.5087209463388
L31_124 V31 V124 -2.624740518294915e-12
C31_124 V31 V124 -1.2102354014427434e-19

R31_125 V31 V125 -707.0770755911263
L31_125 V31 V125 -2.924315582461399e-11
C31_125 V31 V125 -2.874251876561085e-20

R31_126 V31 V126 2709.8796617749554
L31_126 V31 V126 9.046319450995061e-12
C31_126 V31 V126 9.555854765973024e-20

R31_127 V31 V127 667.9993744213134
L31_127 V31 V127 -4.103511106484809e-12
C31_127 V31 V127 -2.688618056749662e-19

R31_128 V31 V128 976.8369727814536
L31_128 V31 V128 8.255323367812482e-12
C31_128 V31 V128 1.2323573115027975e-19

R31_129 V31 V129 586.5193802543123
L31_129 V31 V129 -8.185594969248623e-12
C31_129 V31 V129 6.931089019430452e-20

R31_130 V31 V130 1774.097113611288
L31_130 V31 V130 9.199907688813314e-11
C31_130 V31 V130 -1.7347156034180714e-20

R31_131 V31 V131 -1336.5813603420977
L31_131 V31 V131 5.801302895796049e-12
C31_131 V31 V131 1.733686644453519e-20

R31_132 V31 V132 -1311.9783519593625
L31_132 V31 V132 9.76962036852402e-12
C31_132 V31 V132 -1.10668088776542e-19

R31_133 V31 V133 1236.46901544902
L31_133 V31 V133 9.070068107100757e-12
C31_133 V31 V133 -1.4869203253583518e-21

R31_134 V31 V134 -2961.7908358021455
L31_134 V31 V134 2.2470322191759323e-11
C31_134 V31 V134 -2.03567451759141e-20

R31_135 V31 V135 -2568.955646860163
L31_135 V31 V135 8.097292212521053e-12
C31_135 V31 V135 4.53794214472375e-19

R31_136 V31 V136 -1667.6531382608332
L31_136 V31 V136 -4.790874711534778e-12
C31_136 V31 V136 -1.4377586684986542e-19

R31_137 V31 V137 -544.5120272078927
L31_137 V31 V137 2.8849439331526177e-12
C31_137 V31 V137 -3.2410423882281263e-20

R31_138 V31 V138 5202.764276403992
L31_138 V31 V138 3.69574864442798e-11
C31_138 V31 V138 6.876894383400574e-20

R31_139 V31 V139 1637.6591797013157
L31_139 V31 V139 1.2085623996220073e-11
C31_139 V31 V139 -6.217357354435639e-19

R31_140 V31 V140 862.9200156350515
L31_140 V31 V140 2.6590546462437138e-12
C31_140 V31 V140 2.086044209885401e-19

R31_141 V31 V141 -1204.95393247752
L31_141 V31 V141 -2.673707494658831e-12
C31_141 V31 V141 2.5856888378009262e-20

R31_142 V31 V142 1852.8407446558986
L31_142 V31 V142 -9.079923339328283e-12
C31_142 V31 V142 -6.323945212642843e-21

R31_143 V31 V143 -1398.5270753362518
L31_143 V31 V143 -2.2830603549375166e-12
C31_143 V31 V143 1.089693482951825e-19

R31_144 V31 V144 -1942.6620230018304
L31_144 V31 V144 -6.631184374094776e-12
C31_144 V31 V144 -4.802190580735264e-20

R31_145 V31 V145 511.73658517433574
L31_145 V31 V145 -2.0184030485389657e-12
C31_145 V31 V145 3.9897890061852566e-20

R31_146 V31 V146 -2538.9893470416814
L31_146 V31 V146 -5.093959219165146e-12
C31_146 V31 V146 -4.274535594520116e-20

R31_147 V31 V147 307.5928369507641
L31_147 V31 V147 -1.1391053245202517e-11
C31_147 V31 V147 3.5134777535288767e-19

R31_148 V31 V148 2325.988315182614
L31_148 V31 V148 -2.172209270260948e-12
C31_148 V31 V148 -9.813607660871166e-20

R31_149 V31 V149 5556.811903647056
L31_149 V31 V149 2.0039417547205423e-12
C31_149 V31 V149 -1.1554927146918673e-19

R31_150 V31 V150 -615.7721681560836
L31_150 V31 V150 5.864816636617916e-12
C31_150 V31 V150 -4.348461273177845e-21

R31_151 V31 V151 -155.65565900984492
L31_151 V31 V151 2.2237797931806224e-12
C31_151 V31 V151 -1.752645147094746e-19

R31_152 V31 V152 -3763.8070426554946
L31_152 V31 V152 5.828416666606321e-12
C31_152 V31 V152 5.689954383492074e-20

R31_153 V31 V153 -1139.7238250658047
L31_153 V31 V153 1.8014591122040925e-12
C31_153 V31 V153 6.68017990118809e-20

R31_154 V31 V154 -100220.16853332763
L31_154 V31 V154 2.493756730161906e-12
C31_154 V31 V154 3.292105506853804e-20

R31_155 V31 V155 93.25458886659611
L31_155 V31 V155 1.0570716136717116e-11
C31_155 V31 V155 -1.951734226815553e-19

R31_156 V31 V156 -1260.0165858540108
L31_156 V31 V156 3.937126713208875e-12
C31_156 V31 V156 8.731471924252893e-20

R31_157 V31 V157 -1419.424512932569
L31_157 V31 V157 -5.230569896520556e-12
C31_157 V31 V157 3.242829417604425e-20

R31_158 V31 V158 -19625.90417221841
L31_158 V31 V158 -4.518071077066424e-12
C31_158 V31 V158 -3.386721690531619e-20

R31_159 V31 V159 -344.56058656929434
L31_159 V31 V159 -1.7795110482616129e-12
C31_159 V31 V159 2.40192088060339e-19

R31_160 V31 V160 5052.3479192592295
L31_160 V31 V160 2.0496385075860247e-11
C31_160 V31 V160 -9.426829166103186e-20

R31_161 V31 V161 2534.969743635009
L31_161 V31 V161 -3.928592091953395e-12
C31_161 V31 V161 -6.871984479136327e-20

R31_162 V31 V162 9557.692165277838
L31_162 V31 V162 -1.0423008628433514e-11
C31_162 V31 V162 -5.1454026309409445e-20

R31_163 V31 V163 -496.48280079953446
L31_163 V31 V163 7.797503905848715e-12
C31_163 V31 V163 -1.1998787063754725e-19

R31_164 V31 V164 -992.459327946893
L31_164 V31 V164 -5.405058619716328e-12
C31_164 V31 V164 1.7009383858903406e-20

R31_165 V31 V165 -5225.698662852371
L31_165 V31 V165 -5.359754461616982e-12
C31_165 V31 V165 2.0067084004213098e-20

R31_166 V31 V166 -2374.90277317507
L31_166 V31 V166 1.5754025959273987e-11
C31_166 V31 V166 9.633987063967151e-21

R31_167 V31 V167 -732.7597954471387
L31_167 V31 V167 1.7606649874798158e-12
C31_167 V31 V167 -3.291768163340615e-20

R31_168 V31 V168 561.5191277533226
L31_168 V31 V168 -9.166224264977732e-12
C31_168 V31 V168 -1.925229443083234e-20

R31_169 V31 V169 -1215.0364568741645
L31_169 V31 V169 3.940268670784382e-12
C31_169 V31 V169 8.647123770857536e-20

R31_170 V31 V170 -1927.1454708555423
L31_170 V31 V170 -7.53277853506789e-11
C31_170 V31 V170 8.298284325934594e-21

R31_171 V31 V171 238.40053499377214
L31_171 V31 V171 -2.5781183107770565e-12
C31_171 V31 V171 9.718280477761244e-20

R31_172 V31 V172 10204.345132512532
L31_172 V31 V172 2.8244588156106145e-11
C31_172 V31 V172 2.732065718071627e-20

R31_173 V31 V173 2622.104029746989
L31_173 V31 V173 1.6956657871662545e-11
C31_173 V31 V173 -6.570464574914835e-20

R31_174 V31 V174 641.6192069014079
L31_174 V31 V174 5.948673005019615e-12
C31_174 V31 V174 1.2240231650306739e-20

R31_175 V31 V175 -484.3285373967143
L31_175 V31 V175 -1.3116493392281244e-11
C31_175 V31 V175 -1.840888770290744e-19

R31_176 V31 V176 25142.877495173907
L31_176 V31 V176 2.779044387161385e-12
C31_176 V31 V176 8.458290769135136e-20

R31_177 V31 V177 -1164.5417741102888
L31_177 V31 V177 -3.341773503360911e-11
C31_177 V31 V177 1.1712627338632872e-20

R31_178 V31 V178 -971.6552770800893
L31_178 V31 V178 -1.0057183132023911e-11
C31_178 V31 V178 9.473885135444311e-21

R31_179 V31 V179 476.9498995874406
L31_179 V31 V179 2.87369642629734e-12
C31_179 V31 V179 1.3188646008317125e-19

R31_180 V31 V180 -1439.8523984499216
L31_180 V31 V180 -4.594257366609391e-12
C31_180 V31 V180 -5.54356344782208e-20

R31_181 V31 V181 1815.7482173613344
L31_181 V31 V181 -1.4818407671942223e-11
C31_181 V31 V181 -9.947811825938502e-21

R31_182 V31 V182 1218.5284686359491
L31_182 V31 V182 -4.608142997970098e-11
C31_182 V31 V182 -4.482085192915887e-20

R31_183 V31 V183 -375.2934888499207
L31_183 V31 V183 -5.9891296211608e-12
C31_183 V31 V183 -1.713518240075803e-20

R31_184 V31 V184 -3423.764045787722
L31_184 V31 V184 -1.4082710417406362e-11
C31_184 V31 V184 4.5249696425338784e-20

R31_185 V31 V185 14423.370526173514
L31_185 V31 V185 -1.1900557342798764e-11
C31_185 V31 V185 -1.8352939727193996e-20

R31_186 V31 V186 1910.771158893191
L31_186 V31 V186 -8.711607987946417e-12
C31_186 V31 V186 5.1254668995582703e-20

R31_187 V31 V187 2269.1434890953396
L31_187 V31 V187 -5.8088030973025045e-12
C31_187 V31 V187 -1.6831524249585416e-19

R31_188 V31 V188 498.57966697523034
L31_188 V31 V188 7.582447897981186e-12
C31_188 V31 V188 -3.029446496726957e-20

R31_189 V31 V189 -1750.4490365515821
L31_189 V31 V189 4.780198278502118e-12
C31_189 V31 V189 3.9848687601125136e-20

R31_190 V31 V190 -1172.6046260243552
L31_190 V31 V190 4.219684641151915e-11
C31_190 V31 V190 -6.642993802509936e-23

R31_191 V31 V191 682.6662223264943
L31_191 V31 V191 3.668139412037244e-12
C31_191 V31 V191 1.9026930138393926e-19

R31_192 V31 V192 -4062.062056971448
L31_192 V31 V192 4.214829648822633e-11
C31_192 V31 V192 -2.8668625951218396e-20

R31_193 V31 V193 3269.7049691213892
L31_193 V31 V193 1.5688902680366897e-10
C31_193 V31 V193 1.0431419528269756e-21

R31_194 V31 V194 3031.391123232132
L31_194 V31 V194 5.76462983672832e-12
C31_194 V31 V194 4.045170699142083e-20

R31_195 V31 V195 -654.9945656175033
L31_195 V31 V195 -4.026755892090485e-12
C31_195 V31 V195 -2.9780412845839637e-19

R31_196 V31 V196 -393.9707490974272
L31_196 V31 V196 4.574293952490232e-12
C31_196 V31 V196 2.082112376175351e-19

R31_197 V31 V197 -3627.3540481318373
L31_197 V31 V197 -1.0296233111666621e-11
C31_197 V31 V197 -1.523579978764132e-20

R31_198 V31 V198 -2767.114954981387
L31_198 V31 V198 -2.2816124686866873e-11
C31_198 V31 V198 -2.0644281285136683e-20

R31_199 V31 V199 30393.22901227689
L31_199 V31 V199 1.0392287413060285e-11
C31_199 V31 V199 -6.485332705809549e-21

R31_200 V31 V200 1108.8475224144731
L31_200 V31 V200 -5.969136048590051e-12
C31_200 V31 V200 -1.0929489660524312e-19

R32_32 V32 0 113.012002052738
L32_32 V32 0 1.3950776204505593e-12
C32_32 V32 0 -1.6033021029549177e-18

R32_33 V32 V33 7969.035136141817
L32_33 V32 V33 -1.0866544117840278e-11
C32_33 V32 V33 -1.3936489354045646e-19

R32_34 V32 V34 2763.5945104550306
L32_34 V32 V34 -4.015719438326895e-12
C32_34 V32 V34 -1.5286104934958532e-19

R32_35 V32 V35 2916.445236009215
L32_35 V32 V35 2.939764133785664e-11
C32_35 V32 V35 -3.8248921056443497e-20

R32_36 V32 V36 833.9639630660567
L32_36 V32 V36 1.5210274491259263e-12
C32_36 V32 V36 1.8672507194960123e-19

R32_37 V32 V37 3558.723394151955
L32_37 V32 V37 2.591234522286792e-12
C32_37 V32 V37 9.570780653192942e-20

R32_38 V32 V38 4785.649560933542
L32_38 V32 V38 2.2303713051976825e-12
C32_38 V32 V38 1.8437691530201046e-19

R32_39 V32 V39 1434.197358961764
L32_39 V32 V39 6.056262572692521e-12
C32_39 V32 V39 1.280528275244913e-19

R32_40 V32 V40 522.3111673605276
L32_40 V32 V40 2.2471384038010407e-12
C32_40 V32 V40 3.800480694986721e-19

R32_41 V32 V41 -4982.561346423485
L32_41 V32 V41 -1.483069343854399e-11
C32_41 V32 V41 -2.3097941213045922e-20

R32_42 V32 V42 -10153.230533247435
L32_42 V32 V42 -8.17594074220446e-12
C32_42 V32 V42 -4.520650248336237e-20

R32_43 V32 V43 -4340.950730715821
L32_43 V32 V43 -1.894707763236919e-11
C32_43 V32 V43 -1.1285670554982577e-19

R32_44 V32 V44 -42275.14359138048
L32_44 V32 V44 -1.8955736019233603e-12
C32_44 V32 V44 -6.013966681064575e-19

R32_45 V32 V45 -2814.436357953815
L32_45 V32 V45 -4.7390409723118494e-11
C32_45 V32 V45 2.0764694924314137e-19

R32_46 V32 V46 -2933.506142584992
L32_46 V32 V46 -4.394321348308827e-12
C32_46 V32 V46 6.890989938685626e-20

R32_47 V32 V47 -2032.7717218974215
L32_47 V32 V47 -2.0146453211813998e-11
C32_47 V32 V47 1.3993104345886838e-19

R32_48 V32 V48 -601.9694384991642
L32_48 V32 V48 -5.138872892388928e-12
C32_48 V32 V48 2.268732515872358e-19

R32_49 V32 V49 43141.01314264404
L32_49 V32 V49 1.2794575376863528e-10
C32_49 V32 V49 6.601332902626988e-20

R32_50 V32 V50 28291.82453125327
L32_50 V32 V50 2.6837005933751383e-12
C32_50 V32 V50 2.2867421327727333e-19

R32_51 V32 V51 -6480.103714087525
L32_51 V32 V51 1.1628372861129796e-11
C32_51 V32 V51 1.1740136525974898e-19

R32_52 V32 V52 -3445.186974849593
L32_52 V32 V52 1.0011976477703566e-11
C32_52 V32 V52 -3.5783618601603736e-20

R32_53 V32 V53 -4553.64312291446
L32_53 V32 V53 -2.5356062322708693e-12
C32_53 V32 V53 -3.0371815689486463e-19

R32_54 V32 V54 9196.232642153927
L32_54 V32 V54 -5.217256759931725e-12
C32_54 V32 V54 -2.65782121327602e-19

R32_55 V32 V55 23343.34673975256
L32_55 V32 V55 -5.924501271646625e-12
C32_55 V32 V55 -1.9872454262525794e-19

R32_56 V32 V56 926.6292293540622
L32_56 V32 V56 2.6334293143444597e-12
C32_56 V32 V56 -1.4648302145288075e-19

R32_57 V32 V57 4934.068105776189
L32_57 V32 V57 2.302170065380323e-12
C32_57 V32 V57 2.234803353675372e-19

R32_58 V32 V58 -2554.5789757306206
L32_58 V32 V58 -2.01552184549806e-11
C32_58 V32 V58 5.3186764925584957e-20

R32_59 V32 V59 2981.2593034716906
L32_59 V32 V59 1.8953897367376518e-11
C32_59 V32 V59 1.4519256082985255e-19

R32_60 V32 V60 971.0248630866716
L32_60 V32 V60 -7.983803708897182e-12
C32_60 V32 V60 3.0533967291029567e-20

R32_61 V32 V61 -8879.165995347135
L32_61 V32 V61 -1.518054635059036e-11
C32_61 V32 V61 7.080636784101543e-20

R32_62 V32 V62 2596.7601770828983
L32_62 V32 V62 5.067377561470887e-12
C32_62 V32 V62 2.3352643536306984e-19

R32_63 V32 V63 -7892.653903338258
L32_63 V32 V63 4.366374604606492e-12
C32_63 V32 V63 9.122221672253397e-20

R32_64 V32 V64 -2172.8954556282138
L32_64 V32 V64 -3.670400772632707e-12
C32_64 V32 V64 -1.42002314137482e-19

R32_65 V32 V65 -5525.944501602756
L32_65 V32 V65 -4.9848972585377365e-12
C32_65 V32 V65 -2.659003049273561e-20

R32_66 V32 V66 -16890.6105729938
L32_66 V32 V66 -1.1433231166250752e-10
C32_66 V32 V66 -4.7657096481052556e-20

R32_67 V32 V67 -26137.473894608855
L32_67 V32 V67 -8.705009797811598e-12
C32_67 V32 V67 -1.2225265781800931e-19

R32_68 V32 V68 -1099.4235024300049
L32_68 V32 V68 6.718792373354507e-11
C32_68 V32 V68 5.386728617505454e-20

R32_69 V32 V69 1501584.5335309508
L32_69 V32 V69 1.5758699749530475e-11
C32_69 V32 V69 -4.070602921477558e-20

R32_70 V32 V70 -4641.010123738477
L32_70 V32 V70 -9.053216445084257e-12
C32_70 V32 V70 -1.496116015072302e-19

R32_71 V32 V71 -4902.207072757354
L32_71 V32 V71 -5.688878883005712e-12
C32_71 V32 V71 -9.548240355477492e-22

R32_72 V32 V72 -1488.313887458259
L32_72 V32 V72 8.526032548318157e-12
C32_72 V32 V72 2.2951028393895984e-19

R32_73 V32 V73 -3079.6081455451176
L32_73 V32 V73 -2.618524486518128e-11
C32_73 V32 V73 5.1659990923438814e-20

R32_74 V32 V74 3802.183752840284
L32_74 V32 V74 6.93875447545099e-12
C32_74 V32 V74 1.506585056014823e-19

R32_75 V32 V75 -14348.241168175517
L32_75 V32 V75 5.3899936339553285e-12
C32_75 V32 V75 1.3803819593532485e-19

R32_76 V32 V76 582.6860093679387
L32_76 V32 V76 -1.6387056027852778e-10
C32_76 V32 V76 -4.543847312513219e-19

R32_77 V32 V77 2589.7574731652035
L32_77 V32 V77 6.8436191690189795e-12
C32_77 V32 V77 4.921495177411151e-20

R32_78 V32 V78 -2946.4565364506398
L32_78 V32 V78 1.0926698531306324e-11
C32_78 V32 V78 -8.506047001838496e-20

R32_79 V32 V79 1786.72815376528
L32_79 V32 V79 2.589555149628718e-11
C32_79 V32 V79 -6.818128032611004e-20

R32_80 V32 V80 11184.211345168196
L32_80 V32 V80 1.6580953517473845e-11
C32_80 V32 V80 1.2070796392497464e-19

R32_81 V32 V81 -1893.5271402168196
L32_81 V32 V81 -8.795836143356564e-12
C32_81 V32 V81 2.8756677320527866e-20

R32_82 V32 V82 5321.1082692218715
L32_82 V32 V82 -7.71180270429487e-12
C32_82 V32 V82 5.677917557499644e-20

R32_83 V32 V83 -4334.188748168344
L32_83 V32 V83 -1.9032961127891614e-11
C32_83 V32 V83 3.581468266490844e-20

R32_84 V32 V84 -2002.6509967549464
L32_84 V32 V84 5.1934082195935766e-12
C32_84 V32 V84 2.9928568185831734e-19

R32_85 V32 V85 10687.954965865196
L32_85 V32 V85 -2.5746267779840835e-11
C32_85 V32 V85 6.56275030859109e-20

R32_86 V32 V86 -3220.157847735245
L32_86 V32 V86 -2.173834682498634e-11
C32_86 V32 V86 1.3121233775686459e-19

R32_87 V32 V87 -3764.025562790109
L32_87 V32 V87 1.7934025236036537e-11
C32_87 V32 V87 -1.5080357013413065e-20

R32_88 V32 V88 -1025.1556789071597
L32_88 V32 V88 -2.5553201635451376e-12
C32_88 V32 V88 -4.858567822551679e-19

R32_89 V32 V89 -10700.894280068676
L32_89 V32 V89 -1.646088811202207e-11
C32_89 V32 V89 -1.1426250772174554e-19

R32_90 V32 V90 248865.50471456387
L32_90 V32 V90 4.598363183336701e-12
C32_90 V32 V90 -2.0541169540636873e-19

R32_91 V32 V91 -2488.3940538967236
L32_91 V32 V91 -3.7982218945774646e-12
C32_91 V32 V91 4.175430943544393e-20

R32_92 V32 V92 1828.741377909379
L32_92 V32 V92 2.2504705301693304e-12
C32_92 V32 V92 4.478135001509703e-19

R32_93 V32 V93 -2061.668021630851
L32_93 V32 V93 1.1468264165405794e-11
C32_93 V32 V93 -3.3126886135166424e-20

R32_94 V32 V94 3340.589093559297
L32_94 V32 V94 -5.98810304438894e-12
C32_94 V32 V94 3.263299621807065e-20

R32_95 V32 V95 1562.6213554474634
L32_95 V32 V95 1.3932963985573077e-11
C32_95 V32 V95 2.24811993840311e-20

R32_96 V32 V96 412.96469578117075
L32_96 V32 V96 1.447960625414263e-11
C32_96 V32 V96 7.709493913029546e-20

R32_97 V32 V97 1239.2474523886103
L32_97 V32 V97 1.4720841874984042e-11
C32_97 V32 V97 3.06250403584434e-19

R32_98 V32 V98 -3209.7525911494045
L32_98 V32 V98 -2.0982362991887128e-11
C32_98 V32 V98 2.300626719674614e-19

R32_99 V32 V99 23114.31128043549
L32_99 V32 V99 5.3687763634804045e-12
C32_99 V32 V99 -1.5778865420966207e-20

R32_100 V32 V100 -384.45275695365007
L32_100 V32 V100 -1.5863772231350484e-12
C32_100 V32 V100 -6.097057091828053e-19

R32_101 V32 V101 -3454.0710348522725
L32_101 V32 V101 -5.871643431757482e-12
C32_101 V32 V101 -1.054222068226501e-19

R32_102 V32 V102 7875.534207536134
L32_102 V32 V102 6.215101074446004e-12
C32_102 V32 V102 -1.1030293636868211e-19

R32_103 V32 V103 -1913.6348302947122
L32_103 V32 V103 -7.808625462495978e-12
C32_103 V32 V103 -1.996105016797319e-20

R32_104 V32 V104 -4960.4169322184025
L32_104 V32 V104 1.767389989593198e-12
C32_104 V32 V104 4.631530700128903e-19

R32_105 V32 V105 -925.2100531608543
L32_105 V32 V105 -6.4097133502521266e-12
C32_105 V32 V105 -1.0183925335268954e-19

R32_106 V32 V106 -1137.2779509831703
L32_106 V32 V106 -3.9830431504375714e-12
C32_106 V32 V106 -1.9376091093605329e-19

R32_107 V32 V107 -36080.85621825199
L32_107 V32 V107 -1.681839617720662e-11
C32_107 V32 V107 7.39932390081524e-20

R32_108 V32 V108 689.8372324245695
L32_108 V32 V108 7.464024993729647e-11
C32_108 V32 V108 -1.2056760661573211e-19

R32_109 V32 V109 1185.2492733785223
L32_109 V32 V109 1.211739756752822e-11
C32_109 V32 V109 2.0676676847030775e-19

R32_110 V32 V110 1037.540042786803
L32_110 V32 V110 1.0821187428038322e-11
C32_110 V32 V110 9.444041796551322e-20

R32_111 V32 V111 -1847.602008658299
L32_111 V32 V111 -4.218312809442246e-12
C32_111 V32 V111 -6.309916123201632e-20

R32_112 V32 V112 -638.2999013775252
L32_112 V32 V112 -2.2890295994416654e-12
C32_112 V32 V112 1.9954526731691723e-19

R32_113 V32 V113 7076.496792998595
L32_113 V32 V113 4.99366482825305e-12
C32_113 V32 V113 2.930281953348055e-20

R32_114 V32 V114 1214.73116164826
L32_114 V32 V114 4.758774532557379e-12
C32_114 V32 V114 1.7272236353832534e-19

R32_115 V32 V115 666.0716694982408
L32_115 V32 V115 2.594529979282605e-12
C32_115 V32 V115 7.848179103581478e-21

R32_116 V32 V116 745.1026215662914
L32_116 V32 V116 5.5414453238496625e-12
C32_116 V32 V116 -9.642938187743792e-20

R32_117 V32 V117 3950.585536704915
L32_117 V32 V117 -7.402211541081746e-12
C32_117 V32 V117 -9.862069159079651e-20

R32_118 V32 V118 -573.592924847798
L32_118 V32 V118 -2.973213049899202e-12
C32_118 V32 V118 -1.8785274287176745e-19

R32_119 V32 V119 -1225.8939129543853
L32_119 V32 V119 -2.282811982503041e-11
C32_119 V32 V119 -1.4328015179320908e-19

R32_120 V32 V120 -571.9116745509541
L32_120 V32 V120 3.768499608986354e-12
C32_120 V32 V120 -3.545885721900185e-19

R32_121 V32 V121 -5603.502865167154
L32_121 V32 V121 -5.4553040624696866e-11
C32_121 V32 V121 2.3969794998470666e-20

R32_122 V32 V122 3720.4804467325666
L32_122 V32 V122 1.1898160101544798e-10
C32_122 V32 V122 -7.623092148384005e-20

R32_123 V32 V123 -1283.6371622059974
L32_123 V32 V123 -2.9178181708264024e-12
C32_123 V32 V123 3.3295043252072096e-20

R32_124 V32 V124 5727.2361653215075
L32_124 V32 V124 -2.8888982294544077e-12
C32_124 V32 V124 7.295246699635813e-19

R32_125 V32 V125 -589.3490064659702
L32_125 V32 V125 -6.615018852609537e-11
C32_125 V32 V125 -8.86018091229796e-21

R32_126 V32 V126 2440.162545956573
L32_126 V32 V126 6.2398913014669066e-12
C32_126 V32 V126 1.2599776097779417e-19

R32_127 V32 V127 724.28608455059
L32_127 V32 V127 2.9145267706451843e-12
C32_127 V32 V127 2.2093637193109185e-19

R32_128 V32 V128 572.2863191985737
L32_128 V32 V128 -3.4563922681465163e-12
C32_128 V32 V128 -1.987940611177557e-19

R32_129 V32 V129 495.53003817110067
L32_129 V32 V129 -5.213312101491148e-12
C32_129 V32 V129 1.1363271661066708e-19

R32_130 V32 V130 2056.305466516466
L32_130 V32 V130 -3.749663386895157e-11
C32_130 V32 V130 -5.624155570921003e-20

R32_131 V32 V131 -772.3173439607566
L32_131 V32 V131 -6.711751574329972e-12
C32_131 V32 V131 -2.243605769807803e-19

R32_132 V32 V132 -523.0383670430838
L32_132 V32 V132 3.2762506500087022e-12
C32_132 V32 V132 -2.3002540525504085e-19

R32_133 V32 V133 1732.8876431109877
L32_133 V32 V133 7.0720672201580795e-12
C32_133 V32 V133 -1.2195424767510428e-19

R32_134 V32 V134 -1233.758506658109
L32_134 V32 V134 3.5849272129178105e-11
C32_134 V32 V134 -2.1097898791344638e-19

R32_135 V32 V135 -10269.503442776448
L32_135 V32 V135 -4.661371911964849e-12
C32_135 V32 V135 -1.4114693017861248e-19

R32_136 V32 V136 -2959.3627638354733
L32_136 V32 V136 -1.1778983637179502e-11
C32_136 V32 V136 5.581123202346574e-19

R32_137 V32 V137 -559.6780778354755
L32_137 V32 V137 2.1925780965901604e-12
C32_137 V32 V137 6.217676482098462e-20

R32_138 V32 V138 1584.341396365804
L32_138 V32 V138 1.8464221591147756e-11
C32_138 V32 V138 2.0214729358879938e-19

R32_139 V32 V139 600.2617891031789
L32_139 V32 V139 1.964846496417782e-12
C32_139 V32 V139 2.0710669326388402e-19

R32_140 V32 V140 -20659.18907984661
L32_140 V32 V140 2.1319981435970166e-12
C32_140 V32 V140 -6.375532850628268e-19

R32_141 V32 V141 -1539.4997017262363
L32_141 V32 V141 -2.0423251198238687e-12
C32_141 V32 V141 4.379552672934016e-20

R32_142 V32 V142 1067.9691170034125
L32_142 V32 V142 -4.394122486209311e-11
C32_142 V32 V142 3.077966268930879e-20

R32_143 V32 V143 -784.115395631751
L32_143 V32 V143 -4.269553811756107e-12
C32_143 V32 V143 -1.375045523343442e-20

R32_144 V32 V144 343.35977931365784
L32_144 V32 V144 -2.485311269858438e-12
C32_144 V32 V144 1.0582159937316572e-19

R32_145 V32 V145 524.6301094366816
L32_145 V32 V145 -1.7377624720185025e-12
C32_145 V32 V145 -2.833391345580224e-20

R32_146 V32 V146 -3163.949959699497
L32_146 V32 V146 -2.7322098711268343e-12
C32_146 V32 V146 -9.726171980840317e-20

R32_147 V32 V147 733.6172380931793
L32_147 V32 V147 -2.3634580375503407e-12
C32_147 V32 V147 1.81856450498652e-20

R32_148 V32 V148 -204.55813444171702
L32_148 V32 V148 -4.348094525614203e-12
C32_148 V32 V148 3.320769961398033e-19

R32_149 V32 V149 2743.827372638562
L32_149 V32 V149 1.60582231080888e-12
C32_149 V32 V149 -2.9602091954741787e-20

R32_150 V32 V150 -471.8487941320213
L32_150 V32 V150 4.852398329303536e-12
C32_150 V32 V150 8.892101042119286e-20

R32_151 V32 V151 -933.0569914793505
L32_151 V32 V151 1.4485262723033872e-11
C32_151 V32 V151 1.2588862000275282e-20

R32_152 V32 V152 841.3040182787581
L32_152 V32 V152 3.0835260799044117e-12
C32_152 V32 V152 -1.0469516590146973e-19

R32_153 V32 V153 -1776.5432894767077
L32_153 V32 V153 1.6242357696126962e-12
C32_153 V32 V153 3.119996302680021e-20

R32_154 V32 V154 747.3934358287364
L32_154 V32 V154 2.2695583630233914e-12
C32_154 V32 V154 3.220447060353028e-20

R32_155 V32 V155 308.60927206944467
L32_155 V32 V155 2.050444699769593e-12
C32_155 V32 V155 -3.109641370614704e-21

R32_156 V32 V156 -479.6446125072426
L32_156 V32 V156 2.4774954601947923e-12
C32_156 V32 V156 -2.8607470040519573e-19

R32_157 V32 V157 -594.281488921513
L32_157 V32 V157 -5.580606678125491e-12
C32_157 V32 V157 1.7769465295326044e-19

R32_158 V32 V158 -905.5151057574678
L32_158 V32 V158 -4.4091684293655e-12
C32_158 V32 V158 -2.8230324001857625e-20

R32_159 V32 V159 -315.3292759639948
L32_159 V32 V159 -1.3349229986809102e-11
C32_159 V32 V159 -3.657659460198373e-20

R32_160 V32 V160 249.89712958876
L32_160 V32 V160 -1.4958892740864578e-12
C32_160 V32 V160 1.757062574499435e-19

R32_161 V32 V161 1092.314414577354
L32_161 V32 V161 -2.862457776894716e-12
C32_161 V32 V161 -1.4646808674645415e-19

R32_162 V32 V162 4359.586183551149
L32_162 V32 V162 -8.176990121819329e-12
C32_162 V32 V162 -2.775485826282137e-20

R32_163 V32 V163 -13484.970244406606
L32_163 V32 V163 -9.114777973502374e-12
C32_163 V32 V163 4.5039639730314473e-20

R32_164 V32 V164 -188.8611343960624
L32_164 V32 V164 -1.3976894847069427e-11
C32_164 V32 V164 -1.097399694802554e-19

R32_165 V32 V165 -822.8989067318391
L32_165 V32 V165 -3.881773235548022e-12
C32_165 V32 V165 4.8728881535826064e-20

R32_166 V32 V166 -1232.0705220867221
L32_166 V32 V166 1.5110252612577233e-11
C32_166 V32 V166 8.717976060138936e-20

R32_167 V32 V167 -776.407869722949
L32_167 V32 V167 -5.301434987017545e-12
C32_167 V32 V167 -4.4214225317117466e-20

R32_168 V32 V168 248.31212589834468
L32_168 V32 V168 1.571819462716091e-12
C32_168 V32 V168 -4.7995911978681947e-20

R32_169 V32 V169 -1937.2432830473135
L32_169 V32 V169 3.5391902859556814e-12
C32_169 V32 V169 2.0345916356148594e-19

R32_170 V32 V170 -4567.15187534523
L32_170 V32 V170 -8.783769802436009e-11
C32_170 V32 V170 -2.356269443284723e-21

R32_171 V32 V171 631.9883591572344
L32_171 V32 V171 1.0919724003850159e-11
C32_171 V32 V171 2.7250811780875516e-20

R32_172 V32 V172 1726.8748979315874
L32_172 V32 V172 -3.3468929699783054e-12
C32_172 V32 V172 7.701142339921741e-20

R32_173 V32 V173 2520.152372476144
L32_173 V32 V173 8.047603252723741e-12
C32_173 V32 V173 -1.2710644972574403e-19

R32_174 V32 V174 557.4340401259938
L32_174 V32 V174 4.384950011313621e-12
C32_174 V32 V174 2.5167983827068823e-20

R32_175 V32 V175 -2852.2536188555223
L32_175 V32 V175 2.892563435432581e-12
C32_175 V32 V175 2.418517600743959e-20

R32_176 V32 V176 -577.78104550064
L32_176 V32 V176 5.538129544029343e-12
C32_176 V32 V176 -2.1994912959399126e-19

R32_177 V32 V177 -972.4013380048864
L32_177 V32 V177 -9.358467172303424e-12
C32_177 V32 V177 3.4672364142411243e-20

R32_178 V32 V178 -808.9301361319942
L32_178 V32 V178 -6.7561007506786265e-12
C32_178 V32 V178 6.879847405629613e-21

R32_179 V32 V179 9998.422449489346
L32_179 V32 V179 -5.243992636321154e-12
C32_179 V32 V179 2.1510555241928012e-20

R32_180 V32 V180 1927.6843682263122
L32_180 V32 V180 4.210829245990872e-12
C32_180 V32 V180 1.7724058471186902e-19

R32_181 V32 V181 1496.1394488031935
L32_181 V32 V181 -2.206707498362768e-11
C32_181 V32 V181 -1.9104230986202936e-20

R32_182 V32 V182 999.7483333253203
L32_182 V32 V182 4.141069998133097e-11
C32_182 V32 V182 -3.7056919557473055e-21

R32_183 V32 V183 -1183.711103916584
L32_183 V32 V183 -2.8784996342882764e-11
C32_183 V32 V183 5.2603193609719824e-20

R32_184 V32 V184 -878.0614721138627
L32_184 V32 V184 -4.367898803528606e-12
C32_184 V32 V184 -2.0869943017933833e-20

R32_185 V32 V185 -5788.040366006111
L32_185 V32 V185 -1.0550338744277135e-11
C32_185 V32 V185 -2.3588118659403152e-20

R32_186 V32 V186 17163.95014841589
L32_186 V32 V186 -7.132831968687182e-12
C32_186 V32 V186 -4.72497202759101e-21

R32_187 V32 V187 1971.9661033932884
L32_187 V32 V187 7.969361483088734e-12
C32_187 V32 V187 -6.174109410398084e-20

R32_188 V32 V188 316.35816715858596
L32_188 V32 V188 -6.616655413029912e-12
C32_188 V32 V188 -2.0988680300698263e-19

R32_189 V32 V189 -4563.8787940483835
L32_189 V32 V189 3.886154849032031e-12
C32_189 V32 V189 6.517152125770721e-20

R32_190 V32 V190 -931.2530376533043
L32_190 V32 V190 1.1319396786580796e-10
C32_190 V32 V190 3.176868670831712e-20

R32_191 V32 V191 1220.8819292690825
L32_191 V32 V191 2.441213541886268e-11
C32_191 V32 V191 -5.1703205694890654e-20

R32_192 V32 V192 -11459.481458140546
L32_192 V32 V192 3.083465185862405e-12
C32_192 V32 V192 3.120811550230671e-19

R32_193 V32 V193 1168.8462594127807
L32_193 V32 V193 7.270299739967665e-11
C32_193 V32 V193 4.5667353940823126e-20

R32_194 V32 V194 51802.17688654049
L32_194 V32 V194 4.303941948601198e-12
C32_194 V32 V194 2.1189140004803595e-19

R32_195 V32 V195 -721.8485793419322
L32_195 V32 V195 2.1823165283188665e-10
C32_195 V32 V195 2.5145537801763533e-19

R32_196 V32 V196 -351.61525690120703
L32_196 V32 V196 -5.309953170394656e-12
C32_196 V32 V196 -4.596738244528342e-19

R32_197 V32 V197 -51239.24987937271
L32_197 V32 V197 -8.421170765442729e-12
C32_197 V32 V197 -7.707377947813255e-20

R32_198 V32 V198 -1610.6951549905266
L32_198 V32 V198 -3.735502978762739e-11
C32_198 V32 V198 8.019602378416156e-20

R32_199 V32 V199 -430.2143506431471
L32_199 V32 V199 -4.995123934496243e-11
C32_199 V32 V199 1.53990946564166e-20

R32_200 V32 V200 358.0579816270706
L32_200 V32 V200 -6.215832909351739e-11
C32_200 V32 V200 -2.3688230143884618e-20

R33_33 V33 0 140.7363441652566
L33_33 V33 0 2.658230567797815e-12
C33_33 V33 0 -9.108946247006527e-19

R33_34 V33 V34 -5867.9391804808
L33_34 V33 V34 -2.5232602538432657e-12
C33_34 V33 V34 -4.6715745057871994e-20

R33_35 V33 V35 -17678.94451419416
L33_35 V33 V35 -2.0861976175239396e-12
C33_35 V33 V35 -1.6385805368663384e-19

R33_36 V33 V36 -11229.64580086417
L33_36 V33 V36 -1.5231477396961206e-12
C33_36 V33 V36 -2.693002307806295e-19

R33_37 V33 V37 1792.1211958037268
L33_37 V33 V37 1.5362219773975548e-12
C33_37 V33 V37 2.9823887115408187e-19

R33_38 V33 V38 144897.20599418395
L33_38 V33 V38 1.631681144113115e-11
C33_38 V33 V38 3.4296847941120045e-20

R33_39 V33 V39 -17953.331945445494
L33_39 V33 V39 2.6678566470320957e-12
C33_39 V33 V39 2.228223351645847e-19

R33_40 V33 V40 -10192.004366040646
L33_40 V33 V40 1.9494204904884338e-12
C33_40 V33 V40 2.910671530512129e-19

R33_41 V33 V41 8496.749654600842
L33_41 V33 V41 3.931118840899567e-12
C33_41 V33 V41 1.5855829176816105e-19

R33_42 V33 V42 7463.0612658058235
L33_42 V33 V42 3.587171801644179e-11
C33_42 V33 V42 1.429437399349184e-20

R33_43 V33 V43 4805.152553145796
L33_43 V33 V43 -1.522036385642472e-11
C33_43 V33 V43 -6.554337820026418e-20

R33_44 V33 V44 3695.487357027809
L33_44 V33 V44 2.9927184339339885e-09
C33_44 V33 V44 -6.386685067685527e-20

R33_45 V33 V45 -2768.146102642017
L33_45 V33 V45 3.656390606325322e-11
C33_45 V33 V45 -1.0417325738205958e-19

R33_46 V33 V46 4158.220766360779
L33_46 V33 V46 2.0803180188570036e-12
C33_46 V33 V46 1.2062400529205994e-19

R33_47 V33 V47 4781.967515246909
L33_47 V33 V47 6.84567010652865e-12
C33_47 V33 V47 -2.0024007085814463e-20

R33_48 V33 V48 3602.5857008305743
L33_48 V33 V48 3.5400142192284862e-12
C33_48 V33 V48 1.9777743103959853e-20

R33_49 V33 V49 -1617.7795517419984
L33_49 V33 V49 2.30232296160549e-11
C33_49 V33 V49 1.4414138455562443e-19

R33_50 V33 V50 56715.92653623384
L33_50 V33 V50 -2.7714280021577544e-12
C33_50 V33 V50 -7.771321159665745e-20

R33_51 V33 V51 32965.15110339827
L33_51 V33 V51 -9.751944677489834e-12
C33_51 V33 V51 1.2618172541493874e-21

R33_52 V33 V52 20273.7782282821
L33_52 V33 V52 -8.399833908558897e-12
C33_52 V33 V52 -2.6254987797803364e-20

R33_53 V33 V53 -1722.109136600581
L33_53 V33 V53 -1.3852991757600763e-12
C33_53 V33 V53 -2.186821545549735e-19

R33_54 V33 V54 -3952.6867510447787
L33_54 V33 V54 -3.1589816849906156e-12
C33_54 V33 V54 -8.04600927849687e-20

R33_55 V33 V55 -4218.529755585652
L33_55 V33 V55 -4.469493467332504e-12
C33_55 V33 V55 -5.940659193200908e-20

R33_56 V33 V56 -2841.3393981449713
L33_56 V33 V56 -2.4227348550048717e-12
C33_56 V33 V56 -1.2509333638023232e-19

R33_57 V33 V57 -2886.469774245972
L33_57 V33 V57 9.454040426746412e-12
C33_57 V33 V57 1.707810353834884e-19

R33_58 V33 V58 3908.6714007897426
L33_58 V33 V58 9.996217838478982e-12
C33_58 V33 V58 1.363257030197528e-20

R33_59 V33 V59 4169.246358618348
L33_59 V33 V59 3.0623180158620686e-12
C33_59 V33 V59 1.2055998659643772e-19

R33_60 V33 V60 3231.4300248402023
L33_60 V33 V60 2.2670689163205596e-12
C33_60 V33 V60 1.5602755088466126e-19

R33_61 V33 V61 3162.705988035672
L33_61 V33 V61 4.852806273035116e-12
C33_61 V33 V61 9.191077498342055e-21

R33_62 V33 V62 -33844.53469941722
L33_62 V33 V62 3.996710406712701e-12
C33_62 V33 V62 1.0819675650691089e-19

R33_63 V33 V63 30767.30471209796
L33_63 V33 V63 -2.87077347097059e-11
C33_63 V33 V63 -5.1384063176752284e-20

R33_64 V33 V64 13113.354173387028
L33_64 V33 V64 9.553141404401389e-12
C33_64 V33 V64 -4.301693627400727e-20

R33_65 V33 V65 -4305.291595352819
L33_65 V33 V65 -2.0236219834977534e-11
C33_65 V33 V65 -1.6139327883285204e-20

R33_66 V33 V66 11160.363668142905
L33_66 V33 V66 -1.6262862457896748e-11
C33_66 V33 V66 2.470969997922216e-20

R33_67 V33 V67 15531.9849892422
L33_67 V33 V67 -3.693493811291942e-12
C33_67 V33 V67 -8.862661248499515e-20

R33_68 V33 V68 6716.6216685517065
L33_68 V33 V68 -5.366636173027042e-12
C33_68 V33 V68 -7.713168045258158e-20

R33_69 V33 V69 -1387.9966423724259
L33_69 V33 V69 -1.129580442306491e-11
C33_69 V33 V69 3.198194610240715e-20

R33_70 V33 V70 13770.587253510343
L33_70 V33 V70 -5.0979516863150115e-12
C33_70 V33 V70 -1.11108982692395e-19

R33_71 V33 V71 7208.793204518572
L33_71 V33 V71 3.4565968948648376e-12
C33_71 V33 V71 1.1072720777499424e-19

R33_72 V33 V72 8213.313768697382
L33_72 V33 V72 6.427741899953101e-12
C33_72 V33 V72 8.32240208559979e-20

R33_73 V33 V73 86607.20299089365
L33_73 V33 V73 -4.07725030632668e-12
C33_73 V33 V73 -1.0995654868996741e-19

R33_74 V33 V74 -15068.808581314614
L33_74 V33 V74 1.1442157212185053e-11
C33_74 V33 V74 2.8715636991117534e-20

R33_75 V33 V75 420618.47366482037
L33_75 V33 V75 1.1857956699145167e-11
C33_75 V33 V75 1.4524717355500686e-21

R33_76 V33 V76 -6326.3101544468
L33_76 V33 V76 -6.631679012498485e-12
C33_76 V33 V76 -7.34059771274461e-20

R33_77 V33 V77 8705.219193294652
L33_77 V33 V77 3.9639072124542606e-11
C33_77 V33 V77 9.163925023137763e-20

R33_78 V33 V78 -6210.399275354819
L33_78 V33 V78 -6.971230690689603e-12
C33_78 V33 V78 -7.251157365408195e-20

R33_79 V33 V79 -2970.82455631023
L33_79 V33 V79 -5.6944268730294335e-12
C33_79 V33 V79 -6.84238942630956e-21

R33_80 V33 V80 -3978.9911897619772
L33_80 V33 V80 1.231662943337059e-11
C33_80 V33 V80 5.648517392086041e-20

R33_81 V33 V81 -800.94680605867
L33_81 V33 V81 4.331395117001464e-12
C33_81 V33 V81 1.6867250256362445e-19

R33_82 V33 V82 4603.198217029296
L33_82 V33 V82 3.970210112378494e-12
C33_82 V33 V82 1.6632163728577563e-19

R33_83 V33 V83 2244.2744840416253
L33_83 V33 V83 2.3163626507869913e-11
C33_83 V33 V83 -2.0603481896195218e-20

R33_84 V33 V84 1868.9338651382018
L33_84 V33 V84 3.0278891790819076e-12
C33_84 V33 V84 3.825010098726672e-20

R33_85 V33 V85 7426.973063262408
L33_85 V33 V85 -7.881562045996478e-12
C33_85 V33 V85 -1.5994391321857484e-19

R33_86 V33 V86 1339.6402599938385
L33_86 V33 V86 4.717649941456908e-12
C33_86 V33 V86 2.4952873818700285e-20

R33_87 V33 V87 3239.705932261485
L33_87 V33 V87 -1.201002124554322e-11
C33_87 V33 V87 -8.628526829543998e-20

R33_88 V33 V88 2985.9592751857695
L33_88 V33 V88 -3.5582517641724173e-12
C33_88 V33 V88 -1.266918828964201e-19

R33_89 V33 V89 52875.63713132314
L33_89 V33 V89 -2.132253057860436e-12
C33_89 V33 V89 -1.0051810284881054e-19

R33_90 V33 V90 -1877.6057321320611
L33_90 V33 V90 -1.605633653745659e-12
C33_90 V33 V90 -2.798793433198066e-19

R33_91 V33 V91 -4449.425471776995
L33_91 V33 V91 1.89254497802538e-12
C33_91 V33 V91 1.9951183873409378e-19

R33_92 V33 V92 -3646.0114760617093
L33_92 V33 V92 2.2895430297710482e-12
C33_92 V33 V92 1.1198485580516984e-19

R33_93 V33 V93 -1135.6183986105368
L33_93 V33 V93 3.0240352596584167e-12
C33_93 V33 V93 1.7905193027719689e-19

R33_94 V33 V94 -2744.75722499311
L33_94 V33 V94 1.683269650754077e-11
C33_94 V33 V94 1.38436703868091e-19

R33_95 V33 V95 -4937.073098619422
L33_95 V33 V95 -9.00819159469556e-12
C33_95 V33 V95 4.209685113460598e-20

R33_96 V33 V96 -2526.3517666017588
L33_96 V33 V96 -6.096690191319962e-12
C33_96 V33 V96 6.567960243032858e-20

R33_97 V33 V97 -1986.9822038981727
L33_97 V33 V97 -4.404372136288886e-11
C33_97 V33 V97 7.67658593455443e-20

R33_98 V33 V98 1008.0323154070496
L33_98 V33 V98 2.4384086346254706e-12
C33_98 V33 V98 1.1178754848442535e-19

R33_99 V33 V99 1733.7133179872878
L33_99 V33 V99 -1.672101387925764e-12
C33_99 V33 V99 -2.545666887664558e-19

R33_100 V33 V100 1140.007619256435
L33_100 V33 V100 -6.401915899189375e-12
C33_100 V33 V100 -1.49374775256229e-19

R33_101 V33 V101 1738.232560532967
L33_101 V33 V101 -3.1401992567410687e-12
C33_101 V33 V101 -5.85607948894453e-20

R33_102 V33 V102 -12510.121706264312
L33_102 V33 V102 -4.5646874546319575e-12
C33_102 V33 V102 -1.2439319709747118e-19

R33_103 V33 V103 8221.749017772017
L33_103 V33 V103 3.5157197746577037e-12
C33_103 V33 V103 2.275439224946669e-20

R33_104 V33 V104 3921.0165524763534
L33_104 V33 V104 2.7190908499359165e-12
C33_104 V33 V104 1.575665180030775e-20

R33_105 V33 V105 -602.5511188353798
L33_105 V33 V105 -5.199256810383238e-12
C33_105 V33 V105 -1.635968769933963e-19

R33_106 V33 V106 37376.763672563015
L33_106 V33 V106 -3.470606153074056e-12
C33_106 V33 V106 -6.210421152028459e-20

R33_107 V33 V107 127447.16553702386
L33_107 V33 V107 2.9409440794135887e-12
C33_107 V33 V107 1.7780401979733308e-19

R33_108 V33 V108 -2938.3088806491933
L33_108 V33 V108 -4.199682673382455e-12
C33_108 V33 V108 1.4146253296595976e-20

R33_109 V33 V109 36497.67106480824
L33_109 V33 V109 1.2948614557537398e-11
C33_109 V33 V109 1.2781821032054383e-19

R33_110 V33 V110 33634.969353400804
L33_110 V33 V110 5.517628771450679e-12
C33_110 V33 V110 5.1019781469158675e-20

R33_111 V33 V111 6764.488642918744
L33_111 V33 V111 3.124720599452937e-11
C33_111 V33 V111 4.237255385567852e-20

R33_112 V33 V112 3788.379903595051
L33_112 V33 V112 4.593557640074078e-12
C33_112 V33 V112 9.113294502820578e-20

R33_113 V33 V113 2996.6406981162195
L33_113 V33 V113 2.3241976158565353e-12
C33_113 V33 V113 2.924398771131538e-19

R33_114 V33 V114 -182925.8766287108
L33_114 V33 V114 3.748335075634471e-12
C33_114 V33 V114 1.2156453672082749e-19

R33_115 V33 V115 -4749.572008019195
L33_115 V33 V115 -1.819383412932428e-12
C33_115 V33 V115 -2.1415375280286498e-19

R33_116 V33 V116 -12311.660553103131
L33_116 V33 V116 -3.9342357683031235e-12
C33_116 V33 V116 -7.896098471307407e-20

R33_117 V33 V117 -984.3418824906478
L33_117 V33 V117 -2.405516006566233e-12
C33_117 V33 V117 -2.3247268224647734e-19

R33_118 V33 V118 3940.8206587019768
L33_118 V33 V118 -3.862229977411702e-12
C33_118 V33 V118 -1.7506589350100864e-19

R33_119 V33 V119 3218.5545496865075
L33_119 V33 V119 2.768571894129751e-11
C33_119 V33 V119 -4.2097186840358614e-20

R33_120 V33 V120 2391.2019647455245
L33_120 V33 V120 -8.33296003885742e-12
C33_120 V33 V120 -1.4199635690865292e-19

R33_121 V33 V121 -3273.6436670032517
L33_121 V33 V121 -2.0749539639379368e-12
C33_121 V33 V121 -3.269024225223016e-20

R33_122 V33 V122 -47312.02511877627
L33_122 V33 V122 -5.769464009946258e-11
C33_122 V33 V122 6.466851851913498e-20

R33_123 V33 V123 -39092.858223294126
L33_123 V33 V123 2.1900988314333086e-12
C33_123 V33 V123 2.252586367744514e-19

R33_124 V33 V124 -5644.257965660083
L33_124 V33 V124 1.838085862978495e-12
C33_124 V33 V124 2.615134315069183e-19

R33_125 V33 V125 4931.531389210446
L33_125 V33 V125 1.9706541561509973e-12
C33_125 V33 V125 5.91182112840505e-20

R33_126 V33 V126 9418.430087251323
L33_126 V33 V126 2.458798501223252e-12
C33_126 V33 V126 1.1663239256483978e-19

R33_127 V33 V127 -6838.479535306498
L33_127 V33 V127 -1.1271689174254261e-11
C33_127 V33 V127 -3.14254718309088e-20

R33_128 V33 V128 -3744.6694172954844
L33_128 V33 V128 -4.788675963736516e-12
C33_128 V33 V128 8.606183155944452e-21

R33_129 V33 V129 -1588.5101043564894
L33_129 V33 V129 -8.130558109775056e-12
C33_129 V33 V129 6.571954481945122e-20

R33_130 V33 V130 -6731.756692394815
L33_130 V33 V130 -2.409484021832997e-12
C33_130 V33 V130 -1.7675725339294015e-19

R33_131 V33 V131 4059.4682338281877
L33_131 V33 V131 -5.69760592672242e-12
C33_131 V33 V131 -1.1874931957496703e-19

R33_132 V33 V132 2036.1428382266627
L33_132 V33 V132 -2.9060131355457174e-12
C33_132 V33 V132 -2.5649901800616583e-19

R33_133 V33 V133 -7011.93454121898
L33_133 V33 V133 -7.728117682561825e-12
C33_133 V33 V133 5.737841860510387e-20

R33_134 V33 V134 3062.3679109009654
L33_134 V33 V134 2.6119189545857744e-12
C33_134 V33 V134 1.452015784744009e-19

R33_135 V33 V135 -11871.63613859853
L33_135 V33 V135 3.4335377362619807e-12
C33_135 V33 V135 1.387952344894436e-19

R33_136 V33 V136 -7430.251007905734
L33_136 V33 V136 2.1898487333413782e-12
C33_136 V33 V136 1.946001095270325e-19

R33_137 V33 V137 3575.491302677266
L33_137 V33 V137 3.8898913226381805e-12
C33_137 V33 V137 -1.428137853440257e-19

R33_138 V33 V138 -2860.365023720865
L33_138 V33 V138 6.7198916816868636e-12
C33_138 V33 V138 5.7220977890375974e-21

R33_139 V33 V139 -8844.941714117253
L33_139 V33 V139 -2.0787755190514696e-12
C33_139 V33 V139 -1.6359755706120627e-19

R33_140 V33 V140 14678.087786256901
L33_140 V33 V140 -2.772541260544e-12
C33_140 V33 V140 -1.1329556447435182e-19

R33_141 V33 V141 2076.0861267587657
L33_141 V33 V141 9.845362027338297e-12
C33_141 V33 V141 1.2347295364110998e-19

R33_142 V33 V142 21239.608825012092
L33_142 V33 V142 -1.4976130352808683e-12
C33_142 V33 V142 -8.290691893822952e-20

R33_143 V33 V143 3243.107374200252
L33_143 V33 V143 3.955544300361924e-12
C33_143 V33 V143 1.0547915626334099e-19

R33_144 V33 V144 -26643.746644530616
L33_144 V33 V144 -1.014710250351838e-11
C33_144 V33 V144 1.192979274980774e-20

R33_145 V33 V145 -707.5852434896756
L33_145 V33 V145 -4.586566781424113e-12
C33_145 V33 V145 2.0182551338630141e-19

R33_146 V33 V146 4295.401078165433
L33_146 V33 V146 7.1893784630942115e-12
C33_146 V33 V146 -2.073128759580662e-20

R33_147 V33 V147 -3554.2343007677523
L33_147 V33 V147 3.2564529068291635e-12
C33_147 V33 V147 1.1913243916820995e-19

R33_148 V33 V148 3713.29422181321
L33_148 V33 V148 1.7969789791969396e-12
C33_148 V33 V148 1.0120384090411725e-19

R33_149 V33 V149 2499.9342569300265
L33_149 V33 V149 -1.0338121739142887e-12
C33_149 V33 V149 -4.581821065106503e-19

R33_150 V33 V150 4148.404881555464
L33_150 V33 V150 1.4363243762585745e-12
C33_150 V33 V150 2.2126204180765394e-19

R33_151 V33 V151 19192.338341164235
L33_151 V33 V151 -4.26772676057565e-12
C33_151 V33 V151 -1.1214334278187032e-19

R33_152 V33 V152 -14805.987339087333
L33_152 V33 V152 -5.641474514361297e-12
C33_152 V33 V152 -3.7361023051306e-21

R33_153 V33 V153 -61072.87544530863
L33_153 V33 V153 3.462247859313137e-12
C33_153 V33 V153 -3.291782582701209e-20

R33_154 V33 V154 -4925.837725281901
L33_154 V33 V154 -6.3188663455532665e-12
C33_154 V33 V154 -1.3211446530348095e-19

R33_155 V33 V155 -2911.4046610580276
L33_155 V33 V155 -1.8538108910077525e-12
C33_155 V33 V155 -1.2020973637382667e-19

R33_156 V33 V156 3750.078164801872
L33_156 V33 V156 -1.663034936607332e-11
C33_156 V33 V156 -1.1042509229114905e-19

R33_157 V33 V157 -1753.679155013399
L33_157 V33 V157 8.582467104760694e-13
C33_157 V33 V157 4.878122107188262e-19

R33_158 V33 V158 2728.5595388508286
L33_158 V33 V158 -2.135599409691841e-12
C33_158 V33 V158 -2.3552410678642223e-20

R33_159 V33 V159 1749.9316483917794
L33_159 V33 V159 3.11604851135539e-12
C33_159 V33 V159 4.21683352133678e-20

R33_160 V33 V160 -37000.92952729704
L33_160 V33 V160 -2.3912944939157058e-11
C33_160 V33 V160 -5.443544176590891e-21

R33_161 V33 V161 -5909.361462565756
L33_161 V33 V161 -3.844952063556268e-12
C33_161 V33 V161 -6.361650594757942e-20

R33_162 V33 V162 35580.52287739394
L33_162 V33 V162 -4.467427003254291e-12
C33_162 V33 V162 -6.64454275104901e-20

R33_163 V33 V163 2559.5352568972435
L33_163 V33 V163 3.627466123052963e-12
C33_163 V33 V163 3.1497866977714414e-20

R33_164 V33 V164 1765.22313673266
L33_164 V33 V164 7.307061038842981e-12
C33_164 V33 V164 -5.0084634277231436e-20

R33_165 V33 V165 -814.9975701429876
L33_165 V33 V165 -1.0298473757848252e-12
C33_165 V33 V165 -2.1066478056043758e-19

R33_166 V33 V166 4040.1366429989025
L33_166 V33 V166 2.518928733858346e-12
C33_166 V33 V166 5.729681193252104e-20

R33_167 V33 V167 4422.973125492134
L33_167 V33 V167 -7.720095060675834e-12
C33_167 V33 V167 1.3444143269903862e-20

R33_168 V33 V168 -7360.740107005955
L33_168 V33 V168 -9.076386028267063e-12
C33_168 V33 V168 7.512478117174909e-20

R33_169 V33 V169 2961.5202846202537
L33_169 V33 V169 1.0892875661047228e-11
C33_169 V33 V169 1.4622163674635971e-19

R33_170 V33 V170 -1522.2670149400492
L33_170 V33 V170 -4.364031159436722e-12
C33_170 V33 V170 -9.144232925625586e-20

R33_171 V33 V171 -943.1576798551993
L33_171 V33 V171 -2.001505955337508e-12
C33_171 V33 V171 -1.3324401482738702e-19

R33_172 V33 V172 -1502.534945599652
L33_172 V33 V172 -2.5939325648767636e-11
C33_172 V33 V172 -6.469835091803011e-20

R33_173 V33 V173 -5813.998913560611
L33_173 V33 V173 1.2534345889625776e-12
C33_173 V33 V173 1.3082072916999117e-20

R33_174 V33 V174 5666.062095121217
L33_174 V33 V174 -3.885937382427242e-12
C33_174 V33 V174 1.0044864479076414e-19

R33_175 V33 V175 1292.3441424342639
L33_175 V33 V175 1.336601480760598e-09
C33_175 V33 V175 -7.670384932010973e-20

R33_176 V33 V176 1222.4630934018055
L33_176 V33 V176 -1.2577152274158156e-08
C33_176 V33 V176 -8.50099744769092e-20

R33_177 V33 V177 -1711.0632185102725
L33_177 V33 V177 -1.7011276065062764e-12
C33_177 V33 V177 -1.0204515103444189e-19

R33_178 V33 V178 1760.6462970544574
L33_178 V33 V178 1.7764550404969152e-12
C33_178 V33 V178 6.596616083568371e-20

R33_179 V33 V179 5787.401847340496
L33_179 V33 V179 1.573483320245668e-12
C33_179 V33 V179 2.3774397316063625e-19

R33_180 V33 V180 4194.744954775202
L33_180 V33 V180 2.1550804705949207e-12
C33_180 V33 V180 1.8442527689653728e-19

R33_181 V33 V181 1410.8738598870214
L33_181 V33 V181 3.3880147164669927e-12
C33_181 V33 V181 1.2374514286451114e-19

R33_182 V33 V182 -1823.6349240886984
L33_182 V33 V182 -2.2406062440991273e-12
C33_182 V33 V182 -1.160472570084023e-19

R33_183 V33 V183 -3418.8779524646493
L33_183 V33 V183 3.977236110224731e-12
C33_183 V33 V183 2.6579189975755438e-20

R33_184 V33 V184 -1628.7325396506913
L33_184 V33 V184 1.2745579680474027e-11
C33_184 V33 V184 -1.4375943713966817e-20

R33_185 V33 V185 -15020.43659757174
L33_185 V33 V185 2.885126238700291e-12
C33_185 V33 V185 -1.7070049019167093e-20

R33_186 V33 V186 -2052.109699383041
L33_186 V33 V186 -1.7777582957349295e-12
C33_186 V33 V186 -5.392191215983828e-21

R33_187 V33 V187 -3392.539720343892
L33_187 V33 V187 -1.1836844125095208e-12
C33_187 V33 V187 -2.092349329476492e-19

R33_188 V33 V188 -1786.7587015638167
L33_188 V33 V188 -9.959785320892433e-13
C33_188 V33 V188 -1.574265208232308e-19

R33_189 V33 V189 1527.7613483984633
L33_189 V33 V189 -1.5038757927176134e-12
C33_189 V33 V189 -1.115584842381364e-19

R33_190 V33 V190 1861.4462056804573
L33_190 V33 V190 3.06318453884741e-12
C33_190 V33 V190 1.1490022025874059e-19

R33_191 V33 V191 4383.193847154396
L33_191 V33 V191 -4.165466027118607e-12
C33_191 V33 V191 -4.101307026931242e-20

R33_192 V33 V192 1760.6090129638928
L33_192 V33 V192 3.2046315519502467e-12
C33_192 V33 V192 1.1687376585840909e-20

R33_193 V33 V193 -919.5381631051707
L33_193 V33 V193 3.809250323539359e-12
C33_193 V33 V193 1.2358831165333051e-19

R33_194 V33 V194 1817.532337996262
L33_194 V33 V194 2.417322628187832e-12
C33_194 V33 V194 7.440133057559432e-20

R33_195 V33 V195 4633.172440426632
L33_195 V33 V195 1.3017349858147819e-12
C33_195 V33 V195 1.4880617394194473e-19

R33_196 V33 V196 1931.200609178654
L33_196 V33 V196 1.784193108778906e-12
C33_196 V33 V196 9.124642252405955e-20

R33_197 V33 V197 -7363.371123546328
L33_197 V33 V197 2.8795185395610657e-12
C33_197 V33 V197 -2.157968302814399e-21

R33_198 V33 V198 -2211.2689842638897
L33_198 V33 V198 -3.272039515944128e-12
C33_198 V33 V198 -2.9659838155300635e-20

R33_199 V33 V199 -2963.871314275057
L33_199 V33 V199 -3.904550992541842e-11
C33_199 V33 V199 4.252730310659269e-20

R33_200 V33 V200 -986.5113083337874
L33_200 V33 V200 -4.010882469413108e-12
C33_200 V33 V200 -2.224450897991351e-21

R34_34 V34 0 -1995.5354924680557
L34_34 V34 0 -6.223563570591572e-13
C34_34 V34 0 -5.908473165196484e-19

R34_35 V34 V35 -5381.075871121176
L34_35 V34 V35 -2.484798826473869e-12
C34_35 V34 V35 -1.4168723814156816e-19

R34_36 V34 V36 -3341.6892801933827
L34_36 V34 V36 -1.7269073439523731e-12
C34_36 V34 V36 -2.1653673049189957e-19

R34_37 V34 V37 -9360.982911499808
L34_37 V34 V37 1.8074202055211832e-11
C34_37 V34 V37 2.299883935687737e-20

R34_38 V34 V38 -10253.518160407059
L34_38 V34 V38 2.831163870695589e-12
C34_38 V34 V38 2.312878608856959e-19

R34_39 V34 V39 -4908.430473638767
L34_39 V34 V39 4.232801481672105e-12
C34_39 V34 V39 9.494590112581466e-20

R34_40 V34 V40 -2712.405397680733
L34_40 V34 V40 3.4010597403623215e-12
C34_40 V34 V40 1.1239350121884258e-19

R34_41 V34 V41 9683.006781134165
L34_41 V34 V41 6.32988757769634e-12
C34_41 V34 V41 2.6558279389622898e-20

R34_42 V34 V42 -8344.939110890444
L34_42 V34 V42 8.722402574355968e-13
C34_42 V34 V42 8.392760293079779e-19

R34_43 V34 V43 17248.402454480605
L34_43 V34 V43 6.182001837453767e-12
C34_43 V34 V43 1.4297376326892377e-19

R34_44 V34 V44 11559.347062049823
L34_44 V34 V44 3.4307344037158524e-12
C34_44 V34 V44 2.21553456770813e-19

R34_45 V34 V45 4559.750773888841
L34_45 V34 V45 5.122531183632942e-12
C34_45 V34 V45 5.1353049119464036e-20

R34_46 V34 V46 2190.293626037876
L34_46 V34 V46 2.6560055273959205e-12
C34_46 V34 V46 -8.182083179582902e-20

R34_47 V34 V47 5578.877641909281
L34_47 V34 V47 6.166562280444011e-11
C34_47 V34 V47 -5.172164757949652e-20

R34_48 V34 V48 2815.0492225816583
L34_48 V34 V48 6.700249552805441e-12
C34_48 V34 V48 -8.907745906204578e-23

R34_49 V34 V49 -16919.901439923455
L34_49 V34 V49 -3.6293098005216096e-12
C34_49 V34 V49 -7.87205493392497e-20

R34_50 V34 V50 3107.175708667014
L34_50 V34 V50 -1.114439457199961e-12
C34_50 V34 V50 -5.28857934574404e-19

R34_51 V34 V51 -247506.21156950513
L34_51 V34 V51 -2.8177623372481643e-12
C34_51 V34 V51 -2.0104300525852824e-19

R34_52 V34 V52 -14037.887341098343
L34_52 V34 V52 -1.9831739653779756e-12
C34_52 V34 V52 -2.9548866035220694e-19

R34_53 V34 V53 -28813.42373209113
L34_53 V34 V53 -4.159723891449588e-12
C34_53 V34 V53 -3.651721824334224e-20

R34_54 V34 V54 -2448.818019739246
L34_54 V34 V54 -2.368308963717688e-12
C34_54 V34 V54 2.357407105904993e-20

R34_55 V34 V55 -9804.843830708125
L34_55 V34 V55 8.295251511867134e-12
C34_55 V34 V55 1.413706812956425e-19

R34_56 V34 V56 -3278.981679747177
L34_56 V34 V56 -2.1139602201996895e-11
C34_56 V34 V56 1.018603261066314e-19

R34_57 V34 V57 -14345.70902748913
L34_57 V34 V57 3.4019166006668192e-12
C34_57 V34 V57 1.2565156753214274e-19

R34_58 V34 V58 7523.2025391433435
L34_58 V34 V58 1.2650447517194122e-12
C34_58 V34 V58 3.531402896094299e-19

R34_59 V34 V59 133902.20018976263
L34_59 V34 V59 2.636131772002853e-12
C34_59 V34 V59 1.6484601101938282e-19

R34_60 V34 V60 -27464.01228644245
L34_60 V34 V60 1.8037322040034759e-12
C34_60 V34 V60 2.619135884658315e-19

R34_61 V34 V61 13720.64360313283
L34_61 V34 V61 -2.6790090346028054e-11
C34_61 V34 V61 -7.965057255684678e-20

R34_62 V34 V62 -3298.094838170226
L34_62 V34 V62 -5.102288464301651e-12
C34_62 V34 V62 -1.098487808139228e-19

R34_63 V34 V63 74369.47249650041
L34_63 V34 V63 -4.499141789176784e-12
C34_63 V34 V63 -1.5410325204182722e-19

R34_64 V34 V64 8097.295327989684
L34_64 V34 V64 -4.59658455722436e-12
C34_64 V34 V64 -2.202970007792477e-19

R34_65 V34 V65 7273.879128223239
L34_65 V34 V65 5.821475036826927e-11
C34_65 V34 V65 1.5967112537745466e-20

R34_66 V34 V66 1995.2560978757563
L34_66 V34 V66 2.6336181458542398e-11
C34_66 V34 V66 -4.7817780170192405e-20

R34_67 V34 V67 186460.05772924042
L34_67 V34 V67 -4.913751975292529e-12
C34_67 V34 V67 -7.968918789203594e-20

R34_68 V34 V68 8071.047770156865
L34_68 V34 V68 -8.103596865863852e-12
C34_68 V34 V68 -6.608254925775006e-20

R34_69 V34 V69 -8636.153508677255
L34_69 V34 V69 -1.48035721215168e-11
C34_69 V34 V69 9.666750094812823e-20

R34_70 V34 V70 59687.60393593989
L34_70 V34 V70 3.832919039148839e-12
C34_70 V34 V70 9.853983459592331e-20

R34_71 V34 V71 14326.614109862074
L34_71 V34 V71 4.645692707388155e-12
C34_71 V34 V71 8.563845031422972e-20

R34_72 V34 V72 12346.308492447737
L34_72 V34 V72 5.498222810968408e-12
C34_72 V34 V72 1.162864809827658e-19

R34_73 V34 V73 8990.772804059085
L34_73 V34 V73 -2.3120013843536966e-11
C34_73 V34 V73 -1.1376934654785805e-19

R34_74 V34 V74 -1617.9410935250112
L34_74 V34 V74 -2.2188373645453345e-12
C34_74 V34 V74 -1.367096224521536e-19

R34_75 V34 V75 9624.376602712406
L34_75 V34 V75 4.369806165370243e-12
C34_75 V34 V75 1.0116285578158914e-19

R34_76 V34 V76 -4487.473864450537
L34_76 V34 V76 -1.5799135910585762e-11
C34_76 V34 V76 1.2838101767659651e-20

R34_77 V34 V77 -6100.340990493
L34_77 V34 V77 8.705975001211948e-12
C34_77 V34 V77 1.9490620906702816e-20

R34_78 V34 V78 1233.931052106918
L34_78 V34 V78 -1.985605727699272e-11
C34_78 V34 V78 -9.749755727337757e-20

R34_79 V34 V79 -5388.3667873501645
L34_79 V34 V79 -5.1646553953194095e-12
C34_79 V34 V79 -4.870639635286683e-20

R34_80 V34 V80 -114352.03989267543
L34_80 V34 V80 6.124963642407238e-11
C34_80 V34 V80 -2.6085670842436218e-20

R34_81 V34 V81 2434.489758681029
L34_81 V34 V81 6.547060846459526e-12
C34_81 V34 V81 1.3300709031386977e-19

R34_82 V34 V82 -2712.179287417504
L34_82 V34 V82 1.2838140898631372e-12
C34_82 V34 V82 3.928056915691586e-19

R34_83 V34 V83 -12570.175318804177
L34_83 V34 V83 -7.939311180866032e-12
C34_83 V34 V83 -1.275712067781528e-19

R34_84 V34 V84 14932.653631650197
L34_84 V34 V84 7.852729875598252e-12
C34_84 V34 V84 -5.872150689476374e-20

R34_85 V34 V85 -5216.657366723886
L34_85 V34 V85 -9.930856007794922e-12
C34_85 V34 V85 -7.480294944749894e-20

R34_86 V34 V86 111994.90924162944
L34_86 V34 V86 5.051286599663686e-12
C34_86 V34 V86 -1.0260709840618686e-19

R34_87 V34 V87 6426.430763119929
L34_87 V34 V87 1.1888480371278886e-11
C34_87 V34 V87 8.766647019002961e-20

R34_88 V34 V88 6610.616614010608
L34_88 V34 V88 -1.6248412923985146e-11
C34_88 V34 V88 7.582629483210835e-20

R34_89 V34 V89 -7778.456237907644
L34_89 V34 V89 -3.3976167178789466e-12
C34_89 V34 V89 -6.28682797399855e-20

R34_90 V34 V90 2400.2329177641395
L34_90 V34 V90 -7.114264237201443e-13
C34_90 V34 V90 -4.936068401850425e-19

R34_91 V34 V91 8165.077433602874
L34_91 V34 V91 2.972863945294805e-12
C34_91 V34 V91 1.0627925210838583e-19

R34_92 V34 V92 -4781.653763424685
L34_92 V34 V92 4.7811245081968565e-12
C34_92 V34 V92 1.1706384549318338e-20

R34_93 V34 V93 2462.780941148473
L34_93 V34 V93 5.957355409451955e-12
C34_93 V34 V93 8.288060576335608e-20

R34_94 V34 V94 -1433.6737030589036
L34_94 V34 V94 1.385156471456823e-12
C34_94 V34 V94 5.319877122506538e-19

R34_95 V34 V95 -4849.381493832179
L34_95 V34 V95 -7.167458965661641e-12
C34_95 V34 V95 -7.144120231008967e-20

R34_96 V34 V96 -2860.529473067728
L34_96 V34 V96 -5.747664145175999e-12
C34_96 V34 V96 -6.129411316797371e-20

R34_97 V34 V97 -3016.081563805959
L34_97 V34 V97 3.053497733354104e-12
C34_97 V34 V97 8.788903826113479e-20

R34_98 V34 V98 6032.202451723447
L34_98 V34 V98 1.3436923720501445e-12
C34_98 V34 V98 1.2689306077658813e-19

R34_99 V34 V99 -6322.750381624854
L34_99 V34 V99 -1.998224497070539e-12
C34_99 V34 V99 -1.0136050702760869e-19

R34_100 V34 V100 2588.078603317627
L34_100 V34 V100 -5.113702223210039e-12
C34_100 V34 V100 -6.733873243717796e-21

R34_101 V34 V101 20726.886393957728
L34_101 V34 V101 -2.001526107436283e-12
C34_101 V34 V101 -9.447112263393525e-20

R34_102 V34 V102 1519.5874340111575
L34_102 V34 V102 -9.652896975283933e-13
C34_102 V34 V102 -6.934655853055962e-19

R34_103 V34 V103 6650.6902815601115
L34_103 V34 V103 2.6667709539830363e-12
C34_103 V34 V103 7.382518516901458e-20

R34_104 V34 V104 12327.337998966981
L34_104 V34 V104 1.950426110930759e-12
C34_104 V34 V104 1.0714322532651464e-19

R34_105 V34 V105 4457.556167159505
L34_105 V34 V105 -1.1195730918345546e-11
C34_105 V34 V105 -3.9329051527280627e-20

R34_106 V34 V106 -3776.0353817365763
L34_106 V34 V106 5.062855038183399e-11
C34_106 V34 V106 2.968633430142833e-19

R34_107 V34 V107 7266.85907644016
L34_107 V34 V107 8.875237156728498e-12
C34_107 V34 V107 1.5517657139111712e-20

R34_108 V34 V108 -3113.0304342770673
L34_108 V34 V108 -2.8329209427731958e-12
C34_108 V34 V108 -1.0390781558258092e-19

R34_109 V34 V109 -68862.55890337338
L34_109 V34 V109 2.7397797057426114e-12
C34_109 V34 V109 6.76078499247096e-20

R34_110 V34 V110 -2522.487565098333
L34_110 V34 V110 1.3394939252317612e-12
C34_110 V34 V110 5.56357203987335e-19

R34_111 V34 V111 9077.153865687042
L34_111 V34 V111 -3.873167486509465e-12
C34_111 V34 V111 -3.5287405266168734e-20

R34_112 V34 V112 3622.7601698693
L34_112 V34 V112 -4.658272106904623e-12
C34_112 V34 V112 -9.070474287481445e-20

R34_113 V34 V113 5834.340147102606
L34_113 V34 V113 -9.329759387836757e-12
C34_113 V34 V113 8.006556366209048e-20

R34_114 V34 V114 2794.2128695495294
L34_114 V34 V114 -3.5757087920098994e-12
C34_114 V34 V114 -4.874270595706483e-19

R34_115 V34 V115 -2444.3440824213167
L34_115 V34 V115 -1.3521478408230117e-11
C34_115 V34 V115 -4.5635077223956854e-20

R34_116 V34 V116 -9716.722506095743
L34_116 V34 V116 3.7704514688000874e-12
C34_116 V34 V116 1.1612122464044026e-19

R34_117 V34 V117 -1636.6241179920657
L34_117 V34 V117 -3.5304007043389783e-12
C34_117 V34 V117 -5.320091692736787e-20

R34_118 V34 V118 -1823.9737975017067
L34_118 V34 V118 -1.363135664476858e-12
C34_118 V34 V118 -3.582541951245627e-19

R34_119 V34 V119 19154.7545188695
L34_119 V34 V119 8.188027040736658e-12
C34_119 V34 V119 3.161017216235755e-20

R34_120 V34 V120 116985.6503522587
L34_120 V34 V120 -4.213665237604494e-11
C34_120 V34 V120 -1.3776127649745537e-20

R34_121 V34 V121 2937.702672446174
L34_121 V34 V121 2.567623563743788e-11
C34_121 V34 V121 -6.897205508779775e-20

R34_122 V34 V122 2061.175639809521
L34_122 V34 V122 1.2843927937503822e-12
C34_122 V34 V122 5.622424543625425e-19

R34_123 V34 V123 4039.8603237313937
L34_123 V34 V123 -6.446630557805113e-12
C34_123 V34 V123 -4.092981324164991e-20

R34_124 V34 V124 4949.323496453116
L34_124 V34 V124 -4.940292463953603e-12
C34_124 V34 V124 -1.2405442849091057e-19

R34_125 V34 V125 1053.5917740132256
L34_125 V34 V125 7.591679953993365e-12
C34_125 V34 V125 1.1066379730884095e-20

R34_126 V34 V126 1078.4460875293044
L34_126 V34 V126 1.8624977112678976e-11
C34_126 V34 V126 2.648789695145516e-20

R34_127 V34 V127 -7407945.949025867
L34_127 V34 V127 -2.2505728016653377e-10
C34_127 V34 V127 2.3666022130343052e-21

R34_128 V34 V128 -26286.159115652958
L34_128 V34 V128 -9.409005090927503e-12
C34_128 V34 V128 5.657233244369247e-20

R34_129 V34 V129 -1003.6235921973123
L34_129 V34 V129 -2.6176675782135872e-11
C34_129 V34 V129 1.7221752027725137e-19

R34_130 V34 V130 -700.8596566344826
L34_130 V34 V130 -2.100197924729681e-12
C34_130 V34 V130 -3.5150724075144972e-19

R34_131 V34 V131 -5424.409577884001
L34_131 V34 V131 5.03095863818877e-12
C34_131 V34 V131 4.6211899989891075e-20

R34_132 V34 V132 -2870.4063522837937
L34_132 V34 V132 3.1453479834180044e-12
C34_132 V34 V132 4.20817839146828e-20

R34_133 V34 V133 -1706.5438784479113
L34_133 V34 V133 -5.9287590724807796e-12
C34_133 V34 V133 -1.0843906239159415e-19

R34_134 V34 V134 1743.718681698577
L34_134 V34 V134 3.00434742577173e-12
C34_134 V34 V134 2.55520195608082e-19

R34_135 V34 V135 8439.274614930338
L34_135 V34 V135 -6.829608324071479e-12
C34_135 V34 V135 -3.334796943869864e-20

R34_136 V34 V136 6093.496684606998
L34_136 V34 V136 2.7405293291507178e-11
C34_136 V34 V136 -3.601555643345311e-20

R34_137 V34 V137 632.5852398546637
L34_137 V34 V137 -9.413912218115119e-12
C34_137 V34 V137 -1.6501355501375121e-19

R34_138 V34 V138 1380.697649213028
L34_138 V34 V138 2.1860939004248133e-11
C34_138 V34 V138 -2.432713629235793e-20

R34_139 V34 V139 33580.34766689645
L34_139 V34 V139 -4.5329472134302704e-12
C34_139 V34 V139 -5.098914905386213e-20

R34_140 V34 V140 1557.643855511597
L34_140 V34 V140 -3.3716267747531746e-12
C34_140 V34 V140 -2.5674123290793475e-20

R34_141 V34 V141 -7300.111678733747
L34_141 V34 V141 1.644536110955044e-12
C34_141 V34 V141 2.333621900544919e-19

R34_142 V34 V142 -631.4693128372467
L34_142 V34 V142 5.829663698801955e-12
C34_142 V34 V142 -1.2809685252202348e-20

R34_143 V34 V143 -5062.682421789951
L34_143 V34 V143 3.432774894442579e-12
C34_143 V34 V143 1.0639997947707113e-19

R34_144 V34 V144 -883.2174466091744
L34_144 V34 V144 1.3184797229228017e-11
C34_144 V34 V144 6.297490799641324e-20

R34_145 V34 V145 -635.1786870037748
L34_145 V34 V145 7.2369499283395456e-12
C34_145 V34 V145 1.3779721562928406e-19

R34_146 V34 V146 -5195.288592978318
L34_146 V34 V146 -4.640634123339506e-12
C34_146 V34 V146 -9.88984541455865e-20

R34_147 V34 V147 -2168.045470276411
L34_147 V34 V147 1.1049839379784645e-11
C34_147 V34 V147 -7.327354759598339e-21

R34_148 V34 V148 870.5659866440692
L34_148 V34 V148 2.6471779908182513e-12
C34_148 V34 V148 2.40754654829838e-21

R34_149 V34 V149 11865.103124377038
L34_149 V34 V149 -6.06756045174636e-13
C34_149 V34 V149 -3.6385445700611063e-19

R34_150 V34 V150 568.3815902244291
L34_150 V34 V150 -2.494218156275198e-12
C34_150 V34 V150 1.7255222128378757e-19

R34_151 V34 V151 1931.5432814628002
L34_151 V34 V151 9.726457818299147e-12
C34_151 V34 V151 -3.281896438313072e-20

R34_152 V34 V152 -1273.1991139403758
L34_152 V34 V152 1.797725047309547e-11
C34_152 V34 V152 1.177982642854257e-20

R34_153 V34 V153 602.8344053005384
L34_153 V34 V153 3.77984003361552e-12
C34_153 V34 V153 -4.120570158510456e-20

R34_154 V34 V154 1112.447032567627
L34_154 V34 V154 1.5932216522048753e-12
C34_154 V34 V154 -8.097597836976299e-20

R34_155 V34 V155 -908.7324871984677
L34_155 V34 V155 -3.1015664135419366e-12
C34_155 V34 V155 -7.871074574357162e-20

R34_156 V34 V156 784.8849695721362
L34_156 V34 V156 -7.708325799633036e-11
C34_156 V34 V156 -2.7758052252153705e-20

R34_157 V34 V157 3689.462800557873
L34_157 V34 V157 5.467082107713685e-13
C34_157 V34 V157 2.9080422133003164e-19

R34_158 V34 V158 -440.4792567146318
L34_158 V34 V158 2.1924321837218354e-12
C34_158 V34 V158 2.698702224523357e-20

R34_159 V34 V159 771.7359839301555
L34_159 V34 V159 -6.396345772891658e-12
C34_159 V34 V159 -2.751432681869491e-20

R34_160 V34 V160 -2720.166209881909
L34_160 V34 V160 -2.3014828850353233e-12
C34_160 V34 V160 -7.71153895014896e-20

R34_161 V34 V161 -1603.4735241263766
L34_161 V34 V161 -2.1851139798864435e-12
C34_161 V34 V161 5.3166660896583067e-20

R34_162 V34 V162 -1163.3515577340313
L34_162 V34 V162 -7.715296488800748e-13
C34_162 V34 V162 -9.896791721474259e-20

R34_163 V34 V163 -5456.916988773691
L34_163 V34 V163 4.130904604648941e-12
C34_163 V34 V163 7.894369277766478e-20

R34_164 V34 V164 1474.5630482488443
L34_164 V34 V164 8.30959096801112e-12
C34_164 V34 V164 3.4484801314057575e-20

R34_165 V34 V165 -149567.23735469196
L34_165 V34 V165 -9.108321754518758e-13
C34_165 V34 V165 -1.799280195957319e-19

R34_166 V34 V166 261.56677597899665
L34_166 V34 V166 -3.3124862370760384e-12
C34_166 V34 V166 4.70457442922265e-20

R34_167 V34 V167 -1835.6459806416647
L34_167 V34 V167 4.091670476528394e-12
C34_167 V34 V167 4.2562860765593604e-20

R34_168 V34 V168 -460.71240929599253
L34_168 V34 V168 4.177177553286025e-12
C34_168 V34 V168 9.108439947647475e-20

R34_169 V34 V169 1783.0345655050928
L34_169 V34 V169 2.1989273007415107e-12
C34_169 V34 V169 6.368495025458505e-21

R34_170 V34 V170 -630.5527179050989
L34_170 V34 V170 7.1510896391686e-13
C34_170 V34 V170 -6.705738042500411e-20

R34_171 V34 V171 -9265.669928396283
L34_171 V34 V171 -1.6846550763315887e-12
C34_171 V34 V171 -1.7463286088058797e-19

R34_172 V34 V172 1920.914326017257
L34_172 V34 V172 -3.689617238392835e-12
C34_172 V34 V172 -1.1518662670523284e-19

R34_173 V34 V173 5027.022627469893
L34_173 V34 V173 1.5662932200121407e-12
C34_173 V34 V173 4.84947475126025e-20

R34_174 V34 V174 -270.4332589609454
L34_174 V34 V174 -2.1052381694232935e-12
C34_174 V34 V174 1.2250847051535621e-20

R34_175 V34 V175 1765.5521067761308
L34_175 V34 V175 -4.162794409778445e-11
C34_175 V34 V175 -1.0974266677998099e-20

R34_176 V34 V176 760.1461598621402
L34_176 V34 V176 -3.7664387400597595e-11
C34_176 V34 V176 -1.2752929563660092e-20

R34_177 V34 V177 10424.285557804391
L34_177 V34 V177 -3.0539586082445827e-12
C34_177 V34 V177 -6.160131723725208e-20

R34_178 V34 V178 336.1399364910799
L34_178 V34 V178 -1.2283252264838717e-12
C34_178 V34 V178 1.1232972392919555e-19

R34_179 V34 V179 -4118.560625681427
L34_179 V34 V179 1.37320844259955e-12
C34_179 V34 V179 1.407073126586941e-19

R34_180 V34 V180 -2521.9353664901705
L34_180 V34 V180 1.3351555621366185e-12
C34_180 V34 V180 9.361759553737661e-20

R34_181 V34 V181 -3045.34159006637
L34_181 V34 V181 -1.3927527519563385e-11
C34_181 V34 V181 9.975174371759932e-20

R34_182 V34 V182 6145.734301877385
L34_182 V34 V182 3.376454530933945e-12
C34_182 V34 V182 -9.992991228339172e-20

R34_183 V34 V183 3041.445816259247
L34_183 V34 V183 5.165412631068341e-12
C34_183 V34 V183 3.6340686894028916e-20

R34_184 V34 V184 -12810.65579459572
L34_184 V34 V184 -9.06373404439764e-12
C34_184 V34 V184 2.1372979612628162e-21

R34_185 V34 V185 2088.625866005609
L34_185 V34 V185 2.354878038462659e-12
C34_185 V34 V185 -1.506513563012107e-20

R34_186 V34 V186 -509.7334517071761
L34_186 V34 V186 -9.283545430238321e-12
C34_186 V34 V186 -4.8301424022450564e-20

R34_187 V34 V187 -1900.714372479099
L34_187 V34 V187 -1.368461339987944e-12
C34_187 V34 V187 -1.0173497873014485e-19

R34_188 V34 V188 -1471.8035590644147
L34_188 V34 V188 -1.35892340792419e-12
C34_188 V34 V188 -4.643135679289288e-20

R34_189 V34 V189 3815.9158839714646
L34_189 V34 V189 -2.853372247676744e-12
C34_189 V34 V189 -1.2849722003808608e-19

R34_190 V34 V190 1861.638270446154
L34_190 V34 V190 -3.0980733828053985e-12
C34_190 V34 V190 1.2520431219246708e-19

R34_191 V34 V191 6831.220661725636
L34_191 V34 V191 -2.8461766392209844e-12
C34_191 V34 V191 -1.0972536656444116e-19

R34_192 V34 V192 1608.4439590626464
L34_192 V34 V192 8.759885866085042e-12
C34_192 V34 V192 -1.2954671767610436e-19

R34_193 V34 V193 -1359.4712150928672
L34_193 V34 V193 -6.178711913810452e-12
C34_193 V34 V193 5.805575833823333e-20

R34_194 V34 V194 3442.8990780524123
L34_194 V34 V194 1.4769406176540442e-12
C34_194 V34 V194 -2.5812069386769114e-20

R34_195 V34 V195 1896.4072870960954
L34_195 V34 V195 1.1484992194208386e-12
C34_195 V34 V195 1.7529893558600226e-19

R34_196 V34 V196 1501.2660292547146
L34_196 V34 V196 1.5011393186850011e-12
C34_196 V34 V196 2.3057984502143575e-19

R34_197 V34 V197 5697.806645569057
L34_197 V34 V197 1.6098734478033171e-12
C34_197 V34 V197 1.1168343407933888e-19

R34_198 V34 V198 -3042.201143551481
L34_198 V34 V198 -7.661590051745044e-12
C34_198 V34 V198 -3.300476496463165e-20

R34_199 V34 V199 -6028.565128732993
L34_199 V34 V199 5.029074214904187e-12
C34_199 V34 V199 8.34051055371903e-20

R34_200 V34 V200 -931.5809440001142
L34_200 V34 V200 -1.5795656664181087e-10
C34_200 V34 V200 4.6214177209851105e-20

R35_35 V35 0 -519.0121970008779
L35_35 V35 0 -6.378319272098668e-13
C35_35 V35 0 -8.254739745977683e-19

R35_36 V35 V36 -2882.1981229471558
L35_36 V35 V36 -1.1589077755469785e-12
C35_36 V35 V36 -4.2229079841949047e-19

R35_37 V35 V37 -5008.038736473602
L35_37 V35 V37 -5.917229965813081e-12
C35_37 V35 V37 -6.176011135394796e-20

R35_38 V35 V38 -6339.592215208837
L35_38 V35 V38 -4.100293430028738e-12
C35_38 V35 V38 -1.107779099525078e-19

R35_39 V35 V39 -2656.729716523514
L35_39 V35 V39 8.505300279900519e-13
C35_39 V35 V39 8.232023710914661e-19

R35_40 V35 V40 -2721.5097100165085
L35_40 V35 V40 2.3458262975975624e-12
C35_40 V35 V40 2.9490617258427725e-19

R35_41 V35 V41 10480.372733380687
L35_41 V35 V41 4.460252446874773e-12
C35_41 V35 V41 1.166174125002973e-19

R35_42 V35 V42 252777.7492628096
L35_42 V35 V42 3.5777753606708976e-12
C35_42 V35 V42 1.7473647566207757e-19

R35_43 V35 V43 -18079.92498121572
L35_43 V35 V43 1.324390807742947e-12
C35_43 V35 V43 5.936139411277474e-19

R35_44 V35 V44 11758.915270836967
L35_44 V35 V44 5.9222351926905685e-12
C35_44 V35 V44 1.6128841424277299e-19

R35_45 V35 V45 3248.3223368670187
L35_45 V35 V45 3.896615531761588e-12
C35_45 V35 V45 3.6200882725527424e-20

R35_46 V35 V46 3511.1110510418275
L35_46 V35 V46 2.2621018730774074e-12
C35_46 V35 V46 1.6885745191582447e-19

R35_47 V35 V47 2322.243951805676
L35_47 V35 V47 -2.9525153624244913e-12
C35_47 V35 V47 -5.760519137584738e-19

R35_48 V35 V48 3105.911549803249
L35_48 V35 V48 3.1356102257063047e-12
C35_48 V35 V48 5.2409693510708185e-20

R35_49 V35 V49 15051.863168517977
L35_49 V35 V49 -5.180490554817232e-12
C35_49 V35 V49 -5.417815415136228e-20

R35_50 V35 V50 -157254.61472355385
L35_50 V35 V50 -1.720987302014011e-12
C35_50 V35 V50 -3.1756631368903667e-19

R35_51 V35 V51 2112.147119819844
L35_51 V35 V51 2.810865458791433e-12
C35_51 V35 V51 2.6809006827199267e-19

R35_52 V35 V52 -25553.932616595906
L35_52 V35 V52 -4.142887324102044e-12
C35_52 V35 V52 -1.914787377511861e-19

R35_53 V35 V53 24961.301183473937
L35_53 V35 V53 -4.7255668177052115e-12
C35_53 V35 V53 -7.875022101351535e-20

R35_54 V35 V54 -7643.755787404463
L35_54 V35 V54 -7.154044670373174e-12
C35_54 V35 V54 -1.910088538908685e-20

R35_55 V35 V55 -2450.5897971617787
L35_55 V35 V55 -1.3146811522028824e-12
C35_55 V35 V55 -2.784181197070403e-19

R35_56 V35 V56 -3437.2713777626923
L35_56 V35 V56 -3.6932427089568054e-12
C35_56 V35 V56 -5.568694124945465e-20

R35_57 V35 V57 -17960.74885777466
L35_57 V35 V57 2.687233979055679e-11
C35_57 V35 V57 5.3043068633258394e-20

R35_58 V35 V58 6220.84444353663
L35_58 V35 V58 5.3148092377084164e-12
C35_58 V35 V58 8.467838572045164e-20

R35_59 V35 V59 -2668.9966416184006
L35_59 V35 V59 3.294107003720895e-12
C35_59 V35 V59 9.678806982351722e-20

R35_60 V35 V60 -6867.1107669646035
L35_60 V35 V60 3.519060593688098e-12
C35_60 V35 V60 2.2955268441901283e-19

R35_61 V35 V61 20968.799127267004
L35_61 V35 V61 5.294375480247792e-12
C35_61 V35 V61 6.02480244682511e-20

R35_62 V35 V62 -8407.638175646893
L35_62 V35 V62 9.097257625369765e-12
C35_62 V35 V62 4.18613212431446e-20

R35_63 V35 V63 14363.188588025576
L35_63 V35 V63 5.599803053844809e-12
C35_63 V35 V63 2.5014020313132395e-19

R35_64 V35 V64 5671.707478254624
L35_64 V35 V64 -1.8810231548118843e-11
C35_64 V35 V64 -1.0700094022626384e-19

R35_65 V35 V65 5636.0796626414685
L35_65 V35 V65 1.983774942774053e-11
C35_65 V35 V65 2.1423233774118948e-20

R35_66 V35 V66 14528.805004658872
L35_66 V35 V66 -1.492508109610222e-11
C35_66 V35 V66 2.821063130635822e-21

R35_67 V35 V67 2842.519936749365
L35_67 V35 V67 -4.566271225207975e-12
C35_67 V35 V67 -1.974728688669448e-19

R35_68 V35 V68 8877.518434529602
L35_68 V35 V68 -5.458108023075813e-11
C35_68 V35 V68 -1.0265208971472201e-19

R35_69 V35 V69 35501.12871506256
L35_69 V35 V69 -4.7625658422261715e-12
C35_69 V35 V69 -8.223404903399998e-20

R35_70 V35 V70 23539.66318422176
L35_70 V35 V70 -1.467448003920144e-11
C35_70 V35 V70 -3.050271621469807e-20

R35_71 V35 V71 6331.8300575515805
L35_71 V35 V71 2.627830435584011e-12
C35_71 V35 V71 1.0215555800539816e-20

R35_72 V35 V72 12298.611067371794
L35_72 V35 V72 4.308514249365818e-12
C35_72 V35 V72 1.4533409565781275e-19

R35_73 V35 V73 8248.668945197353
L35_73 V35 V73 5.550667725788181e-12
C35_73 V35 V73 6.108526010686857e-20

R35_74 V35 V74 -10360.706824838855
L35_74 V35 V74 7.783473045133696e-12
C35_74 V35 V74 2.2578034894881887e-20

R35_75 V35 V75 -2495.790182426066
L35_75 V35 V75 -3.714185086504629e-12
C35_75 V35 V75 4.38370552469062e-20

R35_76 V35 V76 -4566.696174964568
L35_76 V35 V76 -3.2216066804612578e-12
C35_76 V35 V76 -6.218543750263258e-20

R35_77 V35 V77 -4048.7158865290057
L35_77 V35 V77 -1.0033037403031197e-11
C35_77 V35 V77 -3.1134142250153434e-21

R35_78 V35 V78 10739.351507755966
L35_78 V35 V78 -2.5074796000171744e-12
C35_78 V35 V78 -1.7729929326054913e-19

R35_79 V35 V79 -26186.629991530943
L35_79 V35 V79 -7.116986008029822e-12
C35_79 V35 V79 4.5768309873557064e-20

R35_80 V35 V80 -6889.429480222563
L35_80 V35 V80 -1.3737658454503623e-11
C35_80 V35 V80 -4.9296090284490576e-20

R35_81 V35 V81 2020.5879803947566
L35_81 V35 V81 1.0261134892572553e-11
C35_81 V35 V81 6.726956490070857e-20

R35_82 V35 V82 -12973.979785124793
L35_82 V35 V82 2.3703615871741725e-12
C35_82 V35 V82 2.3959815427902727e-19

R35_83 V35 V83 -24986.25493579968
L35_83 V35 V83 2.445420654298648e-12
C35_83 V35 V83 4.958379274295355e-20

R35_84 V35 V84 11439.802952822334
L35_84 V35 V84 2.5828031504706363e-12
C35_84 V35 V84 7.296215995870659e-20

R35_85 V35 V85 -10904.343869429846
L35_85 V35 V85 3.3360108313973855e-12
C35_85 V35 V85 1.1510460414390518e-19

R35_86 V35 V86 7270.957502223734
L35_86 V35 V86 1.6598786712579038e-12
C35_86 V35 V86 1.8784710919433086e-19

R35_87 V35 V87 -34498.95181796244
L35_87 V35 V87 -2.2089846902533777e-12
C35_87 V35 V87 -3.5571590388468156e-19

R35_88 V35 V88 13384.718648262802
L35_88 V35 V88 -5.4092204800267375e-12
C35_88 V35 V88 -4.956881776824179e-20

R35_89 V35 V89 -10758.535254134316
L35_89 V35 V89 -2.360981217701039e-12
C35_89 V35 V89 -2.307499559589587e-19

R35_90 V35 V90 -69443.8718854362
L35_90 V35 V90 -8.736995323770643e-13
C35_90 V35 V90 -5.213212265002784e-19

R35_91 V35 V91 937.5722285988538
L35_91 V35 V91 1.73931850205015e-12
C35_91 V35 V91 3.6385589847220265e-19

R35_92 V35 V92 51232.36939726783
L35_92 V35 V92 2.580100140015893e-12
C35_92 V35 V92 9.086845657506574e-20

R35_93 V35 V93 2308.2564345542874
L35_93 V35 V93 -7.283204564832416e-12
C35_93 V35 V93 -1.8212186344796825e-20

R35_94 V35 V94 -4325.129199733774
L35_94 V35 V94 -2.3961059603374233e-11
C35_94 V35 V94 8.347653665517313e-20

R35_95 V35 V95 -1174.3629596971443
L35_95 V35 V95 3.9288243703063966e-12
C35_95 V35 V95 4.186845196783399e-19

R35_96 V35 V96 -2984.521026514724
L35_96 V35 V96 -3.3629491611718244e-12
C35_96 V35 V96 3.995299082656057e-21

R35_97 V35 V97 -6127.340309852159
L35_97 V35 V97 1.7340398067764446e-12
C35_97 V35 V97 3.6186696471291714e-19

R35_98 V35 V98 5015.053765061122
L35_98 V35 V98 1.0667565394286978e-12
C35_98 V35 V98 3.665538123937616e-19

R35_99 V35 V99 -1134.972568920758
L35_99 V35 V99 -1.3658117411319574e-12
C35_99 V35 V99 -6.356149197261726e-19

R35_100 V35 V100 -20208.52997892772
L35_100 V35 V100 -3.2359048978838062e-12
C35_100 V35 V100 -1.7716461468568685e-19

R35_101 V35 V101 -6561.639784080602
L35_101 V35 V101 -1.7633421345983078e-12
C35_101 V35 V101 -2.5096609613140823e-19

R35_102 V35 V102 -88408.2083312426
L35_102 V35 V102 -3.806527930944554e-12
C35_102 V35 V102 -1.325914463246529e-19

R35_103 V35 V103 726.6680402412353
L35_103 V35 V103 -2.875581664912258e-12
C35_103 V35 V103 -4.009832080217546e-19

R35_104 V35 V104 2460.1066463862066
L35_104 V35 V104 1.5434108068774093e-12
C35_104 V35 V104 1.6646070924149645e-19

R35_105 V35 V105 1583.260841279607
L35_105 V35 V105 2.418022436441911e-11
C35_105 V35 V105 -9.317939663114339e-20

R35_106 V35 V106 -21634.15539412263
L35_106 V35 V106 -1.4273894165301777e-12
C35_106 V35 V106 -3.2856538184985535e-19

R35_107 V35 V107 -27361.489068610772
L35_107 V35 V107 1.3458485277622737e-12
C35_107 V35 V107 7.776683065962523e-19

R35_108 V35 V108 -5403.535589063347
L35_108 V35 V108 -2.4970004331669196e-12
C35_108 V35 V108 -1.1145999466836226e-19

R35_109 V35 V109 41655.316631263624
L35_109 V35 V109 1.8084368326168896e-12
C35_109 V35 V109 2.888551469478994e-19

R35_110 V35 V110 -3689.726385382157
L35_110 V35 V110 2.574248988355411e-12
C35_110 V35 V110 2.3960981950452173e-19

R35_111 V35 V111 -2206.8002962338514
L35_111 V35 V111 8.205912474814308e-13
C35_111 V35 V111 3.6616599679753394e-19

R35_112 V35 V112 -13958.771806234925
L35_112 V35 V112 1.1430901986459892e-10
C35_112 V35 V112 -9.734704989542915e-20

R35_113 V35 V113 -8263.631396606206
L35_113 V35 V113 -2.197526415511273e-12
C35_113 V35 V113 2.2955616656182572e-20

R35_114 V35 V114 -36377.28713984972
L35_114 V35 V114 1.851144085791243e-12
C35_114 V35 V114 2.936924001581006e-19

R35_115 V35 V115 -1718.809098530847
L35_115 V35 V115 -6.732417609721766e-13
C35_115 V35 V115 -8.486934795571647e-19

R35_116 V35 V116 -8145.557485123842
L35_116 V35 V116 1.54119504328956e-11
C35_116 V35 V116 1.5096120931162687e-19

R35_117 V35 V117 -1905.248331026282
L35_117 V35 V117 -3.979493527453279e-12
C35_117 V35 V117 -1.582358551772271e-19

R35_118 V35 V118 2247.712256123887
L35_118 V35 V118 -2.765387974337399e-12
C35_118 V35 V118 -2.999363808250618e-19

R35_119 V35 V119 864.7926755436332
L35_119 V35 V119 -1.3217832019331567e-12
C35_119 V35 V119 1.1889674336000404e-20

R35_120 V35 V120 2714.363409915379
L35_120 V35 V120 -4.171415387449245e-12
C35_120 V35 V120 -1.261615555926449e-19

R35_121 V35 V121 1561.7085754486725
L35_121 V35 V121 4.421768467841043e-12
C35_121 V35 V121 1.495980760310606e-20

R35_122 V35 V122 -5989.248351166539
L35_122 V35 V122 -8.271672192304668e-12
C35_122 V35 V122 1.0639731100442568e-20

R35_123 V35 V123 -5140.1152856272065
L35_123 V35 V123 4.769319871340842e-13
C35_123 V35 V123 7.836862758469104e-19

R35_124 V35 V124 -20741.896718583575
L35_124 V35 V124 2.8455291057414814e-12
C35_124 V35 V124 -5.002339921730547e-21

R35_125 V35 V125 762.5859990857324
L35_125 V35 V125 8.607880594735234e-12
C35_125 V35 V125 2.0300282848228265e-21

R35_126 V35 V126 -22890.544578764107
L35_126 V35 V126 2.1276695870331205e-12
C35_126 V35 V126 1.9421528151243328e-19

R35_127 V35 V127 -1161.5315195226792
L35_127 V35 V127 1.8380363290343405e-11
C35_127 V35 V127 -2.6470665742213242e-19

R35_128 V35 V128 -1862.5896746523924
L35_128 V35 V128 1.473721429035926e-11
C35_128 V35 V128 1.0837039151602375e-19

R35_129 V35 V129 -599.4422790665325
L35_129 V35 V129 3.4327460575427366e-11
C35_129 V35 V129 2.0043565180423833e-19

R35_130 V35 V130 -3359.383284411431
L35_130 V35 V130 -3.0257777724903744e-12
C35_130 V35 V130 -1.4407943291776069e-19

R35_131 V35 V131 1866.8673749631848
L35_131 V35 V131 -7.9587605277573e-13
C35_131 V35 V131 -3.6803836810776385e-19

R35_132 V35 V132 1418.8656696432922
L35_132 V35 V132 -1.4354704757031546e-12
C35_132 V35 V132 -2.5495478201077263e-19

R35_133 V35 V133 -1966.2082720624312
L35_133 V35 V133 -3.4025493925217864e-12
C35_133 V35 V133 -1.2239665965103952e-19

R35_134 V35 V134 1726.4184443217655
L35_134 V35 V134 -9.787503362178765e-12
C35_134 V35 V134 1.0558861261122206e-19

R35_135 V35 V135 -72789.41897160327
L35_135 V35 V135 1.1116368440549963e-12
C35_135 V35 V135 5.923188476494678e-19

R35_136 V35 V136 2677.701043648879
L35_136 V35 V136 6.105222565229759e-11
C35_136 V35 V136 3.908724604323308e-20

R35_137 V35 V137 501.7531351708844
L35_137 V35 V137 -4.661506039469582e-12
C35_137 V35 V137 -1.6641975992986785e-19

R35_138 V35 V138 -5203.357038773907
L35_138 V35 V138 2.1725062587002803e-12
C35_138 V35 V138 5.1478241624580547e-20

R35_139 V35 V139 1583.2580636411972
L35_139 V35 V139 -9.65577876954425e-13
C35_139 V35 V139 -5.42488945544174e-19

R35_140 V35 V140 -1965.3120877782528
L35_140 V35 V140 4.371962524910604e-12
C35_140 V35 V140 2.78008042843231e-20

R35_141 V35 V141 11532.323339188004
L35_141 V35 V141 1.1508085416964413e-12
C35_141 V35 V141 3.340194760595107e-19

R35_142 V35 V142 -915.554951873038
L35_142 V35 V142 4.200176803770665e-12
C35_142 V35 V142 -6.389278647791448e-20

R35_143 V35 V143 -1420.2662838793062
L35_143 V35 V143 1.2439931178018531e-12
C35_143 V35 V143 9.544442073531188e-20

R35_144 V35 V144 -6241.019842600883
L35_144 V35 V144 3.2130153100312795e-11
C35_144 V35 V144 1.645853674136148e-21

R35_145 V35 V145 -529.9310402123275
L35_145 V35 V145 2.910369980846546e-12
C35_145 V35 V145 1.5738219276434777e-19

R35_146 V35 V146 12349.757216885266
L35_146 V35 V146 -1.756249903995085e-12
C35_146 V35 V146 -7.438171301740225e-20

R35_147 V35 V147 -475.6327212430365
L35_147 V35 V147 2.774034047154655e-12
C35_147 V35 V147 4.074183898129266e-19

R35_148 V35 V148 -5305.672297304912
L35_148 V35 V148 2.6848610275634106e-12
C35_148 V35 V148 5.337898192594283e-20

R35_149 V35 V149 -5658.798438884319
L35_149 V35 V149 -5.43703763691219e-13
C35_149 V35 V149 -5.824740857710574e-19

R35_150 V35 V150 514.6087892557259
L35_150 V35 V150 1.504758743696381e-11
C35_150 V35 V150 2.302369674226173e-19

R35_151 V35 V151 234.5864628650534
L35_151 V35 V151 -1.3719100671973063e-12
C35_151 V35 V151 -2.1481809514416993e-19

R35_152 V35 V152 -76923.68437672232
L35_152 V35 V152 2.4945313183229618e-11
C35_152 V35 V152 1.6392076361119475e-20

R35_153 V35 V153 520.9192903797089
L35_153 V35 V153 -1.135194516733681e-11
C35_153 V35 V153 2.4649030582107366e-20

R35_154 V35 V154 3167.5809445948853
L35_154 V35 V154 4.922085341132349e-12
C35_154 V35 V154 -9.433343622549453e-20

R35_155 V35 V155 -233.01079234022504
L35_155 V35 V155 -1.111377522900993e-12
C35_155 V35 V155 -2.5666239277044083e-19

R35_156 V35 V156 1379.077361076715
L35_156 V35 V156 -6.425921237638397e-12
C35_156 V35 V156 -5.9675314986912e-20

R35_157 V35 V157 1153.72437235
L35_157 V35 V157 5.677664805682126e-13
C35_157 V35 V157 4.49706136151978e-19

R35_158 V35 V158 -1340.9600725096725
L35_158 V35 V158 -5.945501350871867e-12
C35_158 V35 V158 -7.809392346949098e-20

R35_159 V35 V159 -2350.8870662945233
L35_159 V35 V159 6.281054091339489e-13
C35_159 V35 V159 2.148308044796212e-19

R35_160 V35 V160 15314.299362156396
L35_160 V35 V160 -2.8093195367121457e-12
C35_160 V35 V160 -4.98458587614871e-20

R35_161 V35 V161 -1267.418759812567
L35_161 V35 V161 -2.0646637637130405e-12
C35_161 V35 V161 -5.793222849090176e-20

R35_162 V35 V162 -2668.471131770019
L35_162 V35 V162 -1.3257587250999764e-12
C35_162 V35 V162 -1.2142548462678666e-19

R35_163 V35 V163 5977.336708297739
L35_163 V35 V163 -9.243091332846493e-13
C35_163 V35 V163 -1.3359289281203153e-19

R35_164 V35 V164 239561.6789298642
L35_164 V35 V164 1.952364038653938e-11
C35_164 V35 V164 -4.328485203335633e-20

R35_165 V35 V165 -4728.412212392568
L35_165 V35 V165 -1.4916348174938026e-12
C35_165 V35 V165 -1.4024338930288548e-19

R35_166 V35 V166 1301.8124445412743
L35_166 V35 V166 2.3742904562272816e-12
C35_166 V35 V166 1.1741611772300861e-19

R35_167 V35 V167 334.11633703926407
L35_167 V35 V167 -3.985393179800165e-12
C35_167 V35 V167 7.374249301946667e-20

R35_168 V35 V168 -711.2130968423685
L35_168 V35 V168 -1.3280792968269961e-11
C35_168 V35 V168 5.451851549481576e-20

R35_169 V35 V169 1254.0433703289718
L35_169 V35 V169 2.550699657078557e-12
C35_169 V35 V169 1.0865710194691355e-19

R35_170 V35 V170 -4081.905141383905
L35_170 V35 V170 -2.960451516164903e-11
C35_170 V35 V170 -1.3673678613607692e-19

R35_171 V35 V171 -379.5588589808177
L35_171 V35 V171 1.0386559957787498e-12
C35_171 V35 V171 -7.591381470449854e-20

R35_172 V35 V172 4947.080642863277
L35_172 V35 V172 7.105253086053024e-12
C35_172 V35 V172 -4.433746113550228e-20

R35_173 V35 V173 -63006.099970450254
L35_173 V35 V173 4.021194771997626e-12
C35_173 V35 V173 -3.743770433990434e-20

R35_174 V35 V174 -1430.9202969441349
L35_174 V35 V174 -3.18979978130395e-12
C35_174 V35 V174 1.1987604345018756e-19

R35_175 V35 V175 -2060.1229604337495
L35_175 V35 V175 -9.464786098943866e-13
C35_175 V35 V175 -3.2775831068174464e-19

R35_176 V35 V176 6529.758196119825
L35_176 V35 V176 -7.220535872217236e-12
C35_176 V35 V176 -4.2028802914041013e-20

R35_177 V35 V177 3994.2927262459257
L35_177 V35 V177 -7.914025171112808e-12
C35_177 V35 V177 -1.0577869200761044e-20

R35_178 V35 V178 1181.2802121583713
L35_178 V35 V178 2.0167780564637075e-12
C35_178 V35 V178 6.227954697206879e-20

R35_179 V35 V179 3698.025192263934
L35_179 V35 V179 -3.621258676841113e-12
C35_179 V35 V179 4.294524932072705e-19

R35_180 V35 V180 2378.274073995587
L35_180 V35 V180 2.2566443602778787e-12
C35_180 V35 V180 1.4764460260093867e-19

R35_181 V35 V181 -2858.810584918272
L35_181 V35 V181 -7.2731809159526414e-12
C35_181 V35 V181 8.067567671494843e-20

R35_182 V35 V182 -2123.008695719485
L35_182 V35 V182 -2.1495546219589647e-12
C35_182 V35 V182 -1.4835809870036725e-19

R35_183 V35 V183 728.1064076337848
L35_183 V35 V183 6.505371684231448e-13
C35_183 V35 V183 3.6945672325612985e-21

R35_184 V35 V184 21343.600077976153
L35_184 V35 V184 3.808081362563869e-12
C35_184 V35 V184 3.255174834638538e-20

R35_185 V35 V185 2575.2061898100596
L35_185 V35 V185 3.648619322397931e-12
C35_185 V35 V185 -5.374038446130117e-20

R35_186 V35 V186 -1895.421778356159
L35_186 V35 V186 -1.802408606900577e-11
C35_186 V35 V186 9.8104645549456e-20

R35_187 V35 V187 -987.8759159589443
L35_187 V35 V187 -9.124720960666438e-13
C35_187 V35 V187 -3.798018482212074e-19

R35_188 V35 V188 -957.1850977366495
L35_188 V35 V188 -1.2009187522456756e-12
C35_188 V35 V188 -1.4257771401348185e-19

R35_189 V35 V189 -21750.762408659997
L35_189 V35 V189 -6.2711605524522295e-12
C35_189 V35 V189 -5.450187081614428e-20

R35_190 V35 V190 1529.177393708428
L35_190 V35 V190 9.056876989266355e-12
C35_190 V35 V190 9.092321837153429e-20

R35_191 V35 V191 -1885.95114320067
L35_191 V35 V191 -1.0872036402320279e-12
C35_191 V35 V191 1.2484199543805702e-19

R35_192 V35 V192 3471.452409384958
L35_192 V35 V192 -9.346807939063334e-12
C35_192 V35 V192 -5.66630518843484e-20

R35_193 V35 V193 -2569.7662606019558
L35_193 V35 V193 -4.89246075445455e-12
C35_193 V35 V193 6.306421971731224e-20

R35_194 V35 V194 5648.493544292021
L35_194 V35 V194 3.997271289336613e-12
C35_194 V35 V194 6.736479646022375e-20

R35_195 V35 V195 971.2978749636522
L35_195 V35 V195 7.56668452461345e-13
C35_195 V35 V195 -7.578383423857352e-20

R35_196 V35 V196 752.6000545345224
L35_196 V35 V196 1.290880526173194e-12
C35_196 V35 V196 2.6068456274280065e-19

R35_197 V35 V197 2839.5626530329
L35_197 V35 V197 3.4337752383375575e-12
C35_197 V35 V197 4.167818566485815e-20

R35_198 V35 V198 -5474.984662330085
L35_198 V35 V198 -7.807461805198003e-12
C35_198 V35 V198 -3.7494200608253923e-20

R35_199 V35 V199 -3339.4077700125667
L35_199 V35 V199 2.7081279726597357e-11
C35_199 V35 V199 -2.6636633576391327e-21

R35_200 V35 V200 -1166.4553187945908
L35_200 V35 V200 -1.2213074571867954e-11
C35_200 V35 V200 -5.842970563637187e-20

R36_36 V36 0 -130.6989335961353
L36_36 V36 0 -2.3663519106601297e-13
C36_36 V36 0 -2.2295232535551413e-18

R36_37 V36 V37 -3289.1229648967696
L36_37 V36 V37 -3.1927205743124934e-12
C36_37 V36 V37 -1.0056343606647228e-19

R36_38 V36 V38 -3776.4052626981734
L36_38 V36 V38 -2.922281236182002e-12
C36_38 V36 V38 -1.819721943004664e-19

R36_39 V36 V39 -2311.1979287942445
L36_39 V36 V39 3.8678492535145784e-12
C36_39 V36 V39 2.4532322502132155e-19

R36_40 V36 V40 -1186.539297586889
L36_40 V36 V40 7.38845652168394e-13
C36_40 V36 V40 1.0645154830852018e-18

R36_41 V36 V41 6286.665700048021
L36_41 V36 V41 3.4279802295557354e-12
C36_41 V36 V41 2.15555985190348e-19

R36_42 V36 V42 41411.81100186107
L36_42 V36 V42 2.5769596582124924e-12
C36_42 V36 V42 3.05806823128436e-19

R36_43 V36 V43 14907.150557034207
L36_43 V36 V43 3.094093668102695e-11
C36_43 V36 V43 6.413006574126593e-20

R36_44 V36 V44 -47065.650346134425
L36_44 V36 V44 9.420254709796972e-13
C36_44 V36 V44 6.616182286944358e-19

R36_45 V36 V45 2098.5582913854805
L36_45 V36 V45 2.065198283733029e-12
C36_45 V36 V45 1.5531454923105867e-19

R36_46 V36 V46 2170.9286197957076
L36_46 V36 V46 1.5039300492667689e-12
C36_46 V36 V46 3.6691095014531017e-19

R36_47 V36 V47 2494.942551951636
L36_47 V36 V47 4.316119144731631e-12
C36_47 V36 V47 3.71135492808053e-20

R36_48 V36 V48 1030.0695919652544
L36_48 V36 V48 1.3709464046891001e-11
C36_48 V36 V48 -3.5606602590901377e-19

R36_49 V36 V49 10516.697980453298
L36_49 V36 V49 -4.322693965270913e-12
C36_49 V36 V49 -6.578120867218561e-20

R36_50 V36 V50 -53568.226646718664
L36_50 V36 V50 -1.4554965422114903e-12
C36_50 V36 V50 -4.018618755291398e-19

R36_51 V36 V51 12038.712518100027
L36_51 V36 V51 -3.772192982264541e-12
C36_51 V36 V51 -2.0207524125269097e-19

R36_52 V36 V52 3020.1196829843593
L36_52 V36 V52 5.156148742088206e-12
C36_52 V36 V52 1.0647199497964304e-19

R36_53 V36 V53 12932.793830036031
L36_53 V36 V53 -3.3605989433666664e-12
C36_53 V36 V53 -1.7608392040365991e-19

R36_54 V36 V54 -4420.82502920845
L36_54 V36 V54 -3.3952931388607937e-12
C36_54 V36 V54 -1.48397088687027e-19

R36_55 V36 V55 -7874.517249435911
L36_55 V36 V55 -7.749942484211907e-12
C36_55 V36 V55 -4.400481678196471e-20

R36_56 V36 V56 -1034.9415753887963
L36_56 V36 V56 -7.093322204385929e-13
C36_56 V36 V56 -6.763092301761548e-19

R36_57 V36 V57 -11958.960195416324
L36_57 V36 V57 -3.9622098607514485e-10
C36_57 V36 V57 1.6803330844290845e-19

R36_58 V36 V58 3547.8871136909956
L36_58 V36 V58 3.0245704936883233e-12
C36_58 V36 V58 2.4201326966739083e-19

R36_59 V36 V59 -6440.610419000954
L36_59 V36 V59 2.4902391650369585e-12
C36_59 V36 V59 3.7572201266333745e-19

R36_60 V36 V60 -1518.693135191897
L36_60 V36 V60 1.913471962405622e-12
C36_60 V36 V60 2.924328300016439e-19

R36_61 V36 V61 10662.092507836434
L36_61 V36 V61 3.2742703582378696e-12
C36_61 V36 V61 9.016469300435144e-20

R36_62 V36 V62 -6048.977577090126
L36_62 V36 V62 4.9144246734580496e-12
C36_62 V36 V62 1.4529345140889076e-19

R36_63 V36 V63 10905.31108264539
L36_63 V36 V63 -3.784203065772199e-12
C36_63 V36 V63 -1.860251532768966e-19

R36_64 V36 V64 2209.2599020476246
L36_64 V36 V64 2.7483561413902163e-12
C36_64 V36 V64 2.2867481510347167e-19

R36_65 V36 V65 3786.8840485461355
L36_65 V36 V65 7.596838440596469e-12
C36_65 V36 V65 9.217455669053635e-20

R36_66 V36 V66 12356.717263447132
L36_66 V36 V66 -8.596195435686401e-12
C36_66 V36 V66 -1.4412113662271935e-20

R36_67 V36 V67 -14527.216711978386
L36_67 V36 V67 -2.9554854309228197e-12
C36_67 V36 V67 -2.1355232816209939e-19

R36_68 V36 V68 1800.6279377331555
L36_68 V36 V68 -1.4350071068854861e-11
C36_68 V36 V68 -1.1283169789589713e-19

R36_69 V36 V69 -28711.076225180255
L36_69 V36 V69 -3.045310430819751e-12
C36_69 V36 V69 -2.3763182651035728e-19

R36_70 V36 V70 24301.323780027662
L36_70 V36 V70 -8.305171080778104e-12
C36_70 V36 V70 -1.4153391337164148e-19

R36_71 V36 V71 5154.483514766683
L36_71 V36 V71 1.7499602922968661e-12
C36_71 V36 V71 2.731705292266756e-19

R36_72 V36 V72 4559.374596231692
L36_72 V36 V72 2.1923238243773966e-12
C36_72 V36 V72 -5.600654957205722e-21

R36_73 V36 V73 4302.783625631483
L36_73 V36 V73 3.6010976478713274e-12
C36_73 V36 V73 1.544141777186495e-19

R36_74 V36 V74 -7009.846625511266
L36_74 V36 V74 5.3893743533048396e-12
C36_74 V36 V74 1.12871362391494e-19

R36_75 V36 V75 8059.805861463896
L36_75 V36 V75 6.160881779889512e-12
C36_75 V36 V75 1.2831380489965574e-19

R36_76 V36 V76 -860.5061104391656
L36_76 V36 V76 -8.359562876989871e-13
C36_76 V36 V76 -4.2748508997452514e-19

R36_77 V36 V77 -3354.6628607203825
L36_77 V36 V77 -6.284702328431853e-12
C36_77 V36 V77 5.2545482567924754e-20

R36_78 V36 V78 4283.1876631059
L36_78 V36 V78 -2.1305142349544757e-12
C36_78 V36 V78 -3.047317422033647e-19

R36_79 V36 V79 -2268.41462765954
L36_79 V36 V79 -1.8158553518863396e-12
C36_79 V36 V79 -2.2832217276512024e-19

R36_80 V36 V80 2382.417595075579
L36_80 V36 V80 1.739144299237028e-12
C36_80 V36 V80 3.6921868862926575e-19

R36_81 V36 V81 1331.2316324407523
L36_81 V36 V81 3.4820019304354763e-12
C36_81 V36 V81 1.4768776219163883e-19

R36_82 V36 V82 -6622.857053960303
L36_82 V36 V82 1.8070738454498443e-12
C36_82 V36 V82 3.89169936432628e-19

R36_83 V36 V83 23671.603075578892
L36_83 V36 V83 6.733714749042655e-12
C36_83 V36 V83 4.29409476199187e-20

R36_84 V36 V84 8265.767023760736
L36_84 V36 V84 1.1776541877443108e-12
C36_84 V36 V84 2.605130452833082e-19

R36_85 V36 V85 -8649.508288918825
L36_85 V36 V85 2.5256478015939623e-12
C36_85 V36 V85 1.7678823766102402e-19

R36_86 V36 V86 4721.2472833739475
L36_86 V36 V86 1.3650631882040469e-12
C36_86 V36 V86 3.3337678006335277e-19

R36_87 V36 V87 9091.051274851548
L36_87 V36 V87 -1.3893607861706512e-11
C36_87 V36 V87 -9.33685014267019e-20

R36_88 V36 V88 -5578.349692329396
L36_88 V36 V88 -1.201610408872712e-12
C36_88 V36 V88 -6.683524445978049e-19

R36_89 V36 V89 -4600.230160261426
L36_89 V36 V89 -1.386908475159989e-12
C36_89 V36 V89 -4.621766266420192e-19

R36_90 V36 V90 -9296.200593688583
L36_90 V36 V90 -6.304373412679038e-13
C36_90 V36 V90 -8.948583991506884e-19

R36_91 V36 V91 2162.2323057445487
L36_91 V36 V91 1.4404213699357507e-12
C36_91 V36 V91 3.4421918330943946e-19

R36_92 V36 V92 937.1503411482836
L36_92 V36 V92 2.3273177634593495e-12
C36_92 V36 V92 3.6202300301382327e-19

R36_93 V36 V93 1633.2773047548378
L36_93 V36 V93 -1.1160929309836838e-11
C36_93 V36 V93 1.4014042839829926e-20

R36_94 V36 V94 -2715.050596982334
L36_94 V36 V94 1.654268944025222e-11
C36_94 V36 V94 2.138896867735117e-19

R36_95 V36 V95 -2356.713061504878
L36_95 V36 V95 -4.7331533436899914e-12
C36_95 V36 V95 4.380228910054328e-20

R36_96 V36 V96 -701.6699376501117
L36_96 V36 V96 4.122584490407402e-11
C36_96 V36 V96 5.24652728422318e-19

R36_97 V36 V97 -6050.190102798099
L36_97 V36 V97 1.2385102715061081e-12
C36_97 V36 V97 7.228179154031714e-19

R36_98 V36 V98 2074.380761874328
L36_98 V36 V98 8.040846318367862e-13
C36_98 V36 V98 6.181080400497134e-19

R36_99 V36 V99 -2287.2579078294393
L36_99 V36 V99 -1.0986638368647401e-12
C36_99 V36 V99 -5.195949767027269e-19

R36_100 V36 V100 -2473.2725507146206
L36_100 V36 V100 -3.3903115980654665e-11
C36_100 V36 V100 -6.815513266754138e-19

R36_101 V36 V101 -4727.824513794116
L36_101 V36 V101 -1.548462345375089e-12
C36_101 V36 V101 -3.5962008793806445e-19

R36_102 V36 V102 111909.66454094237
L36_102 V36 V102 -2.14593544157004e-12
C36_102 V36 V102 -3.087928182698522e-19

R36_103 V36 V103 1820.1992420169388
L36_103 V36 V103 1.5938807598522194e-12
C36_103 V36 V103 2.3852672126327847e-19

R36_104 V36 V104 687.9060820419353
L36_104 V36 V104 -4.415367556247179e-12
C36_104 V36 V104 -2.821225279378181e-19

R36_105 V36 V105 1165.5629001780087
L36_105 V36 V105 -8.654943147123359e-11
C36_105 V36 V105 -2.456491204302782e-19

R36_106 V36 V106 -7292.8912701644
L36_106 V36 V106 -1.2848769106955424e-12
C36_106 V36 V106 -4.6104206959158535e-19

R36_107 V36 V107 15759.628606424934
L36_107 V36 V107 2.7680961132903764e-12
C36_107 V36 V107 2.866076552758545e-19

R36_108 V36 V108 -3178.5345602529055
L36_108 V36 V108 -1.710571026335999e-11
C36_108 V36 V108 5.345951473244914e-19

R36_109 V36 V109 -12978.63453387261
L36_109 V36 V109 1.702153887007746e-12
C36_109 V36 V109 5.099948500888608e-19

R36_110 V36 V110 -2610.9818699908196
L36_110 V36 V110 2.9601742201412565e-12
C36_110 V36 V110 2.748383531180382e-19

R36_111 V36 V111 -11140.15662798717
L36_111 V36 V111 -9.653426350699726e-12
C36_111 V36 V111 -1.2923833373814319e-19

R36_112 V36 V112 -2717.761976910945
L36_112 V36 V112 6.361413104811821e-13
C36_112 V36 V112 6.106200114895176e-19

R36_113 V36 V113 74230.58495648426
L36_113 V36 V113 -2.834519049107944e-12
C36_113 V36 V113 8.781516306181593e-20

R36_114 V36 V114 169403.76363872067
L36_114 V36 V114 1.4193503689740733e-12
C36_114 V36 V114 4.656819130763836e-19

R36_115 V36 V115 -1667.4687851292063
L36_115 V36 V115 -2.2626485692100845e-12
C36_115 V36 V115 -1.217964968940142e-19

R36_116 V36 V116 -1226.5829182978673
L36_116 V36 V116 -8.983460852910443e-13
C36_116 V36 V116 -7.533035307431187e-19

R36_117 V36 V117 -1254.463612415937
L36_117 V36 V117 -2.623865037170651e-12
C36_117 V36 V117 -2.8266637949214165e-19

R36_118 V36 V118 1779.2571942811824
L36_118 V36 V118 -2.141417205941451e-12
C36_118 V36 V118 -5.370904565727873e-19

R36_119 V36 V119 1669.2330999912638
L36_119 V36 V119 -9.483943682683949e-12
C36_119 V36 V119 -2.0370747340126563e-19

R36_120 V36 V120 488.27375052745066
L36_120 V36 V120 -7.950741754204303e-13
C36_120 V36 V120 -4.567798376397972e-19

R36_121 V36 V121 1226.2732986628491
L36_121 V36 V121 6.382366331603996e-12
C36_121 V36 V121 5.76257873732082e-20

R36_122 V36 V122 -8594.131869234881
L36_122 V36 V122 -4.316310040057228e-12
C36_122 V36 V122 7.408486629379774e-21

R36_123 V36 V123 9924.961812166108
L36_123 V36 V123 3.181646566942721e-12
C36_123 V36 V123 1.7344122134950782e-19

R36_124 V36 V124 -1372.3215033975177
L36_124 V36 V124 3.831152223020406e-13
C36_124 V36 V124 1.425203409949481e-18

R36_125 V36 V125 516.3504002246681
L36_125 V36 V125 5.061651109801725e-12
C36_125 V36 V125 1.5203624585153046e-20

R36_126 V36 V126 18092.537025595277
L36_126 V36 V126 1.8038869164901645e-12
C36_126 V36 V126 3.145892885151921e-19

R36_127 V36 V127 -1677.9137305932063
L36_127 V36 V127 1.0029225146795076e-11
C36_127 V36 V127 2.265696876442437e-19

R36_128 V36 V128 -657.2157220298094
L36_128 V36 V128 1.6364303457656956e-11
C36_128 V36 V128 -2.417498736410628e-19

R36_129 V36 V129 -416.04223542659486
L36_129 V36 V129 8.073465406138295e-12
C36_129 V36 V129 3.3434629218200083e-19

R36_130 V36 V130 -1656.809126506977
L36_130 V36 V130 -2.3654427705266065e-12
C36_130 V36 V130 -2.9995393594263276e-19

R36_131 V36 V131 1269.4972648102805
L36_131 V36 V131 -5.1388880419583995e-12
C36_131 V36 V131 -2.9274161051020086e-19

R36_132 V36 V132 646.0008719744447
L36_132 V36 V132 -5.041471502158648e-13
C36_132 V36 V132 -8.658339720936288e-19

R36_133 V36 V133 -1772.479474743949
L36_133 V36 V133 -1.9905259918648658e-12
C36_133 V36 V133 -3.414284208925458e-19

R36_134 V36 V134 979.6271154915111
L36_134 V36 V134 -4.2225006152428855e-12
C36_134 V36 V134 -7.112910627420861e-20

R36_135 V36 V135 13197.096248508826
L36_135 V36 V135 -3.705587418105737e-12
C36_135 V36 V135 -7.567692118451748e-20

R36_136 V36 V136 8343.832782131305
L36_136 V36 V136 1.0250812720526024e-12
C36_136 V36 V136 1.0315280929061584e-18

R36_137 V36 V137 403.85634468757746
L36_137 V36 V137 -3.246592719086515e-12
C36_137 V36 V137 -1.2781713131697499e-19

R36_138 V36 V138 -2181.005886007441
L36_138 V36 V138 1.6117491911326487e-12
C36_138 V36 V138 2.2745839841573576e-19

R36_139 V36 V139 -1185.6297899703504
L36_139 V36 V139 1.291666674706774e-11
C36_139 V36 V139 4.2468426183890695e-20

R36_140 V36 V140 954.5424888298857
L36_140 V36 V140 -2.8988709192277873e-12
C36_140 V36 V140 -8.692506174267003e-19

R36_141 V36 V141 5625.191015803636
L36_141 V36 V141 9.03267602797714e-13
C36_141 V36 V141 5.383566542191267e-19

R36_142 V36 V142 -662.3013533079347
L36_142 V36 V142 3.2997714716530837e-12
C36_142 V36 V142 -2.2095568270768325e-20

R36_143 V36 V143 2727.569429458128
L36_143 V36 V143 2.5371921697355326e-12
C36_143 V36 V143 1.3382189972675597e-19

R36_144 V36 V144 -329.40693958865796
L36_144 V36 V144 1.147318621913474e-11
C36_144 V36 V144 6.708772285107462e-20

R36_145 V36 V145 -420.9039684615137
L36_145 V36 V145 2.143560060510917e-12
C36_145 V36 V145 1.2416774538091186e-19

R36_146 V36 V146 -8198.484304781821
L36_146 V36 V146 -1.1832485400472437e-12
C36_146 V36 V146 -1.951880148009458e-19

R36_147 V36 V147 -768.8169868983779
L36_147 V36 V147 5.97720716728282e-12
C36_147 V36 V147 1.7883034253385447e-19

R36_148 V36 V148 360.32957724830896
L36_148 V36 V148 7.143708335247448e-13
C36_148 V36 V148 6.990906143359913e-19

R36_149 V36 V149 -2065.278292607543
L36_149 V36 V149 -4.583400082049688e-13
C36_149 V36 V149 -7.1772506218115405e-19

R36_150 V36 V150 360.88067153863756
L36_150 V36 V150 4.214124292630485e-12
C36_150 V36 V150 4.346718539802155e-19

R36_151 V36 V151 814.7830090846013
L36_151 V36 V151 -3.011857238681431e-11
C36_151 V36 V151 -1.0278503513189646e-19

R36_152 V36 V152 -11796.824245869228
L36_152 V36 V152 -7.58117937286605e-13
C36_152 V36 V152 -1.9917040985528136e-19

R36_153 V36 V153 438.4205302986432
L36_153 V36 V153 -2.9040112948783846e-12
C36_153 V36 V153 -5.036010018132706e-20

R36_154 V36 V154 -4232.017757994195
L36_154 V36 V154 9.511220326692116e-12
C36_154 V36 V154 -1.3322344384465386e-19

R36_155 V36 V155 -441.899363138803
L36_155 V36 V155 -1.4728227425903487e-12
C36_155 V36 V155 -1.957236376431472e-19

R36_156 V36 V156 319.3842300965524
L36_156 V36 V156 2.5367736589536194e-12
C36_156 V36 V156 -4.809058433789446e-19

R36_157 V36 V157 528.0684420257043
L36_157 V36 V157 4.0240308468822473e-13
C36_157 V36 V157 8.482375228065554e-19

R36_158 V36 V158 -2392.4873520105375
L36_158 V36 V158 -2.941673882781914e-10
C36_158 V36 V158 -8.89018435727669e-20

R36_159 V36 V159 415.67757736383214
L36_159 V36 V159 5.866368534614149e-11
C36_159 V36 V159 1.8117349275297607e-20

R36_160 V36 V160 -217.4525695025881
L36_160 V36 V160 1.5025633235603944e-12
C36_160 V36 V160 2.268873443042747e-19

R36_161 V36 V161 -730.9883254943128
L36_161 V36 V161 -1.689413522158811e-12
C36_161 V36 V161 -1.6013658482211865e-19

R36_162 V36 V162 -1953.7124673013584
L36_162 V36 V162 -1.0437173173002183e-12
C36_162 V36 V162 -1.3766524718398595e-19

R36_163 V36 V163 -4305.721433035158
L36_163 V36 V163 1.3063647325135828e-11
C36_163 V36 V163 1.0786670708343021e-19

R36_164 V36 V164 460.0140057820959
L36_164 V36 V164 -1.3046356970035489e-12
C36_164 V36 V164 -2.5362043313226214e-19

R36_165 V36 V165 2284.6890416548094
L36_165 V36 V165 -1.4948918806133805e-12
C36_165 V36 V165 -1.5823893469872733e-19

R36_166 V36 V166 657.853471267898
L36_166 V36 V166 1.4768897131670887e-12
C36_166 V36 V166 2.783041157517173e-19

R36_167 V36 V167 3984.6848947629082
L36_167 V36 V167 2.965456087505018e-12
C36_167 V36 V167 -3.43038981071181e-20

R36_168 V36 V168 -57288.46627980372
L36_168 V36 V168 -1.347415174226037e-12
C36_168 V36 V168 1.4542104623811665e-19

R36_169 V36 V169 1071.2661319095018
L36_169 V36 V169 3.0643470990139546e-12
C36_169 V36 V169 2.7991307899317575e-19

R36_170 V36 V170 -2046.4513996988696
L36_170 V36 V170 -1.3313535483493534e-11
C36_170 V36 V170 -2.1164858465489628e-19

R36_171 V36 V171 -1091.0329424700444
L36_171 V36 V171 -1.6542203279439511e-12
C36_171 V36 V171 -1.6087043771915088e-19

R36_172 V36 V172 -1230.0531960378814
L36_172 V36 V172 5.404429455630946e-13
C36_172 V36 V172 -4.74140902590242e-20

R36_173 V36 V173 -10931.707352144216
L36_173 V36 V173 2.6300640418651837e-12
C36_173 V36 V173 -1.0190034540676016e-19

R36_174 V36 V174 -803.023619878935
L36_174 V36 V174 -2.0490089613097955e-12
C36_174 V36 V174 1.7243562261036278e-19

R36_175 V36 V175 1448.8150752907861
L36_175 V36 V175 -5.868478506254661e-10
C36_175 V36 V175 -6.143368605322646e-20

R36_176 V36 V176 -1851.5684982365412
L36_176 V36 V176 -6.700884207311437e-13
C36_176 V36 V176 -5.584252168954522e-19

R36_177 V36 V177 2560.9079793324454
L36_177 V36 V177 -1.2762413728041207e-11
C36_177 V36 V177 -1.4742474648886941e-21

R36_178 V36 V178 843.41192710596
L36_178 V36 V178 1.4985004617147966e-12
C36_178 V36 V178 7.774890262140821e-20

R36_179 V36 V179 -2774.9900706001554
L36_179 V36 V179 1.0634499167269804e-12
C36_179 V36 V179 3.0145676414119336e-19

R36_180 V36 V180 944.0941088140861
L36_180 V36 V180 -2.3805363933822116e-12
C36_180 V36 V180 6.229117324169094e-19

R36_181 V36 V181 -1864.2833227898866
L36_181 V36 V181 -9.045469299669626e-12
C36_181 V36 V181 1.1860055682080052e-19

R36_182 V36 V182 -1514.1644566341745
L36_182 V36 V182 -2.7349680761061353e-12
C36_182 V36 V182 -1.3681944720569137e-19

R36_183 V36 V183 1611.3009827849164
L36_183 V36 V183 3.5017162688658754e-12
C36_183 V36 V183 1.3272271088557336e-19

R36_184 V36 V184 1325.4682112798864
L36_184 V36 V184 5.491344781999708e-13
C36_184 V36 V184 -1.31775899720505e-19

R36_185 V36 V185 1430.4926988264779
L36_185 V36 V185 2.050497184724839e-12
C36_185 V36 V185 -7.779921743901845e-20

R36_186 V36 V186 -3923.6038783427725
L36_186 V36 V186 5.958080023354737e-12
C36_186 V36 V186 2.4769027872640775e-20

R36_187 V36 V187 -6183.719657996978
L36_187 V36 V187 -1.7041525691269878e-12
C36_187 V36 V187 -3.480845100569557e-19

R36_188 V36 V188 -334.39574555077115
L36_188 V36 V188 -5.004779502908386e-13
C36_188 V36 V188 -3.449599260635531e-19

R36_189 V36 V189 -9131.181105144191
L36_189 V36 V189 -3.5249252094811947e-12
C36_189 V36 V189 -7.178212620140821e-20

R36_190 V36 V190 1054.2240620761672
L36_190 V36 V190 7.553134030562293e-11
C36_190 V36 V190 1.7192734826648063e-19

R36_191 V36 V191 -2751.888729792328
L36_191 V36 V191 -1.3090454997981928e-12
C36_191 V36 V191 -1.3590558487465162e-19

R36_192 V36 V192 1734.3457514753297
L36_192 V36 V192 -2.3389689207543105e-09
C36_192 V36 V192 2.8279444292872376e-19

R36_193 V36 V193 -1117.4987249213234
L36_193 V36 V193 -2.949704512335197e-12
C36_193 V36 V193 1.4493240955295954e-19

R36_194 V36 V194 3096.9218055585957
L36_194 V36 V194 2.003254183773142e-12
C36_194 V36 V194 3.0837306795060023e-19

R36_195 V36 V195 1028.3370373374069
L36_195 V36 V195 7.098339357914683e-13
C36_195 V36 V195 5.41963199655155e-19

R36_196 V36 V196 539.9331930817083
L36_196 V36 V196 1.8214746345143976e-12
C36_196 V36 V196 -4.2646528279586997e-19

R36_197 V36 V197 4261.654470621445
L36_197 V36 V197 2.0764947009679213e-12
C36_197 V36 V197 -2.5350495805613454e-20

R36_198 V36 V198 10968.600085790567
L36_198 V36 V198 -1.1375791062886586e-11
C36_198 V36 V198 3.816918903976887e-20

R36_199 V36 V199 1073.5955613351662
L36_199 V36 V199 3.477815443794518e-11
C36_199 V36 V199 2.8838760619228697e-20

R36_200 V36 V200 -470.5188889304538
L36_200 V36 V200 4.2549077314392254e-12
C36_200 V36 V200 7.34770288462731e-20

R37_37 V37 0 -174.91739972726245
L37_37 V37 0 -1.600037429134001e-13
C37_37 V37 0 -1.187642367984967e-18

R37_38 V37 V38 -6143.818971412955
L37_38 V37 V38 -1.5163436824303046e-12
C37_38 V37 V38 -3.2537854370508597e-19

R37_39 V37 V39 -5029.212718100803
L37_39 V37 V39 -2.293812453936719e-12
C37_39 V37 V39 -1.8551009798570122e-19

R37_40 V37 V40 -3085.0404021099366
L37_40 V37 V40 -1.657725956010663e-12
C37_40 V37 V40 -2.5153307755542045e-19

R37_41 V37 V41 16730.11834955367
L37_41 V37 V41 2.805744026883218e-12
C37_41 V37 V41 5.632870803762919e-19

R37_42 V37 V42 -34230.58313136237
L37_42 V37 V42 1.8269644867301638e-11
C37_42 V37 V42 1.5331668320774484e-19

R37_43 V37 V43 -11808.463294431394
L37_43 V37 V43 -1.520357233943236e-11
C37_43 V37 V43 1.1289898262005747e-19

R37_44 V37 V44 -10694.144326654123
L37_44 V37 V44 7.553413869447868e-11
C37_44 V37 V44 2.0275840035631055e-19

R37_45 V37 V45 993.1358449474101
L37_45 V37 V45 6.594522130227724e-13
C37_45 V37 V45 6.572103279350283e-19

R37_46 V37 V46 19960.862962860985
L37_46 V37 V46 3.747341377291606e-12
C37_46 V37 V46 1.3343601394306683e-19

R37_47 V37 V47 19570.18540403958
L37_47 V37 V47 3.798124679841197e-12
C37_47 V37 V47 9.578074711578779e-20

R37_48 V37 V48 4766.275504744169
L37_48 V37 V48 1.9164862810498895e-12
C37_48 V37 V48 1.9582330836804406e-19

R37_49 V37 V49 1415.6855703161395
L37_49 V37 V49 -1.655904815918842e-12
C37_49 V37 V49 -5.0932304081349e-19

R37_50 V37 V50 -14657.642994274556
L37_50 V37 V50 -1.0325956491846358e-11
C37_50 V37 V50 -7.341741071903097e-20

R37_51 V37 V51 55464.27145877299
L37_51 V37 V51 5.869614533552557e-12
C37_51 V37 V51 2.315389085415955e-20

R37_52 V37 V52 -16998.03360048745
L37_52 V37 V52 2.5258942461090337e-11
C37_52 V37 V52 -3.668143099443707e-20

R37_53 V37 V53 5192.859592536132
L37_53 V37 V53 1.343516107812639e-12
C37_53 V37 V53 1.1536510254775112e-19

R37_54 V37 V54 102454.52303626252
L37_54 V37 V54 2.7229163932529034e-11
C37_54 V37 V54 -6.23328392824641e-20

R37_55 V37 V55 18490.294049434688
L37_55 V37 V55 1.5135391336478407e-11
C37_55 V37 V55 -3.5535169864993294e-20

R37_56 V37 V56 -12654.79126269907
L37_56 V37 V56 -7.572893380438751e-12
C37_56 V37 V56 -1.216612548534085e-19

R37_57 V37 V57 -6280.770716072963
L37_57 V37 V57 -8.919003973750447e-13
C37_57 V37 V57 -5.337515441925607e-19

R37_58 V37 V58 -9244.990996185115
L37_58 V37 V58 -5.255866759776704e-12
C37_58 V37 V58 -2.0790698146892643e-20

R37_59 V37 V59 -3798.7698988055477
L37_59 V37 V59 -2.8895872965845612e-12
C37_59 V37 V59 -8.011829445475944e-20

R37_60 V37 V60 -2579.6742591208217
L37_60 V37 V60 -1.9660250451473036e-12
C37_60 V37 V60 -1.0977963443439455e-19

R37_61 V37 V61 -58925.39710939807
L37_61 V37 V61 1.7396485382604245e-12
C37_61 V37 V61 4.1862951270962845e-19

R37_62 V37 V62 -79531.69131767443
L37_62 V37 V62 -7.867547936707375e-12
C37_62 V37 V62 -6.292408741475088e-20

R37_63 V37 V63 -329771.6794986436
L37_63 V37 V63 -4.8967651954260176e-12
C37_63 V37 V63 -5.770481432095572e-20

R37_64 V37 V64 9335.313781786728
L37_64 V37 V64 -5.123562243736987e-11
C37_64 V37 V64 1.949470323876461e-20

R37_65 V37 V65 1391.7809949288305
L37_65 V37 V65 2.2256744426115936e-12
C37_65 V37 V65 3.731705257888078e-19

R37_66 V37 V66 -18784.492908573862
L37_66 V37 V66 7.924280406172589e-12
C37_66 V37 V66 9.416770817890733e-20

R37_67 V37 V67 -29623.22432550839
L37_67 V37 V67 4.320480450419043e-12
C37_67 V37 V67 1.154312970247851e-19

R37_68 V37 V68 11985.639263635587
L37_68 V37 V68 1.6855804000352087e-12
C37_68 V37 V68 2.8577278674152283e-19

R37_69 V37 V69 2223.274364451909
L37_69 V37 V69 4.860178303565337e-10
C37_69 V37 V69 -3.731590515624458e-19

R37_70 V37 V70 -12218.617123426982
L37_70 V37 V70 9.587728385260483e-12
C37_70 V37 V70 5.2559158240387637e-20

R37_71 V37 V71 -31919.874575904483
L37_71 V37 V71 4.163288406006204e-12
C37_71 V37 V71 8.06304314036382e-20

R37_72 V37 V72 -14036.32518686896
L37_72 V37 V72 7.5647698874041e-12
C37_72 V37 V72 -1.213205986526664e-20

R37_73 V37 V73 -5157.264430779551
L37_73 V37 V73 3.4432388485131327e-12
C37_73 V37 V73 1.4598438856256279e-19

R37_74 V37 V74 -28952.721517029113
L37_74 V37 V74 -2.7361656780265407e-12
C37_74 V37 V74 -2.299431630222217e-19

R37_75 V37 V75 13247.716383983689
L37_75 V37 V75 -3.5581667788086834e-12
C37_75 V37 V75 -9.21929163624421e-20

R37_76 V37 V76 -7125.621232691521
L37_76 V37 V76 -1.4070071618317405e-12
C37_76 V37 V76 -2.7587136663048265e-19

R37_77 V37 V77 -2866.551986721994
L37_77 V37 V77 -1.7731991009543304e-12
C37_77 V37 V77 -2.601659062238698e-19

R37_78 V37 V78 3415.1070058030355
L37_78 V37 V78 3.425885032639465e-12
C37_78 V37 V78 1.4399619966310666e-19

R37_79 V37 V79 17779.950838061704
L37_79 V37 V79 -1.0760940876686261e-10
C37_79 V37 V79 -5.729047387920558e-20

R37_80 V37 V80 5742.032962004239
L37_80 V37 V80 3.793131598567495e-12
C37_80 V37 V80 7.479027936914732e-20

R37_81 V37 V81 573.5768217685167
L37_81 V37 V81 1.839884501396013e-12
C37_81 V37 V81 1.3170924903414854e-19

R37_82 V37 V82 -3568.70284603136
L37_82 V37 V82 1.5530770002037044e-11
C37_82 V37 V82 2.7537298667342113e-20

R37_83 V37 V83 -2162.009325931092
L37_83 V37 V83 -7.660015472111481e-12
C37_83 V37 V83 -2.5210958333303366e-20

R37_84 V37 V84 -2990.918757201244
L37_84 V37 V84 1.0267267298573717e-11
C37_84 V37 V84 1.1871280600969618e-19

R37_85 V37 V85 52600.1376924746
L37_85 V37 V85 1.6133438861407804e-12
C37_85 V37 V85 4.929620591588097e-19

R37_86 V37 V86 -1414.0773106556103
L37_86 V37 V86 -6.515459564552313e-12
C37_86 V37 V86 1.7941477278861995e-20

R37_87 V37 V87 -7366.355740859894
L37_87 V37 V87 -9.752689671296699e-12
C37_87 V37 V87 -1.2737102940014042e-20

R37_88 V37 V88 -5063.59063134883
L37_88 V37 V88 -7.45420123852745e-12
C37_88 V37 V88 -4.120066788429472e-20

R37_89 V37 V89 -2386.443709157386
L37_89 V37 V89 1.6616355759225753e-11
C37_89 V37 V89 -1.223206931640456e-19

R37_90 V37 V90 1855.2469687840974
L37_90 V37 V90 -3.1229335483525615e-12
C37_90 V37 V90 -1.5360866706134933e-19

R37_91 V37 V91 1869.6649623141489
L37_91 V37 V91 1.6086002596955606e-12
C37_91 V37 V91 2.713338004603961e-19

R37_92 V37 V92 3400.947002700304
L37_92 V37 V92 2.5703437479285013e-12
C37_92 V37 V92 1.1710245481746462e-19

R37_93 V37 V93 964.9770660378144
L37_93 V37 V93 -1.7429720580155877e-12
C37_93 V37 V93 -4.920069668238522e-19

R37_94 V37 V94 3733.3252800513687
L37_94 V37 V94 4.071528030726066e-12
C37_94 V37 V94 -2.3506856927996172e-20

R37_95 V37 V95 -16277.846794458457
L37_95 V37 V95 -4.260232138865793e-12
C37_95 V37 V95 -1.0097347131466284e-19

R37_96 V37 V96 -78376.76563387008
L37_96 V37 V96 -3.0920549141828387e-12
C37_96 V37 V96 -1.0406643017657972e-19

R37_97 V37 V97 4222.595772400737
L37_97 V37 V97 2.4183820404134077e-12
C37_97 V37 V97 1.7871751509076201e-19

R37_98 V37 V98 -1144.932534451439
L37_98 V37 V98 2.5786331386339617e-11
C37_98 V37 V98 1.9950373281609203e-19

R37_99 V37 V99 -1105.7784197737185
L37_99 V37 V99 -1.5514436471050318e-12
C37_99 V37 V99 -3.0772186398114563e-19

R37_100 V37 V100 -1377.242925517402
L37_100 V37 V100 -3.066246166659303e-12
C37_100 V37 V100 -1.5096046649069428e-19

R37_101 V37 V101 -2241.540247928993
L37_101 V37 V101 1.515544658768834e-11
C37_101 V37 V101 1.8616241661204104e-19

R37_102 V37 V102 113904.95062521104
L37_102 V37 V102 -2.6260621598126383e-12
C37_102 V37 V102 -1.3866499426057886e-19

R37_103 V37 V103 6336.489936993037
L37_103 V37 V103 8.768244165152356e-12
C37_103 V37 V103 9.567428533244237e-20

R37_104 V37 V104 19237.567676960734
L37_104 V37 V104 1.2521889899140423e-11
C37_104 V37 V104 1.2608311254000053e-19

R37_105 V37 V105 456.6089751838493
L37_105 V37 V105 1.906880743174517e-12
C37_105 V37 V105 1.2843421371020479e-19

R37_106 V37 V106 -32829.0570964769
L37_106 V37 V106 1.1104814086728691e-11
C37_106 V37 V106 -8.702424166513064e-20

R37_107 V37 V107 6423.469973960332
L37_107 V37 V107 3.016132721049935e-12
C37_107 V37 V107 2.273656115426135e-19

R37_108 V37 V108 9087.113497509286
L37_108 V37 V108 5.329442751221028e-12
C37_108 V37 V108 1.2172858973389165e-19

R37_109 V37 V109 -1878.5550965587408
L37_109 V37 V109 1.6605892162669244e-12
C37_109 V37 V109 1.1189253076263261e-19

R37_110 V37 V110 -21233.201019735305
L37_110 V37 V110 -1.2810122842249345e-10
C37_110 V37 V110 1.3129023666052028e-19

R37_111 V37 V111 -22872.82334776741
L37_111 V37 V111 3.1301041705799375e-12
C37_111 V37 V111 -1.9847968523365636e-21

R37_112 V37 V112 -9205.49695481287
L37_112 V37 V112 5.151253013107638e-12
C37_112 V37 V112 -6.193151929336398e-20

R37_113 V37 V113 -2770.80877687817
L37_113 V37 V113 -1.1636064879231513e-12
C37_113 V37 V113 -5.032518073243166e-19

R37_114 V37 V114 -8238.235562605138
L37_114 V37 V114 -2.7096352807339703e-11
C37_114 V37 V114 2.2535423652927734e-20

R37_115 V37 V115 -3280.469124415098
L37_115 V37 V115 -1.7869273042126315e-12
C37_115 V37 V115 -2.1240748771063081e-19

R37_116 V37 V116 -5170.402139726744
L37_116 V37 V116 -2.1507551224222997e-12
C37_116 V37 V116 -1.673301735773003e-19

R37_117 V37 V117 1133.9697555985763
L37_117 V37 V117 -2.9091176917018428e-12
C37_117 V37 V117 -3.5159680649526976e-20

R37_118 V37 V118 10970.29808600519
L37_118 V37 V118 -3.47131598999895e-11
C37_118 V37 V118 -8.796475911988165e-20

R37_119 V37 V119 -12260.958335590098
L37_119 V37 V119 5.055197940244618e-10
C37_119 V37 V119 7.925207101905786e-20

R37_120 V37 V120 -6128.979305355188
L37_120 V37 V120 -9.569670673171133e-12
C37_120 V37 V120 4.702317374140419e-20

R37_121 V37 V121 3578.135564868502
L37_121 V37 V121 9.20849348160385e-13
C37_121 V37 V121 4.0843264506049866e-19

R37_122 V37 V122 -5013.519904884484
L37_122 V37 V122 1.0236586425116863e-11
C37_122 V37 V122 3.228839363005538e-20

R37_123 V37 V123 5530.885225499257
L37_123 V37 V123 4.523057755452073e-12
C37_123 V37 V123 -7.766921393166153e-21

R37_124 V37 V124 3911.449331753735
L37_124 V37 V124 2.215816751509963e-12
C37_124 V37 V124 1.2106444518972034e-19

R37_125 V37 V125 1011.1473463678049
L37_125 V37 V125 4.667297106428272e-12
C37_125 V37 V125 1.016354645763398e-19

R37_126 V37 V126 21824.740673235043
L37_126 V37 V126 6.890192723573998e-12
C37_126 V37 V126 1.8749514245741632e-19

R37_127 V37 V127 -90859.36117759575
L37_127 V37 V127 -1.4405458109357795e-11
C37_127 V37 V127 9.495078724345054e-20

R37_128 V37 V128 13021.251483493215
L37_128 V37 V128 -3.345982929685312e-11
C37_128 V37 V128 6.03437106899751e-20

R37_129 V37 V129 -2782.396921123327
L37_129 V37 V129 4.229051739431276e-12
C37_129 V37 V129 1.480418799682297e-19

R37_130 V37 V130 -85992.01021748858
L37_130 V37 V130 -3.0798640103280184e-12
C37_130 V37 V130 -1.6998141900923702e-19

R37_131 V37 V131 -10535.547751456352
L37_131 V37 V131 5.1873251132179966e-11
C37_131 V37 V131 -9.216361656775872e-20

R37_132 V37 V132 -2291.2224685049614
L37_132 V37 V132 -4.3689999078484e-12
C37_132 V37 V132 -2.0398250337532146e-19

R37_133 V37 V133 -1254.8566094903474
L37_133 V37 V133 -1.1244765571378563e-12
C37_133 V37 V133 -6.95317947959504e-19

R37_134 V37 V134 -2544.319352468121
L37_134 V37 V134 1.6464576129060576e-11
C37_134 V37 V134 -1.9169946006449475e-20

R37_135 V37 V135 9362.797099186815
L37_135 V37 V135 -7.87891743146432e-11
C37_135 V37 V135 -5.504692792151627e-20

R37_136 V37 V136 4182.378727764571
L37_136 V37 V136 1.0344643692251066e-11
C37_136 V37 V136 -1.8215744522309045e-20

R37_137 V37 V137 862.761694628141
L37_137 V37 V137 -1.3381706795900314e-12
C37_137 V37 V137 -1.3575675585630793e-19

R37_138 V37 V138 1525.0455762574736
L37_138 V37 V138 4.567937228888176e-11
C37_138 V37 V138 8.357115307619998e-20

R37_139 V37 V139 -3335.902452484748
L37_139 V37 V139 -7.086327655567218e-12
C37_139 V37 V139 3.000444159308679e-20

R37_140 V37 V140 -7079.82737083225
L37_140 V37 V140 -2.943799327095925e-12
C37_140 V37 V140 -6.066140550411078e-20

R37_141 V37 V141 -3823.442728581914
L37_141 V37 V141 5.876922408805439e-13
C37_141 V37 V141 8.511667093376812e-19

R37_142 V37 V142 -1985.0831258989804
L37_142 V37 V142 3.816971877422763e-11
C37_142 V37 V142 5.292946597123019e-20

R37_143 V37 V143 -8655.106774703108
L37_143 V37 V143 1.2332596070567483e-10
C37_143 V37 V143 -3.006037217569986e-20

R37_144 V37 V144 -2097.439231737731
L37_144 V37 V144 5.064118877148411e-12
C37_144 V37 V144 1.5894123764065366e-19

R37_145 V37 V145 1209.460417269037
L37_145 V37 V145 1.5007869004953056e-12
C37_145 V37 V145 2.0070917646046537e-20

R37_146 V37 V146 -2039.864375763001
L37_146 V37 V146 4.791163420404836e-12
C37_146 V37 V146 -1.0121677336735635e-19

R37_147 V37 V147 6193.539194535688
L37_147 V37 V147 2.7809954672210855e-12
C37_147 V37 V147 2.2057398577807065e-19

R37_148 V37 V148 1197.6810233656965
L37_148 V37 V148 1.7520509685780047e-12
C37_148 V37 V148 1.4505280733733577e-19

R37_149 V37 V149 -479.97253875938793
L37_149 V37 V149 -7.325259735098094e-13
C37_149 V37 V149 -3.8206133857462807e-19

R37_150 V37 V150 1225.0249340775226
L37_150 V37 V150 9.72800554125904e-12
C37_150 V37 V150 1.8113328296492212e-19

R37_151 V37 V151 1917.6163053836167
L37_151 V37 V151 3.2557418096509685e-12
C37_151 V37 V151 -3.4133479679362686e-20

R37_152 V37 V152 -2661.9178187626303
L37_152 V37 V152 -5.7013752471064505e-12
C37_152 V37 V152 -9.91736488479643e-20

R37_153 V37 V153 662.9761898295495
L37_153 V37 V153 -1.5558538239406366e-12
C37_153 V37 V153 -2.574325027617971e-19

R37_154 V37 V154 -9099.969303227259
L37_154 V37 V154 -2.514766565140854e-12
C37_154 V37 V154 -1.5575817545847662e-19

R37_155 V37 V155 -913.7675346411772
L37_155 V37 V155 -1.869443149124481e-12
C37_155 V37 V155 -1.2178860966022133e-20

R37_156 V37 V156 10415.390738559234
L37_156 V37 V156 -3.254959564723094e-12
C37_156 V37 V156 -1.7690347838836556e-19

R37_157 V37 V157 812.6289954372228
L37_157 V37 V157 1.3997687970259564e-12
C37_157 V37 V157 -2.7823703421960514e-20

R37_158 V37 V158 -4430.512989866334
L37_158 V37 V158 -3.4458192675850356e-11
C37_158 V37 V158 -1.85393609523643e-20

R37_159 V37 V159 3333.429029845598
L37_159 V37 V159 -3.1182197535123675e-12
C37_159 V37 V159 -1.6073995843989309e-19

R37_160 V37 V160 -2456.8449323260998
L37_160 V37 V160 -3.2709522959394298e-12
C37_160 V37 V160 1.5306668566587974e-20

R37_161 V37 V161 1682.7624576470641
L37_161 V37 V161 5.2734348714622726e-12
C37_161 V37 V161 4.617212291552762e-19

R37_162 V37 V162 -2603.0383275404247
L37_162 V37 V162 -4.967298048131656e-12
C37_162 V37 V162 -1.7686994402866113e-19

R37_163 V37 V163 -2022.2688871008784
L37_163 V37 V163 -7.227893575226497e-12
C37_163 V37 V163 -6.115960089794248e-20

R37_164 V37 V164 10678.009412963578
L37_164 V37 V164 4.354045037417865e-12
C37_164 V37 V164 -1.1685909149480729e-21

R37_165 V37 V165 2070.8866878796034
L37_165 V37 V165 7.601012755300484e-13
C37_165 V37 V165 1.6408421702051193e-19

R37_166 V37 V166 -2534.5862668169916
L37_166 V37 V166 1.499840621992633e-12
C37_166 V37 V166 2.230292215382824e-19

R37_167 V37 V167 6566.9609520514905
L37_167 V37 V167 1.9590133245742957e-12
C37_167 V37 V167 1.5572509489984265e-19

R37_168 V37 V168 -1394.555515589257
L37_168 V37 V168 2.823002470989316e-12
C37_168 V37 V168 2.9611795456418127e-19

R37_169 V37 V169 9721.735445312113
L37_169 V37 V169 -2.0474516646251198e-12
C37_169 V37 V169 -3.5024680584677533e-19

R37_170 V37 V170 874.6248358927036
L37_170 V37 V170 -4.6641225318039515e-12
C37_170 V37 V170 -2.7957055915359266e-20

R37_171 V37 V171 1648.0445266953004
L37_171 V37 V171 8.952433971197217e-12
C37_171 V37 V171 6.384109282096079e-20

R37_172 V37 V172 1802.5488591137623
L37_172 V37 V172 4.8185268760958115e-11
C37_172 V37 V172 -8.611459727875758e-20

R37_173 V37 V173 1034.512973466938
L37_173 V37 V173 -7.555153121530671e-13
C37_173 V37 V173 -2.6630898203888656e-19

R37_174 V37 V174 -1153.274873027728
L37_174 V37 V174 -1.1569788160935253e-12
C37_174 V37 V174 -2.552397063216331e-19

R37_175 V37 V175 -1265.292072280502
L37_175 V37 V175 -1.340859439339862e-12
C37_175 V37 V175 -3.491645035506181e-19

R37_176 V37 V176 -1623.7992592094463
L37_176 V37 V176 -9.943564398693631e-13
C37_176 V37 V176 -4.448117031891003e-19

R37_177 V37 V177 -2392.5304687168623
L37_177 V37 V177 8.627530096472319e-13
C37_177 V37 V177 3.254889843205727e-19

R37_178 V37 V178 5823.64812565543
L37_178 V37 V178 3.223198641209669e-12
C37_178 V37 V178 6.16638747541994e-20

R37_179 V37 V179 -20848.09411317008
L37_179 V37 V179 5.187147456840469e-12
C37_179 V37 V179 1.3710571791289212e-19

R37_180 V37 V180 4036.637640930582
L37_180 V37 V180 2.0124972209605456e-12
C37_180 V37 V180 2.4352664848550883e-19

R37_181 V37 V181 -2268.364986603492
L37_181 V37 V181 -3.51188574271572e-12
C37_181 V37 V181 3.382025321596175e-19

R37_182 V37 V182 4536.839319089533
L37_182 V37 V182 1.4838224557643635e-11
C37_182 V37 V182 1.7396210631118372e-21

R37_183 V37 V183 2300.6497917815236
L37_183 V37 V183 3.2945155327935776e-12
C37_183 V37 V183 7.253020095113355e-20

R37_184 V37 V184 2967.097821068415
L37_184 V37 V184 1.6902298137722208e-12
C37_184 V37 V184 1.1491261815492887e-19

R37_185 V37 V185 575.390028765644
L37_185 V37 V185 -1.0800432352069688e-11
C37_185 V37 V185 -3.904895247917203e-19

R37_186 V37 V186 -1208.1237090545803
L37_186 V37 V186 1.033210124186839e-12
C37_186 V37 V186 3.1858903128928473e-19

R37_187 V37 V187 -3487.279879597095
L37_187 V37 V187 2.8988185071281388e-12
C37_187 V37 V187 -4.529947089984162e-21

R37_188 V37 V188 -2326.197714879091
L37_188 V37 V188 4.092743387754282e-11
C37_188 V37 V188 2.949848574837105e-20

R37_189 V37 V189 -541.9892112216271
L37_189 V37 V189 5.0904330254246214e-12
C37_189 V37 V189 -2.959293284464066e-20

R37_190 V37 V190 4081.676296710971
L37_190 V37 V190 -2.098513123455818e-12
C37_190 V37 V190 -6.488835766538429e-20

R37_191 V37 V191 1881.100880671163
L37_191 V37 V191 -2.5845106328169754e-12
C37_191 V37 V191 -8.727973509801691e-20

R37_192 V37 V192 2385.4373412676237
L37_192 V37 V192 -1.8041210115386259e-12
C37_192 V37 V192 -2.3656617804925795e-19

R37_193 V37 V193 -2011.6706895103887
L37_193 V37 V193 -1.651817017920105e-12
C37_193 V37 V193 -1.8221037742609087e-19

R37_194 V37 V194 1077.8226442211198
L37_194 V37 V194 -9.9424720795854e-13
C37_194 V37 V194 -2.3190954554777593e-19

R37_195 V37 V195 5200.56716190406
L37_195 V37 V195 5.2304020800559674e-12
C37_195 V37 V195 1.2350225425750697e-19

R37_196 V37 V196 2995.358250379126
L37_196 V37 V196 -5.02089939230445e-12
C37_196 V37 V196 -2.1309502424899206e-20

R37_197 V37 V197 632.4273529484191
L37_197 V37 V197 2.1238984759245967e-12
C37_197 V37 V197 3.997024717586604e-19

R37_198 V37 V198 -1410.7740478206692
L37_198 V37 V198 1.807364318404683e-12
C37_198 V37 V198 3.8370715184910953e-20

R37_199 V37 V199 -953.2453600189261
L37_199 V37 V199 3.2502423361748924e-12
C37_199 V37 V199 -1.1879837559109418e-19

R37_200 V37 V200 -983.3116276051023
L37_200 V37 V200 1.2889711172197847e-12
C37_200 V37 V200 2.3226808720138057e-19

R38_38 V38 0 -282.6861700747924
L38_38 V38 0 -2.6979822137963206e-13
C38_38 V38 0 -7.844387742709948e-19

R38_39 V38 V39 -12002.850647519454
L38_39 V38 V39 -4.5151862189875134e-12
C38_39 V38 V39 -7.07800401080731e-20

R38_40 V38 V40 -6698.666860069911
L38_40 V38 V40 -4.3279220296392986e-12
C38_40 V38 V40 -5.3957866051042524e-20

R38_41 V38 V41 11693.333174131947
L38_41 V38 V41 9.904740257267188e-12
C38_41 V38 V41 2.0957335570065335e-19

R38_42 V38 V42 -9246.513687192566
L38_42 V38 V42 2.4523209449591055e-12
C38_42 V38 V42 4.1781119737087874e-19

R38_43 V38 V43 -73247.59219813524
L38_43 V38 V43 -2.1778859293133217e-11
C38_43 V38 V43 8.443391450425845e-20

R38_44 V38 V44 -78089.25711649694
L38_44 V38 V44 -3.0686949392797426e-10
C38_44 V38 V44 1.156455075491613e-19

R38_45 V38 V45 4963.536036355373
L38_45 V38 V45 3.081545678506283e-12
C38_45 V38 V45 6.393112212203661e-20

R38_46 V38 V46 2617.912552584885
L38_46 V38 V46 1.0801665537313831e-12
C38_46 V38 V46 5.316109459758402e-19

R38_47 V38 V47 18176.100132878197
L38_47 V38 V47 5.236982990894951e-12
C38_47 V38 V47 5.221874303951565e-20

R38_48 V38 V48 5947.3336323523745
L38_48 V38 V48 2.9295893843503025e-12
C38_48 V38 V48 1.0411534411041563e-19

R38_49 V38 V49 11509.899892535856
L38_49 V38 V49 8.145347553240887e-11
C38_49 V38 V49 -5.260320904316642e-20

R38_50 V38 V50 7068.69394472582
L38_50 V38 V50 -1.7255046924176487e-12
C38_50 V38 V50 -3.1932299107979507e-19

R38_51 V38 V51 30473.27133770295
L38_51 V38 V51 3.934172215785668e-11
C38_51 V38 V51 -5.24183219068323e-20

R38_52 V38 V52 -10653947.755680356
L38_52 V38 V52 -3.873322320802986e-11
C38_52 V38 V52 -1.133296449192953e-19

R38_53 V38 V53 27503.63537099325
L38_53 V38 V53 2.2938023893152785e-12
C38_53 V38 V53 1.7396349452809932e-19

R38_54 V38 V54 -4960.304125995808
L38_54 V38 V54 -2.1856628867369956e-12
C38_54 V38 V54 -3.1641264652734023e-19

R38_55 V38 V55 -18235.66506374489
L38_55 V38 V55 -5.654305964494477e-11
C38_55 V38 V55 2.8566023750632663e-21

R38_56 V38 V56 -5210.021720234595
L38_56 V38 V56 -6.016638684753664e-12
C38_56 V38 V56 -7.59241366036615e-20

R38_57 V38 V57 -16324.114992136307
L38_57 V38 V57 -1.4164282010112128e-12
C38_57 V38 V57 -3.0741199791133616e-19

R38_58 V38 V58 22074.47655753731
L38_58 V38 V58 -4.185238939977105e-11
C38_58 V38 V58 -4.139359057958384e-22

R38_59 V38 V59 -30890.98601397203
L38_59 V38 V59 -1.3801585264072191e-11
C38_59 V38 V59 7.061710253622502e-20

R38_60 V38 V60 -11446.99803704891
L38_60 V38 V60 -9.51272324185501e-12
C38_60 V38 V60 7.771699472593436e-20

R38_61 V38 V61 15336.28734162315
L38_61 V38 V61 4.6923594310253464e-12
C38_61 V38 V61 1.1888156947997925e-19

R38_62 V38 V62 -8180.994823048167
L38_62 V38 V62 1.3048710017388615e-12
C38_62 V38 V62 4.434984188208082e-19

R38_63 V38 V63 2959355.9041793896
L38_63 V38 V63 -4.275228097603641e-12
C38_63 V38 V63 -1.4309517551234628e-19

R38_64 V38 V64 11024.960619169135
L38_64 V38 V64 -8.130780375196678e-12
C38_64 V38 V64 -1.238130906290368e-19

R38_65 V38 V65 6599.580772104041
L38_65 V38 V65 2.548073986751701e-12
C38_65 V38 V65 2.458430872987239e-19

R38_66 V38 V66 7163.651412058819
L38_66 V38 V66 -2.2274525168651856e-12
C38_66 V38 V66 -1.158847187035096e-19

R38_67 V38 V67 -31333.257075930807
L38_67 V38 V67 9.300275515928662e-12
C38_67 V38 V67 2.6434374203168052e-20

R38_68 V38 V68 18194.534031793257
L38_68 V38 V68 2.959231395028482e-12
C38_68 V38 V68 1.0575759490851186e-19

R38_69 V38 V69 -16856.97634089751
L38_69 V38 V69 -1.8921707279629325e-11
C38_69 V38 V69 -1.6327650167351108e-19

R38_70 V38 V70 3365.6986451288803
L38_70 V38 V70 -3.3705845848227813e-12
C38_70 V38 V70 -3.1569557136319637e-19

R38_71 V38 V71 16345.45002343044
L38_71 V38 V71 3.2536838024126852e-12
C38_71 V38 V71 1.4796361383120657e-19

R38_72 V38 V72 24572.084477780783
L38_72 V38 V72 4.0792872928119315e-12
C38_72 V38 V72 1.1497648006215873e-19

R38_73 V38 V73 6707.519210250184
L38_73 V38 V73 6.942058873686537e-11
C38_73 V38 V73 -2.3659291648343586e-20

R38_74 V38 V74 -5482.252876072069
L38_74 V38 V74 1.3556304208835254e-12
C38_74 V38 V74 2.8214988137738073e-19

R38_75 V38 V75 22148.017214083473
L38_75 V38 V75 -3.284503424889852e-12
C38_75 V38 V75 -1.2037101870934194e-19

R38_76 V38 V76 -6459.463198901903
L38_76 V38 V76 -1.6017467194427135e-12
C38_76 V38 V76 -2.8389393071188726e-19

R38_77 V38 V77 -18842.440084184986
L38_77 V38 V77 -4.833728155360179e-12
C38_77 V38 V77 -4.04724916454798e-20

R38_78 V38 V78 -4135.5754525309485
L38_78 V38 V78 -3.203092613196195e-12
C38_78 V38 V78 -8.759092195785189e-20

R38_79 V38 V79 -7989.9246464229755
L38_79 V38 V79 -5.3921378365176324e-11
C38_79 V38 V79 -1.7460769357566362e-20

R38_80 V38 V80 -31752.01569631509
L38_80 V38 V80 4.754097067418943e-12
C38_80 V38 V80 8.480896129373791e-20

R38_81 V38 V81 4797.856814309712
L38_81 V38 V81 4.106243528538614e-12
C38_81 V38 V81 1.1098191176129322e-19

R38_82 V38 V82 5466.641639602103
L38_82 V38 V82 -1.1692130225978467e-11
C38_82 V38 V82 -8.787846183627523e-20

R38_83 V38 V83 -70356.43975434851
L38_83 V38 V83 1.0689554470524167e-11
C38_83 V38 V83 5.94991050209904e-20

R38_84 V38 V84 16396.072800318514
L38_84 V38 V84 3.0792840771273842e-12
C38_84 V38 V84 1.7266925951787293e-19

R38_85 V38 V85 190086.82144916768
L38_85 V38 V85 3.3131096451556563e-12
C38_85 V38 V85 1.329783539821904e-19

R38_86 V38 V86 1501.0494224756505
L38_86 V38 V86 2.2298479736555377e-12
C38_86 V38 V86 2.8845106301539094e-19

R38_87 V38 V87 -19123.60511157152
L38_87 V38 V87 -3.628968563577662e-12
C38_87 V38 V87 -1.6545097920795448e-19

R38_88 V38 V88 -12574.68381890248
L38_88 V38 V88 -2.5243406237416104e-12
C38_88 V38 V88 -2.435894499812792e-19

R38_89 V38 V89 -25333.413613662648
L38_89 V38 V89 -1.4355638309549356e-11
C38_89 V38 V89 -1.1657275068473715e-19

R38_90 V38 V90 -1221.4850567510498
L38_90 V38 V90 -1.459252357488873e-12
C38_90 V38 V90 -3.5013291744125346e-19

R38_91 V38 V91 7137.1214650043485
L38_91 V38 V91 1.7827741978263536e-12
C38_91 V38 V91 2.8909358629020957e-19

R38_92 V38 V92 6271.3442516183095
L38_92 V38 V92 1.7555059730195924e-12
C38_92 V38 V92 2.422346725470156e-19

R38_93 V38 V93 10165.728237174499
L38_93 V38 V93 -2.888956401046781e-12
C38_93 V38 V93 -1.4800149901675584e-19

R38_94 V38 V94 -6811.832968321161
L38_94 V38 V94 1.0393131896784806e-11
C38_94 V38 V94 -2.0161078482684856e-20

R38_95 V38 V95 59283.05824045647
L38_95 V38 V95 -1.3246303204417952e-11
C38_95 V38 V95 5.2446766495029245e-20

R38_96 V38 V96 -10374.778653968158
L38_96 V38 V96 -5.149625738825195e-12
C38_96 V38 V96 6.083749622058763e-20

R38_97 V38 V97 -19792.323146855855
L38_97 V38 V97 4.856739111873645e-12
C38_97 V38 V97 1.565394588692667e-19

R38_98 V38 V98 1523.473472830947
L38_98 V38 V98 1.6723066261952928e-12
C38_98 V38 V98 2.798898589388711e-19

R38_99 V38 V99 -1945.1979963248166
L38_99 V38 V99 -1.4109831791524062e-12
C38_99 V38 V99 -4.0987488584084e-19

R38_100 V38 V100 -2296.9727868077453
L38_100 V38 V100 -2.0673193975818843e-12
C38_100 V38 V100 -3.479548355589725e-19

R38_101 V38 V101 277157.00597842626
L38_101 V38 V101 6.451440659555703e-11
C38_101 V38 V101 1.5241703003093697e-20

R38_102 V38 V102 -1875.1446162189675
L38_102 V38 V102 -1.8491933334998653e-12
C38_102 V38 V102 -1.2356273061845323e-19

R38_103 V38 V103 2545.4978357530804
L38_103 V38 V103 3.344260110998276e-12
C38_103 V38 V103 1.5161216221031658e-19

R38_104 V38 V104 2087.1578200644776
L38_104 V38 V104 2.8826848816683977e-12
C38_104 V38 V104 1.893217724645506e-19

R38_105 V38 V105 2281.4748038732455
L38_105 V38 V105 7.032325682129135e-12
C38_105 V38 V105 -2.000547668940624e-20

R38_106 V38 V106 1214.2280434594293
L38_106 V38 V106 9.615049533760541e-11
C38_106 V38 V106 -1.1498425977157988e-19

R38_107 V38 V107 17888.289988404547
L38_107 V38 V107 4.897924614440113e-12
C38_107 V38 V107 1.914593192605424e-19

R38_108 V38 V108 -240671.30686399795
L38_108 V38 V108 -2.183297257394453e-11
C38_108 V38 V108 5.2629532525474073e-20

R38_109 V38 V109 -3345.7296821010045
L38_109 V38 V109 1.2888577093903919e-11
C38_109 V38 V109 1.288842937798518e-19

R38_110 V38 V110 -1402.8654874182375
L38_110 V38 V110 -6.61739797128943e-12
C38_110 V38 V110 -8.430178509135434e-20

R38_111 V38 V111 -5271.378557115959
L38_111 V38 V111 6.0153292140163775e-12
C38_111 V38 V111 -4.179551376976156e-20

R38_112 V38 V112 -4119.6947503012225
L38_112 V38 V112 3.7037122023728765e-12
C38_112 V38 V112 3.8884869990141783e-20

R38_113 V38 V113 -9570.261904146711
L38_113 V38 V113 -3.704292866378031e-12
C38_113 V38 V113 -1.3934155552629006e-19

R38_114 V38 V114 -1520.2007510781216
L38_114 V38 V114 7.029255864163653e-12
C38_114 V38 V114 3.381705365811984e-19

R38_115 V38 V115 -7545.935022783536
L38_115 V38 V115 -2.154770538347511e-12
C38_115 V38 V115 -1.4289973217617776e-19

R38_116 V38 V116 -7892.714138086343
L38_116 V38 V116 -2.1950081010796646e-12
C38_116 V38 V116 -1.1209090632142092e-19

R38_117 V38 V117 9455.322044807326
L38_117 V38 V117 -9.35952559170483e-12
C38_117 V38 V117 -1.1231562566533544e-19

R38_118 V38 V118 585.5647852450917
L38_118 V38 V118 3.1136918088113246e-12
C38_118 V38 V118 -1.568683359132169e-19

R38_119 V38 V119 3195.850097801655
L38_119 V38 V119 -1.2057502003092451e-11
C38_119 V38 V119 -3.577163865427135e-20

R38_120 V38 V120 3030.8756907476754
L38_120 V38 V120 -3.779714722563272e-12
C38_120 V38 V120 -1.4640550355734202e-19

R38_121 V38 V121 4521.950520911427
L38_121 V38 V121 3.685855694950294e-12
C38_121 V38 V121 2.428555314437666e-19

R38_122 V38 V122 -2570.292522167836
L38_122 V38 V122 -2.258444043766137e-12
C38_122 V38 V122 -1.8527312260321058e-19

R38_123 V38 V123 9891.313562539623
L38_123 V38 V123 1.7644022629654373e-12
C38_123 V38 V123 1.7954947229811542e-19

R38_124 V38 V124 10770.624373540419
L38_124 V38 V124 1.1566115689308035e-12
C38_124 V38 V124 3.744555938029557e-19

R38_125 V38 V125 2437.586787844432
L38_125 V38 V125 1.6246261659904248e-11
C38_125 V38 V125 6.040778998188383e-21

R38_126 V38 V126 -830.6305104806189
L38_126 V38 V126 5.349942208006734e-12
C38_126 V38 V126 4.04290580541765e-19

R38_127 V38 V127 -1628.642432989339
L38_127 V38 V127 -3.9357393674569044e-12
C38_127 V38 V127 2.195763249214309e-20

R38_128 V38 V128 -1523.8536201408158
L38_128 V38 V128 -3.06626851543411e-12
C38_128 V38 V128 -2.1229238038229565e-20

R38_129 V38 V129 -1583.6029228403659
L38_129 V38 V129 1.3677056555683326e-11
C38_129 V38 V129 2.1660235615702326e-20

R38_130 V38 V130 1537.8551542443588
L38_130 V38 V130 8.854261219214884e-12
C38_130 V38 V130 -1.8706102742498967e-19

R38_131 V38 V131 1548.8327448563018
L38_131 V38 V131 -1.3097891866625469e-11
C38_131 V38 V131 -1.6831999171068956e-19

R38_132 V38 V132 1208.4500244970193
L38_132 V38 V132 -3.3604549587895165e-12
C38_132 V38 V132 -3.165653537673391e-19

R38_133 V38 V133 -5931.761347532372
L38_133 V38 V133 -5.123738096126127e-12
C38_133 V38 V133 -1.4884478097561609e-19

R38_134 V38 V134 1296.3978987628586
L38_134 V38 V134 -2.372978612232846e-12
C38_134 V38 V134 -1.5954498377868978e-19

R38_135 V38 V135 3202.41923369289
L38_135 V38 V135 2.684131746108832e-12
C38_135 V38 V135 1.5588892089188007e-19

R38_136 V38 V136 1743.2012875697428
L38_136 V38 V136 1.9130041457444094e-12
C38_136 V38 V136 2.554872140225561e-19

R38_137 V38 V137 1129.023903559385
L38_137 V38 V137 -2.6684967751777763e-12
C38_137 V38 V137 -9.090629286538877e-20

R38_138 V38 V138 -1303.1901574786993
L38_138 V38 V138 2.7714493070563368e-12
C38_138 V38 V138 2.972802652432798e-19

R38_139 V38 V139 -1124.6917420956115
L38_139 V38 V139 -1.567418838156401e-12
C38_139 V38 V139 -1.4878180051548906e-19

R38_140 V38 V140 -891.5165967996246
L38_140 V38 V140 -1.36561106860782e-12
C38_140 V38 V140 -2.0909781428555088e-19

R38_141 V38 V141 8176.020473237175
L38_141 V38 V141 1.6496780606664766e-12
C38_141 V38 V141 3.212041494608621e-19

R38_142 V38 V142 -801.6269367847732
L38_142 V38 V142 9.667359214654302e-12
C38_142 V38 V142 -8.314024945214284e-20

R38_143 V38 V143 2602.431594317798
L38_143 V38 V143 4.538255510142092e-12
C38_143 V38 V143 -1.6252172588214358e-21

R38_144 V38 V144 -19635.09145020673
L38_144 V38 V144 4.344070732743648e-12
C38_144 V38 V144 5.51063205461935e-20

R38_145 V38 V145 -1614.6007535662545
L38_145 V38 V145 1.6221903848457026e-12
C38_145 V38 V145 1.0435956806399013e-19

R38_146 V38 V146 523.6260350429352
L38_146 V38 V146 3.1104996291083415e-12
C38_146 V38 V146 -7.165450164805168e-20

R38_147 V38 V147 -19215.055103205967
L38_147 V38 V147 1.6709050489742304e-12
C38_147 V38 V147 3.144078166749954e-19

R38_148 V38 V148 1043.3361139633528
L38_148 V38 V148 1.3427193436863293e-12
C38_148 V38 V148 2.3355393693711467e-19

R38_149 V38 V149 -2995.968701253585
L38_149 V38 V149 -1.27064184719181e-12
C38_149 V38 V149 -3.2084971838200217e-19

R38_150 V38 V150 1021.6210343338939
L38_150 V38 V150 -7.434105289980647e-12
C38_150 V38 V150 1.6933150196092064e-19

R38_151 V38 V151 -7942.836280614688
L38_151 V38 V151 -9.04507692389203e-12
C38_151 V38 V151 -1.3611869661452865e-19

R38_152 V38 V152 -745.3984637715449
L38_152 V38 V152 -2.8181071430334445e-12
C38_152 V38 V152 -9.274724630523721e-20

R38_153 V38 V153 1210.6296753895226
L38_153 V38 V153 -1.6111528466462343e-12
C38_153 V38 V153 -1.52194802127241e-19

R38_154 V38 V154 -860.2498956586904
L38_154 V38 V154 -1.6572383080835474e-12
C38_154 V38 V154 -7.15894945193481e-20

R38_155 V38 V155 -1700.5420865232074
L38_155 V38 V155 -1.4536895942238121e-12
C38_155 V38 V155 -6.341221555910342e-20

R38_156 V38 V156 668.602490084156
L38_156 V38 V156 -3.0564743240195235e-12
C38_156 V38 V156 -2.121485493620666e-19

R38_157 V38 V157 3344.4590705096293
L38_157 V38 V157 2.9453646422644244e-12
C38_157 V38 V157 2.235511759556744e-19

R38_158 V38 V158 -5276.495213594178
L38_158 V38 V158 2.2070350876788873e-12
C38_158 V38 V158 -1.2067173053572167e-19

R38_159 V38 V159 755.4584941380449
L38_159 V38 V159 4.892466247644552e-12
C38_159 V38 V159 -1.2824836741741226e-20

R38_160 V38 V160 3231.5875420760954
L38_160 V38 V160 8.969000410907319e-12
C38_160 V38 V160 1.1659515537980195e-19

R38_161 V38 V161 -1368.609516352121
L38_161 V38 V161 4.557052639369139e-12
C38_161 V38 V161 8.844240021376632e-20

R38_162 V38 V162 2603.735730882778
L38_162 V38 V162 2.916880711469052e-12
C38_162 V38 V162 -6.675918007865733e-20

R38_163 V38 V163 -1027.28371887797
L38_163 V38 V163 9.613966751216287e-11
C38_163 V38 V163 -5.611991185099693e-20

R38_164 V38 V164 -1108.713916839644
L38_164 V38 V164 3.992100737172592e-12
C38_164 V38 V164 -7.924304513924824e-20

R38_165 V38 V165 1735.2589238171472
L38_165 V38 V165 1.3810940451471236e-12
C38_165 V38 V165 5.926903188585938e-20

R38_166 V38 V166 1570.3577745216376
L38_166 V38 V166 -2.291843113973126e-12
C38_166 V38 V166 1.5725102124552403e-19

R38_167 V38 V167 5158.920877748194
L38_167 V38 V167 3.740741402475112e-12
C38_167 V38 V167 -2.8405056318025276e-22

R38_168 V38 V168 -2992.4053716642825
L38_168 V38 V168 7.377324845979699e-12
C38_168 V38 V168 9.356327477330925e-20

R38_169 V38 V169 1128.696416056979
L38_169 V38 V169 -3.974984575823298e-12
C38_169 V38 V169 -2.4890536047263446e-20

R38_170 V38 V170 -2162.3409689968007
L38_170 V38 V170 -1.6723940308378775e-11
C38_170 V38 V170 -2.5247566979607684e-20

R38_171 V38 V171 2037.1074924737618
L38_171 V38 V171 1.017571718383709e-11
C38_171 V38 V171 1.0436952251349173e-19

R38_172 V38 V172 1253.7863542187038
L38_172 V38 V172 4.306847541448255e-12
C38_172 V38 V172 4.772326917062123e-20

R38_173 V38 V173 -1786.3017203536997
L38_173 V38 V173 -1.587498526091503e-12
C38_173 V38 V173 -2.1013463347349254e-19

R38_174 V38 V174 -1912.4792211438462
L38_174 V38 V174 1.8672685307414226e-12
C38_174 V38 V174 -7.31421973492745e-20

R38_175 V38 V175 -4194.534558302761
L38_175 V38 V175 -2.312539920586232e-12
C38_175 V38 V175 -2.29249156962581e-19

R38_176 V38 V176 -2431.448648560653
L38_176 V38 V176 -1.3845106274958891e-12
C38_176 V38 V176 -3.005226939985521e-19

R38_177 V38 V177 -16326.41349320754
L38_177 V38 V177 2.1934390140139274e-12
C38_177 V38 V177 1.4883853796005399e-19

R38_178 V38 V178 1698.903320444527
L38_178 V38 V178 -5.842850811067115e-12
C38_178 V38 V178 2.1359605442689806e-20

R38_179 V38 V179 -4235.058595866658
L38_179 V38 V179 5.925173148189994e-12
C38_179 V38 V179 1.6201791296559247e-19

R38_180 V38 V180 21171.311625421364
L38_180 V38 V180 3.1693007707313355e-12
C38_180 V38 V180 2.122005548184752e-19

R38_181 V38 V181 3331.579266363048
L38_181 V38 V181 6.945642347663814e-12
C38_181 V38 V181 1.7433254614722074e-19

R38_182 V38 V182 8276.813830046827
L38_182 V38 V182 -2.362774185021985e-12
C38_182 V38 V182 -4.508045047063243e-20

R38_183 V38 V183 2168.614755979819
L38_183 V38 V183 3.262077510544126e-12
C38_183 V38 V183 2.5772183792068204e-20

R38_184 V38 V184 2784.3601223525316
L38_184 V38 V184 1.9320315237592697e-12
C38_184 V38 V184 5.262807753016919e-20

R38_185 V38 V185 5316.656816556893
L38_185 V38 V185 -8.175890033354905e-12
C38_185 V38 V185 -1.9719379280237612e-19

R38_186 V38 V186 -7983.053887296554
L38_186 V38 V186 1.1758442402159316e-12
C38_186 V38 V186 1.6531507003467052e-19

R38_187 V38 V187 -4632.476353917506
L38_187 V38 V187 6.382114470980798e-12
C38_187 V38 V187 -8.568310143783029e-20

R38_188 V38 V188 -1130.7805862539508
L38_188 V38 V188 -3.0743507781980408e-12
C38_188 V38 V188 -7.987947960269108e-20

R38_189 V38 V189 -4621.049297051856
L38_189 V38 V189 -5.459020716979719e-12
C38_189 V38 V189 5.622903228822903e-22

R38_190 V38 V190 3436.6305072193113
L38_190 V38 V190 -6.5153879576289606e-12
C38_190 V38 V190 -1.787014132203354e-20

R38_191 V38 V191 -6186.90734262195
L38_191 V38 V191 -3.793429703497677e-12
C38_191 V38 V191 2.3078374029834262e-20

R38_192 V38 V192 6072.196229218008
L38_192 V38 V192 -1.4700573812101426e-11
C38_192 V38 V192 3.563444464934524e-20

R38_193 V38 V193 -2755.181452108537
L38_193 V38 V193 -8.340175912514733e-11
C38_193 V38 V193 -1.1340070170714467e-20

R38_194 V38 V194 10980.145672259114
L38_194 V38 V194 -4.967313162994934e-12
C38_194 V38 V194 2.2771174069850023e-20

R38_195 V38 V195 2388.8873283837825
L38_195 V38 V195 1.0255035883238691e-11
C38_195 V38 V195 4.964239293524221e-21

R38_196 V38 V196 1869.0891655079981
L38_196 V38 V196 -3.263099670380869e-12
C38_196 V38 V196 -2.2553421039182696e-19

R38_197 V38 V197 10932.726834437235
L38_197 V38 V197 9.989915074961733e-12
C38_197 V38 V197 8.402457668299246e-20

R38_198 V38 V198 -7923.785164813073
L38_198 V38 V198 6.537830252470392e-12
C38_198 V38 V198 2.1131635161565194e-20

R38_199 V38 V199 -19637.304172716096
L38_199 V38 V199 1.3417617555798178e-11
C38_199 V38 V199 -1.0765703327212658e-19

R38_200 V38 V200 -1735.8967664472445
L38_200 V38 V200 2.386384725808421e-12
C38_200 V38 V200 1.0933426288820886e-19

R39_39 V39 0 -233.6038478457959
L39_39 V39 0 -4.999687247414921e-13
C39_39 V39 0 2.4244727766901285e-19

R39_40 V39 V40 -1127.7678757964065
L39_40 V39 V40 -2.7018634754483286e-12
C39_40 V39 V40 -2.984446471312338e-19

R39_41 V39 V41 5261.510603101501
L39_41 V39 V41 -1.2316896676724567e-11
C39_41 V39 V41 1.4707226109300186e-20

R39_42 V39 V42 9989.449821231126
L39_42 V39 V42 -2.3531770954273404e-11
C39_42 V39 V42 -9.388262732414771e-21

R39_43 V39 V43 -96421.1896371073
L39_43 V39 V43 9.604089210399276e-12
C39_43 V39 V43 2.195577447603899e-19

R39_44 V39 V44 4457.036811045654
L39_44 V39 V44 -1.77557400623599e-11
C39_44 V39 V44 1.0717180052361799e-19

R39_45 V39 V45 4971.272642369002
L39_45 V39 V45 6.029774833588582e-12
C39_45 V39 V45 -1.0766932515095119e-20

R39_46 V39 V46 5850.501415276515
L39_46 V39 V46 -1.8538138302989514e-11
C39_46 V39 V46 -1.160888704354634e-19

R39_47 V39 V47 903.8991204790356
L39_47 V39 V47 1.2841530356367921e-12
C39_47 V39 V47 5.345054647178273e-19

R39_48 V39 V48 1956.4034646452474
L39_48 V39 V48 -2.210642723263587e-11
C39_48 V39 V48 -1.1181291959635132e-19

R39_49 V39 V49 257502.11361047637
L39_49 V39 V49 1.3828810450125886e-11
C39_49 V39 V49 -4.817055181346135e-20

R39_50 V39 V50 24136.928733501798
L39_50 V39 V50 8.162346396021398e-12
C39_50 V39 V50 9.27441709159795e-20

R39_51 V39 V51 2979.87656682788
L39_51 V39 V51 -1.22185572901663e-12
C39_51 V39 V51 -5.62150982236825e-19

R39_52 V39 V52 -35171.43410969072
L39_52 V39 V52 7.566195161919422e-12
C39_52 V39 V52 6.44829455071135e-20

R39_53 V39 V53 5486.794020353776
L39_53 V39 V53 2.054982778876913e-12
C39_53 V39 V53 2.404010814852674e-19

R39_54 V39 V54 40172.848401225514
L39_54 V39 V54 6.0211269072918354e-12
C39_54 V39 V54 1.2412686774928016e-19

R39_55 V39 V55 -3041.2433981521644
L39_55 V39 V55 4.162908577341383e-12
C39_55 V39 V55 1.4050745626237177e-19

R39_56 V39 V56 -3223.876939007108
L39_56 V39 V56 4.337047283462895e-12
C39_56 V39 V56 1.907046246031888e-19

R39_57 V39 V57 -5985.53121478
L39_57 V39 V57 -1.9751741770925625e-12
C39_57 V39 V57 -2.5670601585449307e-19

R39_58 V39 V58 3482.2749599399576
L39_58 V39 V58 -7.207613784452268e-12
C39_58 V39 V58 -9.662019074038004e-20

R39_59 V39 V59 -1708.2753531881062
L39_59 V39 V59 5.507720702909124e-12
C39_59 V39 V59 1.047801693798845e-19

R39_60 V39 V60 -2664.703440631177
L39_60 V39 V60 -3.2149344475532253e-12
C39_60 V39 V60 -1.8452182903996935e-19

R39_61 V39 V61 10921.137703976658
L39_61 V39 V61 7.053274625998516e-11
C39_61 V39 V61 -1.3100697297578755e-20

R39_62 V39 V62 -3116.1273088864664
L39_62 V39 V62 -1.0246538711181364e-11
C39_62 V39 V62 -1.0838177431106911e-19

R39_63 V39 V63 110867.98283855047
L39_63 V39 V63 -1.670972694956696e-11
C39_63 V39 V63 -1.0274847080476018e-19

R39_64 V39 V64 5284.203376596181
L39_64 V39 V64 -6.387409704153566e-12
C39_64 V39 V64 -8.056551769603503e-20

R39_65 V39 V65 6627.606926702627
L39_65 V39 V65 5.074360489233076e-12
C39_65 V39 V65 8.449601376688261e-20

R39_66 V39 V66 12082.164560008456
L39_66 V39 V66 7.561691563873547e-12
C39_66 V39 V66 7.659275783766264e-20

R39_67 V39 V67 2202.642247966503
L39_67 V39 V67 -3.096550001943206e-12
C39_67 V39 V67 -5.264146799888164e-20

R39_68 V39 V68 2997.646706036203
L39_68 V39 V68 3.249077299315408e-12
C39_68 V39 V68 1.7534067805273552e-19

R39_69 V39 V69 -209469.10963948877
L39_69 V39 V69 5.193683660489814e-12
C39_69 V39 V69 6.157185384907799e-20

R39_70 V39 V70 5952.307942748368
L39_70 V39 V70 2.0850468181838842e-10
C39_70 V39 V70 8.718825572913113e-21

R39_71 V39 V71 1645.6791005716475
L39_71 V39 V71 6.369226771684718e-12
C39_71 V39 V71 4.0960928972112584e-20

R39_72 V39 V72 4015.407868156441
L39_72 V39 V72 3.7346562835789364e-11
C39_72 V39 V72 -4.422767187689263e-20

R39_73 V39 V73 3610.193119395339
L39_73 V39 V73 6.294299563585045e-11
C39_73 V39 V73 -4.179540308286064e-20

R39_74 V39 V74 -6267.691376741987
L39_74 V39 V74 -1.0195585313061058e-11
C39_74 V39 V74 -8.883551534737415e-20

R39_75 V39 V75 -1796.0167040203594
L39_75 V39 V75 2.343986426524083e-12
C39_75 V39 V75 1.8160823748054991e-19

R39_76 V39 V76 -1832.4885835681198
L39_76 V39 V76 -4.179125487727611e-12
C39_76 V39 V76 -3.6177184210651514e-20

R39_77 V39 V77 -3966.158467611366
L39_77 V39 V77 -3.9635001771725514e-12
C39_77 V39 V77 -1.336167458449989e-19

R39_78 V39 V78 5443.986207483674
L39_78 V39 V78 4.853092197370748e-12
C39_78 V39 V78 1.8692355768280831e-19

R39_79 V39 V79 -1056.3379573604886
L39_79 V39 V79 -3.2370251763076777e-12
C39_79 V39 V79 -2.206774632518201e-19

R39_80 V39 V80 -3450.213564597023
L39_80 V39 V80 4.831965286165502e-12
C39_80 V39 V80 5.4021863893050707e-20

R39_81 V39 V81 7458.257940364423
L39_81 V39 V81 6.755364730591395e-12
C39_81 V39 V81 5.0491759095819044e-20

R39_82 V39 V82 -7340.854416404642
L39_82 V39 V82 -7.475371557467717e-12
C39_82 V39 V82 -1.519200056738014e-19

R39_83 V39 V83 2421.6967711481725
L39_83 V39 V83 -2.4767656334764562e-12
C39_83 V39 V83 -1.7122883859514448e-19

R39_84 V39 V84 3884.5591785359297
L39_84 V39 V84 -6.527192639122178e-12
C39_84 V39 V84 -7.744710666677896e-20

R39_85 V39 V85 -517653.1766721813
L39_85 V39 V85 4.3405559392652966e-11
C39_85 V39 V85 -1.6134074889279747e-20

R39_86 V39 V86 2781.635629570433
L39_86 V39 V86 -3.87308512687032e-12
C39_86 V39 V86 -1.6630409334179904e-19

R39_87 V39 V87 653.147831927541
L39_87 V39 V87 1.5739663269743451e-12
C39_87 V39 V87 5.680163538659724e-19

R39_88 V39 V88 3516.01683232456
L39_88 V39 V88 -1.1760380964427466e-11
C39_88 V39 V88 5.725827243341856e-20

R39_89 V39 V89 3714.4061553563756
L39_89 V39 V89 3.2285324244027497e-12
C39_89 V39 V89 1.7214294203191477e-19

R39_90 V39 V90 13753.257177906062
L39_90 V39 V90 3.017359391243625e-12
C39_90 V39 V90 3.5160259286794744e-19

R39_91 V39 V91 -761.4981409852415
L39_91 V39 V91 -1.6360241827056978e-12
C39_91 V39 V91 -5.696676490013029e-19

R39_92 V39 V92 -11963.599919663431
L39_92 V39 V92 3.955523058492044e-12
C39_92 V39 V92 2.4566724071522803e-20

R39_93 V39 V93 6548.453398782022
L39_93 V39 V93 -6.210610574173448e-12
C39_93 V39 V93 -4.4001884513394106e-20

R39_94 V39 V94 -3470.165691725349
L39_94 V39 V94 5.404280388546952e-12
C39_94 V39 V94 5.216596778147468e-21

R39_95 V39 V95 -571.2115138905457
L39_95 V39 V95 -1.1805960324495616e-11
C39_95 V39 V95 -3.058184451364917e-19

R39_96 V39 V96 -1251.3798169002466
L39_96 V39 V96 -9.477731966404509e-12
C39_96 V39 V96 -7.091754310622032e-20

R39_97 V39 V97 -1369.1814445702853
L39_97 V39 V97 -3.1017441072858517e-12
C39_97 V39 V97 -3.9591074552412287e-19

R39_98 V39 V98 6276.340090740443
L39_98 V39 V98 -2.2085214279299953e-12
C39_98 V39 V98 -3.278000727336297e-19

R39_99 V39 V99 356.19835524317614
L39_99 V39 V99 1.4935602668734135e-12
C39_99 V39 V99 7.209066836902455e-19

R39_100 V39 V100 2424.9557337722094
L39_100 V39 V100 -7.513629886531485e-12
C39_100 V39 V100 5.34097080795663e-20

R39_101 V39 V101 3734.3198061872968
L39_101 V39 V101 2.6281039572997537e-12
C39_101 V39 V101 2.7123860743700223e-19

R39_102 V39 V102 -10517.27826540461
L39_102 V39 V102 -7.783607356057144e-12
C39_102 V39 V102 2.788476637945113e-20

R39_103 V39 V103 -1283.1843601545788
L39_103 V39 V103 -2.090998752120493e-12
C39_103 V39 V103 -1.35906375841734e-19

R39_104 V39 V104 3422.627975484533
L39_104 V39 V104 -7.219714660638809e-12
C39_104 V39 V104 -7.573922569948004e-20

R39_105 V39 V105 1075.8577924629874
L39_105 V39 V105 6.92990522769187e-12
C39_105 V39 V105 1.718483283740945e-19

R39_106 V39 V106 975.8541645225346
L39_106 V39 V106 1.7038968535631346e-12
C39_106 V39 V106 4.495865580866593e-19

R39_107 V39 V107 -946.3959946490924
L39_107 V39 V107 5.11355034241267e-11
C39_107 V39 V107 -3.217859427979199e-19

R39_108 V39 V108 -6676.842728544225
L39_108 V39 V108 5.298632580940959e-12
C39_108 V39 V108 1.143708445343326e-19

R39_109 V39 V109 -2463.5511985171
L39_109 V39 V109 -4.7883081117701585e-12
C39_109 V39 V109 -2.5063582767068006e-19

R39_110 V39 V110 -1320.090757240512
L39_110 V39 V110 -4.235957636063673e-12
C39_110 V39 V110 -2.354965750672008e-19

R39_111 V39 V111 377.97307283801763
L39_111 V39 V111 -2.841254400795063e-12
C39_111 V39 V111 -1.4624400322802064e-19

R39_112 V39 V112 1485.3082342406863
L39_112 V39 V112 3.641919736175122e-12
C39_112 V39 V112 9.139383790053882e-20

R39_113 V39 V113 -1565.2462188631725
L39_113 V39 V113 3.018264133038738e-11
C39_113 V39 V113 -1.3718544222610917e-19

R39_114 V39 V114 -968.7464749125758
L39_114 V39 V114 -2.1935117793370055e-12
C39_114 V39 V114 -3.537780990048273e-19

R39_115 V39 V115 -619.0353253809003
L39_115 V39 V115 1.6801115703082557e-12
C39_115 V39 V115 4.799552297459302e-19

R39_116 V39 V116 -995.3615237755605
L39_116 V39 V116 -2.3919434799191857e-12
C39_116 V39 V116 -2.205592240531053e-19

R39_117 V39 V117 -8701.550258234713
L39_117 V39 V117 1.9178907397189028e-11
C39_117 V39 V117 1.0534229576730346e-19

R39_118 V39 V118 645.4759281371563
L39_118 V39 V118 3.771454999699485e-12
C39_118 V39 V118 3.1881757129329643e-19

R39_119 V39 V119 13278.656760828568
L39_119 V39 V119 2.3368247458068943e-12
C39_119 V39 V119 5.3399882753456856e-20

R39_120 V39 V120 1901.252459731639
L39_120 V39 V120 -6.494042436060666e-11
C39_120 V39 V120 1.497672986210453e-19

R39_121 V39 V121 2323.6178126615628
L39_121 V39 V121 1.6334579513371113e-11
C39_121 V39 V121 8.169347142049552e-20

R39_122 V39 V122 32248.496894792494
L39_122 V39 V122 5.656742813732724e-12
C39_122 V39 V122 8.407649978040904e-20

R39_123 V39 V123 631.1950282123926
L39_123 V39 V123 -7.148804794111628e-13
C39_123 V39 V123 -7.817720237478881e-19

R39_124 V39 V124 1165.6103804420018
L39_124 V39 V124 2.4611416760026006e-12
C39_124 V39 V124 6.863361823144006e-20

R39_125 V39 V125 880.2974813011415
L39_125 V39 V125 2.5469594014240152e-11
C39_125 V39 V125 7.210954544569445e-20

R39_126 V39 V126 -1834.5094472234332
L39_126 V39 V126 -3.3824480815780113e-12
C39_126 V39 V126 -1.7632848748018461e-19

R39_127 V39 V127 -773.5113664555205
L39_127 V39 V127 2.8267806787579815e-12
C39_127 V39 V127 4.918190655746898e-19

R39_128 V39 V128 -1041.6889967749594
L39_128 V39 V128 -3.300849265472909e-12
C39_128 V39 V128 -1.5563777609164678e-19

R39_129 V39 V129 -746.7760662209922
L39_129 V39 V129 7.585871579126077e-12
C39_129 V39 V129 -1.3430139495185986e-19

R39_130 V39 V130 -2059.2540587703543
L39_130 V39 V130 -3.242299629458286e-11
C39_130 V39 V130 -1.623199446657419e-20

R39_131 V39 V131 1767.6218485330387
L39_131 V39 V131 1.3963639643769724e-12
C39_131 V39 V131 1.8104916598416851e-19

R39_132 V39 V132 2134.6769301396494
L39_132 V39 V132 3.207117457010718e-12
C39_132 V39 V132 2.4055585805111864e-19

R39_133 V39 V133 -1054.9695248942282
L39_133 V39 V133 -7.342057598938465e-12
C39_133 V39 V133 -1.0874089958921694e-19

R39_134 V39 V134 5662.217210167465
L39_134 V39 V134 5.269910452006982e-12
C39_134 V39 V134 1.0732653412963935e-19

R39_135 V39 V135 935.1421157192291
L39_135 V39 V135 -8.312009057326432e-13
C39_135 V39 V135 -8.754706440483065e-19

R39_136 V39 V136 1498.5695314235334
L39_136 V39 V136 2.7565325433553474e-12
C39_136 V39 V136 2.3007723508862722e-20

R39_137 V39 V137 641.7525627505769
L39_137 V39 V137 -2.5639308160423125e-12
C39_137 V39 V137 2.924063711529126e-20

R39_138 V39 V138 -7826.081693168286
L39_138 V39 V138 -3.1392935615954438e-12
C39_138 V39 V138 -1.6499701627617112e-19

R39_139 V39 V139 -479.75150917802335
L39_139 V39 V139 9.118563325892892e-13
C39_139 V39 V139 1.0012036961002576e-18

R39_140 V39 V140 -780.7410688842926
L39_140 V39 V140 -1.3954697726770026e-12
C39_140 V39 V140 -1.2768717675973596e-19

R39_141 V39 V141 933.8858783250031
L39_141 V39 V141 4.125229617677332e-12
C39_141 V39 V141 6.848491232739242e-20

R39_142 V39 V142 -3693.7784648111415
L39_142 V39 V142 -8.005579492405452e-12
C39_142 V39 V142 1.6919785206626148e-20

R39_143 V39 V143 967.4027879339014
L39_143 V39 V143 -1.2905715611678837e-10
C39_143 V39 V143 -1.2020506571996668e-19

R39_144 V39 V144 3447.580564681567
L39_144 V39 V144 6.275801138236972e-12
C39_144 V39 V144 1.136533867701966e-19

R39_145 V39 V145 -613.775755253888
L39_145 V39 V145 2.152560834505438e-12
C39_145 V39 V145 -5.0202140604485086e-20

R39_146 V39 V146 2527.4130873298764
L39_146 V39 V146 1.513793676002682e-12
C39_146 V39 V146 9.035480320950017e-20

R39_147 V39 V147 -743.0493880522637
L39_147 V39 V147 -1.7782973800990514e-12
C39_147 V39 V147 -6.560435977780121e-19

R39_148 V39 V148 3786.777092114058
L39_148 V39 V148 1.5961096245315229e-12
C39_148 V39 V148 7.901032377707755e-21

R39_149 V39 V149 -2412.908893061301
L39_149 V39 V149 1.248536973478944e-11
C39_149 V39 V149 1.9026571472623968e-19

R39_150 V39 V150 743.3758848725643
L39_150 V39 V150 -1.3748040761345948e-11
C39_150 V39 V150 2.843490536427555e-20

R39_151 V39 V151 208.3761180499656
L39_151 V39 V151 -3.582842493215642e-11
C39_151 V39 V151 3.793836852884103e-19

R39_152 V39 V152 7542.372430173012
L39_152 V39 V152 -3.1830350734178278e-12
C39_152 V39 V152 -5.861839927544092e-20

R39_153 V39 V153 2115.5736300588173
L39_153 V39 V153 -1.6896867883947352e-12
C39_153 V39 V153 -1.9745248953427153e-19

R39_154 V39 V154 -2527.642330788135
L39_154 V39 V154 -1.7119836427485551e-12
C39_154 V39 V154 -1.256110396243212e-19

R39_155 V39 V155 -98.84618665648259
L39_155 V39 V155 1.2239932538530275e-12
C39_155 V39 V155 2.407603892622712e-19

R39_156 V39 V156 1460.508467039891
L39_156 V39 V156 -3.298373874849933e-12
C39_156 V39 V156 -7.524719065193533e-20

R39_157 V39 V157 1854.8651050900535
L39_157 V39 V157 -2.5891075102314926e-12
C39_157 V39 V157 -1.691892614278658e-19

R39_158 V39 V158 2383.614570104933
L39_158 V39 V158 4.590921614407565e-12
C39_158 V39 V158 8.989268167076352e-20

R39_159 V39 V159 296.2941112280978
L39_159 V39 V159 -1.6589451281001416e-12
C39_159 V39 V159 -4.674016757711309e-19

R39_160 V39 V160 -1692.3492034463682
L39_160 V39 V160 2.2280221574753247e-11
C39_160 V39 V160 8.209761085613669e-20

R39_161 V39 V161 -16366.479371556328
L39_161 V39 V161 1.860549569731933e-12
C39_161 V39 V161 2.9333054402817683e-19

R39_162 V39 V162 31439.908351231257
L39_162 V39 V162 2.0671510758389905e-12
C39_162 V39 V162 7.846417701506677e-20

R39_163 V39 V163 400.1564681103352
L39_163 V39 V163 6.628048566198861e-12
C39_163 V39 V163 1.9784654494386744e-19

R39_164 V39 V164 698.8348008974016
L39_164 V39 V164 3.565742260287373e-12
C39_164 V39 V164 4.6029542995442284e-20

R39_165 V39 V165 2672.94687011511
L39_165 V39 V165 1.7401801150469501e-12
C39_165 V39 V165 -3.432542145706415e-20

R39_166 V39 V166 2844.0710679955223
L39_166 V39 V166 -1.0118097086884392e-11
C39_166 V39 V166 -3.250751660599709e-20

R39_167 V39 V167 -3200.2099291709983
L39_167 V39 V167 7.390954063768062e-12
C39_167 V39 V167 9.665721228281362e-20

R39_168 V39 V168 -672.9499662400481
L39_168 V39 V168 4.8762360667464754e-12
C39_168 V39 V168 1.089132282806162e-19

R39_169 V39 V169 1488.4787045528783
L39_169 V39 V169 -1.8314602353994896e-12
C39_169 V39 V169 -2.972043847103723e-19

R39_170 V39 V170 1638.497226553542
L39_170 V39 V170 -9.33889428395392e-12
C39_170 V39 V170 1.1087214922441257e-20

R39_171 V39 V171 -312.84322139263264
L39_171 V39 V171 -3.6138956610851307e-12
C39_171 V39 V171 -1.3346094066140732e-19

R39_172 V39 V172 -4297.41269162708
L39_172 V39 V172 -2.3185706898605716e-11
C39_172 V39 V172 -6.46639400015861e-20

R39_173 V39 V173 -2683.221774530306
L39_173 V39 V173 -3.5654335821533062e-12
C39_173 V39 V173 6.430734571511428e-20

R39_174 V39 V174 -619.1698282753528
L39_174 V39 V174 -1.1866082960817794e-11
C39_174 V39 V174 -1.2330241822909795e-19

R39_175 V39 V175 359.16569060779705
L39_175 V39 V175 1.8970696933298938e-12
C39_175 V39 V175 3.288823162381528e-19

R39_176 V39 V176 -50889.02588374981
L39_176 V39 V176 -2.024292123778535e-12
C39_176 V39 V176 -1.7962369693905087e-19

R39_177 V39 V177 1673.5605891811904
L39_177 V39 V177 3.8497595723345075e-12
C39_177 V39 V177 6.673096021659808e-20

R39_178 V39 V178 1073.1116401203037
L39_178 V39 V178 -6.624224841473106e-12
C39_178 V39 V178 1.7187393612402024e-20

R39_179 V39 V179 -400.94244237657205
L39_179 V39 V179 8.775018724634251e-12
C39_179 V39 V179 -3.4439232828332833e-19

R39_180 V39 V180 1901.0446792920554
L39_180 V39 V180 6.084551069014064e-12
C39_180 V39 V180 6.567694644834262e-20

R39_181 V39 V181 -3822.2823876571047
L39_181 V39 V181 6.523034553509542e-12
C39_181 V39 V181 1.0532034996167968e-19

R39_182 V39 V182 -1770.867069019665
L39_182 V39 V182 5.539918590442788e-12
C39_182 V39 V182 9.129563235891817e-20

R39_183 V39 V183 540.7332328720967
L39_183 V39 V183 -1.5600481405472493e-12
C39_183 V39 V183 2.5281958482992406e-20

R39_184 V39 V184 4487.533773913675
L39_184 V39 V184 9.250110509153768e-12
C39_184 V39 V184 -2.0267970382323978e-20

R39_185 V39 V185 -317703.21114636894
L39_185 V39 V185 3.401067470853578e-11
C39_185 V39 V185 -7.558375520623319e-20

R39_186 V39 V186 -1788.699718178843
L39_186 V39 V186 2.3871919768342055e-12
C39_186 V39 V186 -2.16578641860838e-21

R39_187 V39 V187 3051.795419745689
L39_187 V39 V187 1.3056370056885212e-12
C39_187 V39 V187 3.974039385396939e-19

R39_188 V39 V188 -556.4829061286792
L39_188 V39 V188 5.743466895975793e-12
C39_188 V39 V188 8.092361189134708e-20

R39_189 V39 V189 3049.7665140070517
L39_189 V39 V189 -3.674769599984663e-12
C39_189 V39 V189 -1.1063164803024233e-19

R39_190 V39 V190 1393.6167569021045
L39_190 V39 V190 -3.761183733199686e-12
C39_190 V39 V190 -3.8948297205169104e-20

R39_191 V39 V191 -1047.5030956953299
L39_191 V39 V191 4.7494173348962655e-12
C39_191 V39 V191 -3.201860643043272e-19

R39_192 V39 V192 2591.019938560672
L39_192 V39 V192 1.0373337976936894e-11
C39_192 V39 V192 -5.634284973065892e-20

R39_193 V39 V193 -2962.1827826560752
L39_193 V39 V193 -8.739281190574529e-11
C39_193 V39 V193 -3.446420649998522e-20

R39_194 V39 V194 -8907.987061378593
L39_194 V39 V194 -2.3845659320874057e-12
C39_194 V39 V194 -1.9073659641052782e-19

R39_195 V39 V195 1279.5287203197831
L39_195 V39 V195 -1.0252922122301942e-11
C39_195 V39 V195 4.188410891093244e-19

R39_196 V39 V196 475.1109567154006
L39_196 V39 V196 -1.3273341250277987e-12
C39_196 V39 V196 -2.3305953799974505e-19

R39_197 V39 V197 2825.7715961253202
L39_197 V39 V197 4.511836752747017e-12
C39_197 V39 V197 1.9328678787772861e-19

R39_198 V39 V198 2683.7420624649153
L39_198 V39 V198 4.189480950747034e-12
C39_198 V39 V198 1.304149136506274e-20

R39_199 V39 V199 9674.42934667552
L39_199 V39 V199 -1.223208978713622e-11
C39_199 V39 V199 -3.0696289137795774e-20

R39_200 V39 V200 -983.6030535772272
L39_200 V39 V200 2.0493224629281154e-12
C39_200 V39 V200 2.598693519559628e-19

R40_40 V40 0 -114.05352392717715
L40_40 V40 0 -8.796721500262741e-13
C40_40 V40 0 7.257046334531217e-19

R40_41 V40 V41 3775.602098930507
L40_41 V40 V41 -7.5431060658846e-12
C40_41 V40 V41 1.9189865461362476e-20

R40_42 V40 V42 8449.014056563266
L40_42 V40 V42 -1.0355897468245836e-11
C40_42 V40 V42 -3.895767044056632e-20

R40_43 V40 V43 4307.133035175748
L40_43 V40 V43 -2.136439752227269e-11
C40_43 V40 V43 9.859555210096622e-20

R40_44 V40 V44 4679.000479787102
L40_44 V40 V44 1.8484276320428453e-11
C40_44 V40 V44 2.7443509428243356e-19

R40_45 V40 V45 2984.0796210754925
L40_45 V40 V45 4.933489659222802e-12
C40_45 V40 V45 -3.857719394399093e-20

R40_46 V40 V46 3583.815355743841
L40_46 V40 V46 -7.225948511384569e-12
C40_46 V40 V46 -1.919314102512049e-19

R40_47 V40 V47 1576.5237377190165
L40_47 V40 V47 1.3848804147345003e-11
C40_47 V40 V47 -3.632734342504149e-21

R40_48 V40 V48 575.8041474574661
L40_48 V40 V48 1.5808387221510202e-12
C40_48 V40 V48 3.3531801591809683e-19

R40_49 V40 V49 -79315.00040752326
L40_49 V40 V49 1.4491731242730103e-11
C40_49 V40 V49 -8.798532790082388e-20

R40_50 V40 V50 -151875.90905478568
L40_50 V40 V50 7.1271345738776685e-12
C40_50 V40 V50 9.079683560490085e-20

R40_51 V40 V51 4456.335165698724
L40_51 V40 V51 6.2632886464706615e-12
C40_51 V40 V51 -6.490383247961403e-21

R40_52 V40 V52 -20952.345841162292
L40_52 V40 V52 -1.3324581553853813e-12
C40_52 V40 V52 -4.2491956801866234e-19

R40_53 V40 V53 4343.3426304776085
L40_53 V40 V53 1.4370513687379477e-12
C40_53 V40 V53 3.2967070214384996e-19

R40_54 V40 V54 -19049.42527785939
L40_54 V40 V54 3.81202334832837e-12
C40_54 V40 V54 1.8780702835785022e-19

R40_55 V40 V55 -15883.047689023568
L40_55 V40 V55 3.293809061854674e-12
C40_55 V40 V55 1.945703649433561e-19

R40_56 V40 V56 -1040.1157109977441
L40_56 V40 V56 1.973286019052494e-12
C40_56 V40 V56 3.749755375595222e-19

R40_57 V40 V57 -4177.454355233352
L40_57 V40 V57 -1.3850447576714094e-12
C40_57 V40 V57 -3.6191847012303076e-19

R40_58 V40 V58 2299.8704311290126
L40_58 V40 V58 -4.90336364344561e-12
C40_58 V40 V58 -1.4094515302047533e-19

R40_59 V40 V59 -2614.7795297947787
L40_59 V40 V59 -3.479667930628445e-12
C40_59 V40 V59 -1.9387943439131657e-19

R40_60 V40 V60 -1180.4671927203183
L40_60 V40 V60 -5.537284526210717e-12
C40_60 V40 V60 -1.132153773829367e-19

R40_61 V40 V61 7272.029665754991
L40_61 V40 V61 2.4843082076932333e-10
C40_61 V40 V61 -9.297989373225613e-21

R40_62 V40 V62 -2332.217991124928
L40_62 V40 V62 -5.2407849154033206e-12
C40_62 V40 V62 -1.6835562768614007e-19

R40_63 V40 V63 11312.005771617985
L40_63 V40 V63 -5.2229426363888536e-12
C40_63 V40 V63 -6.958738762267459e-20

R40_64 V40 V64 2947.902333669046
L40_64 V40 V64 -7.841625687936872e-12
C40_64 V40 V64 -5.869540672020321e-20

R40_65 V40 V65 4072.632829333254
L40_65 V40 V65 4.042749720840692e-12
C40_65 V40 V65 9.270675580314894e-20

R40_66 V40 V66 16397.479260906344
L40_66 V40 V66 5.729276370590786e-12
C40_66 V40 V66 7.970772095316012e-20

R40_67 V40 V67 7236.901953474968
L40_67 V40 V67 3.0183875757282746e-12
C40_67 V40 V67 1.787864301885778e-19

R40_68 V40 V68 1277.640594446393
L40_68 V40 V68 -2.4991850975720877e-11
C40_68 V40 V68 7.727169174922256e-20

R40_69 V40 V69 -19459.160052920848
L40_69 V40 V69 3.0790318816397537e-12
C40_69 V40 V69 1.0545564028203663e-19

R40_70 V40 V70 4338.424467350046
L40_70 V40 V70 1.6715335115616288e-11
C40_70 V40 V70 5.501078151743478e-20

R40_71 V40 V71 3726.9308539327826
L40_71 V40 V71 -3.190357404804821e-11
C40_71 V40 V71 -7.828733835448673e-20

R40_72 V40 V72 1191.7937446392482
L40_72 V40 V72 -1.0495702258162382e-10
C40_72 V40 V72 -7.447038416575279e-20

R40_73 V40 V73 3075.3792394428096
L40_73 V40 V73 -3.1370851237937467e-11
C40_73 V40 V73 -8.567583186615157e-20

R40_74 V40 V74 -3983.2063562904023
L40_74 V40 V74 -5.738248573636979e-12
C40_74 V40 V74 -1.3793657621714523e-19

R40_75 V40 V75 -93094.2968679355
L40_75 V40 V75 -5.110546677790932e-12
C40_75 V40 V75 -7.706699931744727e-20

R40_76 V40 V76 -631.023623787741
L40_76 V40 V76 1.510535185707534e-12
C40_76 V40 V76 3.4865143018891035e-19

R40_77 V40 V77 -3318.1743166765764
L40_77 V40 V77 -2.5693931714437074e-12
C40_77 V40 V77 -1.9479338294752173e-19

R40_78 V40 V78 2804.794109571706
L40_78 V40 V78 3.633682687672663e-12
C40_78 V40 V78 2.3430772290240897e-19

R40_79 V40 V79 -1585.1015650986344
L40_79 V40 V79 4.1343848619842274e-12
C40_79 V40 V79 7.433488112398954e-20

R40_80 V40 V80 -1662.8660862032982
L40_80 V40 V80 -1.6781856559095886e-12
C40_80 V40 V80 -3.305373964547764e-19

R40_81 V40 V81 2726.216216809976
L40_81 V40 V81 4.419687184365988e-12
C40_81 V40 V81 4.7606572715704945e-20

R40_82 V40 V82 -5952.646993147659
L40_82 V40 V82 -5.873927383459863e-12
C40_82 V40 V82 -2.0404682860685999e-19

R40_83 V40 V83 3637.976055067449
L40_83 V40 V83 -6.288675592497103e-12
C40_83 V40 V83 -8.307164330674022e-20

R40_84 V40 V84 1469.7421131203457
L40_84 V40 V84 -2.1038218466435407e-12
C40_84 V40 V84 -2.3316707303235773e-19

R40_85 V40 V85 -21394.12921488334
L40_85 V40 V85 6.714015046098866e-11
C40_85 V40 V85 -1.59566089213992e-20

R40_86 V40 V86 2937.7430808632635
L40_86 V40 V86 -3.099433939667818e-12
C40_86 V40 V86 -2.1055834851858608e-19

R40_87 V40 V87 1766.6016303569556
L40_87 V40 V87 5.319203143409169e-11
C40_87 V40 V87 1.4961681870416199e-19

R40_88 V40 V88 591.508393503449
L40_88 V40 V88 1.1354923915550431e-12
C40_88 V40 V88 6.632654689065467e-19

R40_89 V40 V89 3448.308575055098
L40_89 V40 V89 1.6770645465295976e-12
C40_89 V40 V89 2.9828093281558096e-19

R40_90 V40 V90 11925.927595918763
L40_90 V40 V90 1.7490245990824533e-12
C40_90 V40 V90 4.9109052048470795e-19

R40_91 V40 V91 8678.946566729821
L40_91 V40 V91 6.846035743077204e-12
C40_91 V40 V91 -1.4525236861289115e-19

R40_92 V40 V92 -527.6263294295536
L40_92 V40 V92 -1.3497838338013093e-12
C40_92 V40 V92 -5.08223776951691e-19

R40_93 V40 V93 2531.230951145016
L40_93 V40 V93 -4.088713922785908e-12
C40_93 V40 V93 -9.369889267867994e-20

R40_94 V40 V94 -5278.274690791983
L40_94 V40 V94 5.5745961024918116e-12
C40_94 V40 V94 -3.9364545045783024e-20

R40_95 V40 V95 -1041.8400836685014
L40_95 V40 V95 -9.723278103802561e-12
C40_95 V40 V95 -1.0290447626006452e-19

R40_96 V40 V96 -403.67695775690964
L40_96 V40 V96 -2.5704390993932736e-10
C40_96 V40 V96 -3.0358206746529855e-19

R40_97 V40 V97 -1003.8780414459819
L40_97 V40 V97 -1.8171782989513082e-12
C40_97 V40 V97 -5.64406703105939e-19

R40_98 V40 V98 12855.937201952256
L40_98 V40 V98 -1.451089043671603e-12
C40_98 V40 V98 -4.273480429830161e-19

R40_99 V40 V99 1619.9980098665826
L40_99 V40 V99 1.1632417516074928e-11
C40_99 V40 V99 2.577105824002685e-19

R40_100 V40 V100 244.72432148917434
L40_100 V40 V100 2.3338022441592204e-12
C40_100 V40 V100 5.959123195894503e-19

R40_101 V40 V101 2421.749447374144
L40_101 V40 V101 1.668684744801623e-12
C40_101 V40 V101 3.81049748255489e-19

R40_102 V40 V102 -5075.187440326473
L40_102 V40 V102 -1.2313372064387827e-11
C40_102 V40 V102 8.808649976567615e-20

R40_103 V40 V103 3146.140488430036
L40_103 V40 V103 -7.188234086255653e-12
C40_103 V40 V103 -1.0452675570948378e-19

R40_104 V40 V104 -1498.5532374560319
L40_104 V40 V104 -2.007249797583978e-12
C40_104 V40 V104 -1.0329056704174215e-19

R40_105 V40 V105 761.3540203874023
L40_105 V40 V105 3.7694371745493975e-12
C40_105 V40 V105 2.481162891795403e-19

R40_106 V40 V106 649.0266421877855
L40_106 V40 V106 1.5445069829781614e-12
C40_106 V40 V106 4.647800255094777e-19

R40_107 V40 V107 -6512.283138060533
L40_107 V40 V107 1.973416245033856e-11
C40_107 V40 V107 -8.7884391966639e-20

R40_108 V40 V108 -480.378108506957
L40_108 V40 V108 2.52547312132258e-12
C40_108 V40 V108 -7.231048487501326e-20

R40_109 V40 V109 -1033.9776751187858
L40_109 V40 V109 -4.464608327851327e-12
C40_109 V40 V109 -3.520464246366963e-19

R40_110 V40 V110 -743.7355632416755
L40_110 V40 V110 -6.122843966131958e-12
C40_110 V40 V110 -1.9422364156539925e-19

R40_111 V40 V111 869.0722845960331
L40_111 V40 V111 4.555840282722039e-12
C40_111 V40 V111 7.916553478474722e-20

R40_112 V40 V112 367.5589215140653
L40_112 V40 V112 -1.5090597838243e-12
C40_112 V40 V112 -4.261732526756119e-19

R40_113 V40 V113 -1788.5624802336692
L40_113 V40 V113 -6.274320228606262e-12
C40_113 V40 V113 -2.1641547003582427e-19

R40_114 V40 V114 -772.0383939596884
L40_114 V40 V114 -1.4899991402011405e-12
C40_114 V40 V114 -4.346245942403934e-19

R40_115 V40 V115 -514.9029594786568
L40_115 V40 V115 -3.3988384944728923e-12
C40_115 V40 V115 -4.7344968887330904e-20

R40_116 V40 V116 -879.0422749744129
L40_116 V40 V116 2.4606426404828264e-12
C40_116 V40 V116 3.5586083484926533e-19

R40_117 V40 V117 -42327.33281258229
L40_117 V40 V117 1.2199590766064502e-11
C40_117 V40 V117 1.8143534499246058e-19

R40_118 V40 V118 418.22232080928654
L40_118 V40 V118 3.4572700458006434e-12
C40_118 V40 V118 3.597262079529096e-19

R40_119 V40 V119 1272.178469294066
L40_119 V40 V119 5.784392976803784e-12
C40_119 V40 V119 2.324936713112165e-19

R40_120 V40 V120 2250.1367820231744
L40_120 V40 V120 1.8618033664771045e-12
C40_120 V40 V120 4.383198861238286e-19

R40_121 V40 V121 5677.190006873091
L40_121 V40 V121 3.530585911459024e-12
C40_121 V40 V121 1.198360016267539e-19

R40_122 V40 V122 -2909.4707459853653
L40_122 V40 V122 3.4857432991148185e-12
C40_122 V40 V122 1.2557303825356415e-19

R40_123 V40 V123 826.8657826107813
L40_123 V40 V123 1.6923827086580895e-11
C40_123 V40 V123 -1.7790444088434211e-19

R40_124 V40 V124 1107.0314757968683
L40_124 V40 V124 -6.494324996256164e-13
C40_124 V40 V124 -1.0996543360825664e-18

R40_125 V40 V125 667.7233290118544
L40_125 V40 V125 -8.098907213540081e-11
C40_125 V40 V125 3.727680783922037e-20

R40_126 V40 V126 -1148.850227020821
L40_126 V40 V126 -2.434940842237737e-12
C40_126 V40 V126 -2.0522536622098843e-19

R40_127 V40 V127 -544.7479536671154
L40_127 V40 V127 -2.202307948910577e-12
C40_127 V40 V127 -1.951008686376865e-19

R40_128 V40 V128 -623.543282430102
L40_128 V40 V128 3.0472905168106526e-12
C40_128 V40 V128 3.0170585336281535e-19

R40_129 V40 V129 -564.1716455600478
L40_129 V40 V129 9.201030836063021e-12
C40_129 V40 V129 -1.7855181832232512e-19

R40_130 V40 V130 -2774.810299905771
L40_130 V40 V130 -2.993709954092246e-11
C40_130 V40 V130 2.50659556663351e-21

R40_131 V40 V131 706.6610356017079
L40_131 V40 V131 2.7025412473398484e-12
C40_131 V40 V131 2.854093089963476e-19

R40_132 V40 V132 659.8769065931884
L40_132 V40 V132 1.0867490145896933e-12
C40_132 V40 V132 5.474762848676509e-19

R40_133 V40 V133 -1039.647589721514
L40_133 V40 V133 -8.575047089010736e-12
C40_133 V40 V133 -2.1723933438828877e-20

R40_134 V40 V134 1717.452828220236
L40_134 V40 V134 3.447101504463572e-12
C40_134 V40 V134 2.491730621436354e-19

R40_135 V40 V135 2599.804584454189
L40_135 V40 V135 5.147341173094881e-12
C40_135 V40 V135 -3.8705533282254053e-20

R40_136 V40 V136 771.4749439188605
L40_136 V40 V136 -1.0923335580288037e-12
C40_136 V40 V136 -8.861302634591942e-19

R40_137 V40 V137 536.1697773574108
L40_137 V40 V137 -1.6664096281325705e-12
C40_137 V40 V137 -6.081533714948544e-20

R40_138 V40 V138 -1697.0513688767699
L40_138 V40 V138 -2.561229910392451e-12
C40_138 V40 V138 -2.7724760690719743e-19

R40_139 V40 V139 -450.27380786350153
L40_139 V40 V139 -2.0767651433120673e-12
C40_139 V40 V139 -3.0411533818019354e-20

R40_140 V40 V140 -520.4273078732481
L40_140 V40 V140 6.830695443232147e-12
C40_140 V40 V140 7.60940431678802e-19

R40_141 V40 V141 913.863787392651
L40_141 V40 V141 2.9695059167119475e-12
C40_141 V40 V141 5.483485197429332e-20

R40_142 V40 V142 -1195.391093548302
L40_142 V40 V142 -4.873764580449085e-12
C40_142 V40 V142 -1.9287335223555505e-20

R40_143 V40 V143 658.2473756025323
L40_143 V40 V143 -2.023368827432312e-11
C40_143 V40 V143 -5.4665111977742e-20

R40_144 V40 V144 -476.3272705570043
L40_144 V40 V144 2.3397802100656055e-12
C40_144 V40 V144 -3.165887166269291e-20

R40_145 V40 V145 -478.86255122265646
L40_145 V40 V145 1.4158685099247764e-12
C40_145 V40 V145 3.0775479532597444e-21

R40_146 V40 V146 1324.9948980461788
L40_146 V40 V146 1.0262790590273556e-12
C40_146 V40 V146 1.4735176173538417e-19

R40_147 V40 V147 -820.3347675258038
L40_147 V40 V147 3.4853180707262615e-12
C40_147 V40 V147 -1.4363652139668376e-19

R40_148 V40 V148 181.19948725784784
L40_148 V40 V148 -1.1395403558001178e-12
C40_148 V40 V148 -5.360992218315246e-19

R40_149 V40 V149 -3468.0664549443836
L40_149 V40 V149 -3.616595920534765e-11
C40_149 V40 V149 2.1225158503373267e-19

R40_150 V40 V150 455.30743913947646
L40_150 V40 V150 -3.815377582155208e-12
C40_150 V40 V150 -2.4346083713517e-20

R40_151 V40 V151 540.8096310553381
L40_151 V40 V151 5.2020281439607955e-12
C40_151 V40 V151 1.0375977740491122e-19

R40_152 V40 V152 -1007.8656341866968
L40_152 V40 V152 2.6112933566856503e-12
C40_152 V40 V152 1.8532422861175913e-19

R40_153 V40 V153 4061.385931713372
L40_153 V40 V153 -1.8405916668050345e-12
C40_153 V40 V153 -1.8580984292953778e-19

R40_154 V40 V154 -588.7445700148278
L40_154 V40 V154 -2.370664753598907e-12
C40_154 V40 V154 -1.2030112777563086e-19

R40_155 V40 V155 -202.23649624364833
L40_155 V40 V155 -6.299301287320243e-12
C40_155 V40 V155 1.0157597717190174e-19

R40_156 V40 V156 -52171.13493345733
L40_156 V40 V156 -3.892861749598953e-12
C40_156 V40 V156 3.7917582347997947e-19

R40_157 V40 V157 796.2164929052537
L40_157 V40 V157 -1.3235846801403075e-12
C40_157 V40 V157 -3.4508823621169173e-19

R40_158 V40 V158 757.8305530702127
L40_158 V40 V158 1.2750106932575878e-11
C40_158 V40 V158 1.0253250105316722e-19

R40_159 V40 V159 293.77549234033023
L40_159 V40 V159 -6.374372772464013e-12
C40_159 V40 V159 -6.066688842189619e-20

R40_160 V40 V160 -336.5946912495053
L40_160 V40 V160 4.8591562144277677e-11
C40_160 V40 V160 -3.7889682379983844e-19

R40_161 V40 V161 -1838.1187057502045
L40_161 V40 V161 1.1231575452736788e-12
C40_161 V40 V161 4.0404487382548393e-19

R40_162 V40 V162 -32047.938600420486
L40_162 V40 V162 1.6569222385878514e-12
C40_162 V40 V162 7.591610911175749e-20

R40_163 V40 V163 2090.9432157067918
L40_163 V40 V163 1.1137350871692287e-11
C40_163 V40 V163 -1.5964228685678492e-20

R40_164 V40 V164 160.71752747247442
L40_164 V40 V164 5.294467241164455e-12
C40_164 V40 V164 2.7752880317741517e-19

R40_165 V40 V165 756.3532683371006
L40_165 V40 V165 1.5647935894490018e-12
C40_165 V40 V165 1.2005961732595788e-20

R40_166 V40 V166 1269.677243715879
L40_166 V40 V166 -5.577824377948187e-12
C40_166 V40 V166 -8.427485854250956e-20

R40_167 V40 V167 602.5010391708008
L40_167 V40 V167 3.865701256229319e-12
C40_167 V40 V167 1.4852081244059235e-19

R40_168 V40 V168 -179.55121299595527
L40_168 V40 V168 1.7818915729600574e-12
C40_168 V40 V168 1.154063480401833e-19

R40_169 V40 V169 1549.8739387903133
L40_169 V40 V169 -1.6298687251703623e-12
C40_169 V40 V169 -3.8495788768105146e-19

R40_170 V40 V170 2346.1094159211993
L40_170 V40 V170 2.177467017858734e-11
C40_170 V40 V170 7.223884054846827e-20

R40_171 V40 V171 -490.5083757760138
L40_171 V40 V171 3.3327572328393527e-12
C40_171 V40 V171 3.7431872466469183e-20

R40_172 V40 V172 -1550.113739564079
L40_172 V40 V172 -1.1406278085099113e-12
C40_172 V40 V172 -1.9694321847340798e-19

R40_173 V40 V173 -1583.4202285394265
L40_173 V40 V173 -2.5236845829025086e-12
C40_173 V40 V173 4.9105470467517044e-20

R40_174 V40 V174 -452.3199207165441
L40_174 V40 V174 -3.958406058109442e-12
C40_174 V40 V174 -1.7823023718075839e-19

R40_175 V40 V175 2604.1806204875047
L40_175 V40 V175 -1.6152230327442642e-12
C40_175 V40 V175 -1.241588897537173e-19

R40_176 V40 V176 357.51983099029286
L40_176 V40 V176 2.504426272101637e-12
C40_176 V40 V176 3.2983731044552237e-19

R40_177 V40 V177 978.4036548248122
L40_177 V40 V177 2.925176338827565e-12
C40_177 V40 V177 1.0213786193901398e-19

R40_178 V40 V178 707.9725148590122
L40_178 V40 V178 -4.401734884842475e-12
C40_178 V40 V178 -1.4334992606134818e-20

R40_179 V40 V179 -2510.564858309286
L40_179 V40 V179 -9.584131854265752e-12
C40_179 V40 V179 -9.634158361355008e-20

R40_180 V40 V180 -909.9376850241371
L40_180 V40 V180 3.156844757142985e-12
C40_180 V40 V180 -3.631739006805716e-19

R40_181 V40 V181 -2176.9266499995265
L40_181 V40 V181 1.006704246283557e-11
C40_181 V40 V181 1.2472894760733729e-19

R40_182 V40 V182 -1142.9747666632227
L40_182 V40 V182 1.1147484933059784e-11
C40_182 V40 V182 5.448732899683108e-20

R40_183 V40 V183 930.9428259593482
L40_183 V40 V183 -2.6368838724606866e-11
C40_183 V40 V183 -8.07896638138734e-20

R40_184 V40 V184 1705.915378572036
L40_184 V40 V184 -1.8105290999701153e-12
C40_184 V40 V184 7.244083815690689e-20

R40_185 V40 V185 19659.72963095544
L40_185 V40 V185 2.210649040162554e-11
C40_185 V40 V185 -9.724931112673836e-20

R40_186 V40 V186 -1972.9588763783067
L40_186 V40 V186 2.802314136806842e-12
C40_186 V40 V186 1.0606338501184007e-19

R40_187 V40 V187 -1303.0428508211075
L40_187 V40 V187 3.906076156708663e-12
C40_187 V40 V187 1.7801665455896335e-19

R40_188 V40 V188 -486.1328046564879
L40_188 V40 V188 8.195853238230433e-13
C40_188 V40 V188 3.6939581995348385e-19

R40_189 V40 V189 4892.832168925453
L40_189 V40 V189 -2.8300440497327757e-12
C40_189 V40 V189 -1.1576302631616587e-19

R40_190 V40 V190 886.6407571954078
L40_190 V40 V190 -4.194699564125751e-12
C40_190 V40 V190 -3.7357986479493414e-20

R40_191 V40 V191 -1833.8688506658523
L40_191 V40 V191 2.27478616392833e-12
C40_191 V40 V191 6.485783929153867e-20

R40_192 V40 V192 -36131.33687952002
L40_192 V40 V192 -1.8060914324725043e-12
C40_192 V40 V192 -4.778743705157364e-19

R40_193 V40 V193 -1132.6543194240219
L40_193 V40 V193 -9.08909587552651e-12
C40_193 V40 V193 -1.4649853406365687e-19

R40_194 V40 V194 7442.728376368231
L40_194 V40 V194 -1.1812492309072942e-12
C40_194 V40 V194 -3.740237717598474e-19

R40_195 V40 V195 766.718475146044
L40_195 V40 V195 -1.2475898611509565e-12
C40_195 V40 V195 -2.944965868066254e-19

R40_196 V40 V196 377.7493398509269
L40_196 V40 V196 2.849947665438457e-12
C40_196 V40 V196 5.935792924155473e-19

R40_197 V40 V197 8886.050601601757
L40_197 V40 V197 3.0939034004462037e-12
C40_197 V40 V197 2.646859733149044e-19

R40_198 V40 V198 1347.888981803845
L40_198 V40 V198 3.818304948758801e-12
C40_198 V40 V198 -1.6768224689119878e-20

R40_199 V40 V199 460.37681191934325
L40_199 V40 V199 4.41767018762787e-12
C40_199 V40 V199 1.099353072204779e-19

R40_200 V40 V200 -352.90316766054616
L40_200 V40 V200 -2.6817570161628183e-10
C40_200 V40 V200 -5.192574227118494e-20

R41_41 V41 0 -2053.662573114257
L41_41 V41 0 2.8784110725341106e-12
C41_41 V41 0 8.847816732914868e-19

R41_42 V41 V42 -9790.957072809537
L41_42 V41 V42 -3.756834057166959e-12
C41_42 V41 V42 -2.2824710181199103e-19

R41_43 V41 V43 -7495.5689814467505
L41_43 V41 V43 -4.926709384835896e-12
C41_43 V41 V43 -1.6111360855160173e-19

R41_44 V41 V44 -5338.163884302913
L41_44 V41 V44 -2.9547571295316853e-12
C41_44 V41 V44 -2.391559525927284e-19

R41_45 V41 V45 4224.787928146793
L41_45 V41 V45 4.8548708651167576e-12
C41_45 V41 V45 -3.8162438202222246e-20

R41_46 V41 V46 -5793.385099146412
L41_46 V41 V46 -4.625545397784402e-12
C41_46 V41 V46 -1.3733847667671409e-19

R41_47 V41 V47 -4951.952571974019
L41_47 V41 V47 8.503640830777728e-11
C41_47 V41 V47 1.4988751187681237e-20

R41_48 V41 V48 -3578.549727261995
L41_48 V41 V48 -1.8134445543581743e-11
C41_48 V41 V48 -4.5947003415708815e-20

R41_49 V41 V49 4203.879873166138
L41_49 V41 V49 1.5064264337791995e-12
C41_49 V41 V49 3.935618515415529e-19

R41_50 V41 V50 -22910.533439052644
L41_50 V41 V50 2.294285805582417e-12
C41_50 V41 V50 2.2085420221716223e-19

R41_51 V41 V51 -25427.468098280664
L41_51 V41 V51 5.683814543175202e-12
C41_51 V41 V51 6.668622351085283e-20

R41_52 V41 V52 39211.19569668282
L41_52 V41 V52 5.1367255125648665e-12
C41_52 V41 V52 1.3731573213525112e-19

R41_53 V41 V53 2990.459771142008
L41_53 V41 V53 -6.894561323579137e-12
C41_53 V41 V53 -1.761907042223629e-19

R41_54 V41 V54 4718.471698739711
L41_54 V41 V54 1.0101872512971647e-11
C41_54 V41 V54 3.3012898621957167e-20

R41_55 V41 V55 5848.301089795067
L41_55 V41 V55 1.901404628460361e-11
C41_55 V41 V55 -1.0259355244965665e-20

R41_56 V41 V56 3155.133998605168
L41_56 V41 V56 8.334240766797076e-12
C41_56 V41 V56 7.519229575578563e-20

R41_57 V41 V57 54023.47186983308
L41_57 V41 V57 -3.376074318941479e-12
C41_57 V41 V57 1.5855154766832165e-19

R41_58 V41 V58 -4652.796910744787
L41_58 V41 V58 -4.559624692743573e-12
C41_58 V41 V58 -1.0851308540299386e-19

R41_59 V41 V59 -22439.589368454188
L41_59 V41 V59 -5.479538797202871e-12
C41_59 V41 V59 -7.637404339374336e-20

R41_60 V41 V60 -17568.44627249663
L41_60 V41 V60 -3.7177179613678346e-12
C41_60 V41 V60 -8.330799121873161e-20

R41_61 V41 V61 -3236.2272183263935
L41_61 V41 V61 8.150804584564684e-12
C41_61 V41 V61 -1.3755631592748314e-19

R41_62 V41 V62 16489.968344925022
L41_62 V41 V62 -1.160983063201935e-10
C41_62 V41 V62 6.1387002821075046e-21

R41_63 V41 V63 -19766.47791874335
L41_63 V41 V63 1.5127921575862116e-10
C41_63 V41 V63 4.1894355739295526e-20

R41_64 V41 V64 -7731.612205648452
L41_64 V41 V64 -2.2578172729017483e-11
C41_64 V41 V64 2.0283822331162523e-21

R41_65 V41 V65 -23729.618584159558
L41_65 V41 V65 -1.7291733733261022e-10
C41_65 V41 V65 -1.129840396209305e-19

R41_66 V41 V66 -12478.984183289931
L41_66 V41 V66 9.653381818600622e-12
C41_66 V41 V66 1.0055836395543582e-20

R41_67 V41 V67 -155198.57152996655
L41_67 V41 V67 5.821248882807659e-12
C41_67 V41 V67 6.678326218381383e-20

R41_68 V41 V68 -12476.607728239636
L41_68 V41 V68 9.86186844917308e-12
C41_68 V41 V68 -4.253262943103399e-21

R41_69 V41 V69 2619.430843652509
L41_69 V41 V69 7.538841196101354e-12
C41_69 V41 V69 7.949849485446945e-20

R41_70 V41 V70 -9422.578650919548
L41_70 V41 V70 1.7512822188142547e-11
C41_70 V41 V70 3.8396389896536255e-21

R41_71 V41 V71 -6181.216221628444
L41_71 V41 V71 -2.0640813937388458e-11
C41_71 V41 V71 -7.538976322822394e-20

R41_72 V41 V72 -6494.096501878071
L41_72 V41 V72 1.907734342088907e-11
C41_72 V41 V72 -9.582203559051457e-21

R41_73 V41 V73 26309.126053688262
L41_73 V41 V73 -2.259669146059349e-11
C41_73 V41 V73 -5.0372037388354076e-20

R41_74 V41 V74 5972.305886976112
L41_74 V41 V74 7.946829876168818e-11
C41_74 V41 V74 2.987231805298818e-21

R41_75 V41 V75 30383.774521753592
L41_75 V41 V75 -7.801217008962086e-12
C41_75 V41 V75 -9.011796823135784e-20

R41_76 V41 V76 3833.1989796835355
L41_76 V41 V76 1.1968623153188337e-10
C41_76 V41 V76 3.645076284099721e-20

R41_77 V41 V77 -9957.256012467393
L41_77 V41 V77 3.2971976043355354e-11
C41_77 V41 V77 1.7354498917174856e-19

R41_78 V41 V78 -22615.649415274424
L41_78 V41 V78 -1.7608624258667134e-11
C41_78 V41 V78 -6.353714124874721e-21

R41_79 V41 V79 4897.92170107097
L41_79 V41 V79 7.664836142032765e-11
C41_79 V41 V79 7.897303682766169e-20

R41_80 V41 V80 15060.124289398578
L41_80 V41 V80 -6.170378128468649e-12
C41_80 V41 V80 -1.1455939281920095e-20

R41_81 V41 V81 3348.8403313376407
L41_81 V41 V81 9.674299866479473e-12
C41_81 V41 V81 -5.525048240636283e-20

R41_82 V41 V82 -21913.22481575344
L41_82 V41 V82 2.2279602444574734e-11
C41_82 V41 V82 1.703934245461502e-20

R41_83 V41 V83 -7192.991576307244
L41_83 V41 V83 5.600371328249259e-12
C41_83 V41 V83 1.0769962519924878e-19

R41_84 V41 V84 -4711.597765967575
L41_84 V41 V84 3.7640402791578143e-11
C41_84 V41 V84 4.0627418981489355e-20

R41_85 V41 V85 -5088.702381435464
L41_85 V41 V85 -2.9606962390185e-12
C41_85 V41 V85 -3.1005924419381816e-19

R41_86 V41 V86 -2561.9037066618243
L41_86 V41 V86 1.9392676290664925e-11
C41_86 V41 V86 -5.81298106746743e-20

R41_87 V41 V87 -4613.384114607351
L41_87 V41 V87 -8.914206523587625e-11
C41_87 V41 V87 -3.564424463718955e-20

R41_88 V41 V88 -5039.853957050435
L41_88 V41 V88 7.978379534401714e-12
C41_88 V41 V88 1.0724105091540218e-20

R41_89 V41 V89 11228.859245749994
L41_89 V41 V89 2.3029057279755547e-12
C41_89 V41 V89 1.1199083496862348e-19

R41_90 V41 V90 3276.880427225503
L41_90 V41 V90 6.368368297367183e-12
C41_90 V41 V90 8.272037763217761e-20

R41_91 V41 V91 10699.598551292633
L41_91 V41 V91 -4.104156194905063e-12
C41_91 V41 V91 -2.0040421875562345e-19

R41_92 V41 V92 4962.884304828001
L41_92 V41 V92 -3.8989076941871e-12
C41_92 V41 V92 -1.3109593175506519e-19

R41_93 V41 V93 3304.675240300756
L41_93 V41 V93 -3.4925235472658917e-11
C41_93 V41 V93 2.3302489313167976e-19

R41_94 V41 V94 4084.5638670711655
L41_94 V41 V94 -5.110822916957385e-12
C41_94 V41 V94 -7.340848297955112e-21

R41_95 V41 V95 3327.6996008506308
L41_95 V41 V95 2.6867664300783985e-11
C41_95 V41 V95 6.977549008483065e-20

R41_96 V41 V96 2457.5483770490196
L41_96 V41 V96 1.602987114185374e-11
C41_96 V41 V96 6.562305140180684e-20

R41_97 V41 V97 4104.215754259812
L41_97 V41 V97 -1.7324997504893634e-12
C41_97 V41 V97 -1.5344862638296054e-19

R41_98 V41 V98 -2071.173891428288
L41_98 V41 V98 1.1500923378425881e-11
C41_98 V41 V98 -6.409579797669964e-20

R41_99 V41 V99 -3027.3870724148046
L41_99 V41 V99 3.872758291555693e-12
C41_99 V41 V99 2.1608400954941361e-19

R41_100 V41 V100 -1794.971728346746
L41_100 V41 V100 3.988387513270962e-11
C41_100 V41 V100 1.66188752465001e-19

R41_101 V41 V101 -2916.681509489405
L41_101 V41 V101 1.5992890538798953e-12
C41_101 V41 V101 -4.402277138641987e-20

R41_102 V41 V102 13893.95204608336
L41_102 V41 V102 7.434223916828488e-12
C41_102 V41 V102 6.543628356711293e-20

R41_103 V41 V103 -8573.891567390412
L41_103 V41 V103 -2.0340526905809462e-11
C41_103 V41 V103 -7.056976799689539e-20

R41_104 V41 V104 -5398.88440610504
L41_104 V41 V104 -9.885162790051795e-12
C41_104 V41 V104 -1.134870247235078e-19

R41_105 V41 V105 3091.413087331448
L41_105 V41 V105 1.2380987757537107e-11
C41_105 V41 V105 1.6377985110566802e-20

R41_106 V41 V106 -3484.073821681666
L41_106 V41 V106 -5.624459732362902e-12
C41_106 V41 V106 1.559982237730819e-20

R41_107 V41 V107 57811.647945814126
L41_107 V41 V107 -5.910052189143199e-12
C41_107 V41 V107 -1.759714905623855e-19

R41_108 V41 V108 3692.733492367367
L41_108 V41 V108 6.927470952499022e-12
C41_108 V41 V108 -7.851191986041517e-20

R41_109 V41 V109 7839.425945161749
L41_109 V41 V109 -3.3374132685361404e-12
C41_109 V41 V109 -1.14921505994972e-19

R41_110 V41 V110 3434.6470535732365
L41_110 V41 V110 7.827033066719217e-12
C41_110 V41 V110 -2.844506290624407e-20

R41_111 V41 V111 -6049.976381181031
L41_111 V41 V111 -1.727415175731718e-11
C41_111 V41 V111 5.918485354420615e-21

R41_112 V41 V112 -5801.52900270347
L41_112 V41 V112 -5.50613551569535e-12
C41_112 V41 V112 1.8055916450082008e-21

R41_113 V41 V113 -18373.523712634444
L41_113 V41 V113 -4.772666454533126e-10
C41_113 V41 V113 8.448073618748161e-20

R41_114 V41 V114 4694.323190917591
L41_114 V41 V114 -1.4134681118363196e-11
C41_114 V41 V114 -4.7995625480643826e-20

R41_115 V41 V115 2492.2318514035956
L41_115 V41 V115 3.4340804340532592e-12
C41_115 V41 V115 1.8078759405220027e-19

R41_116 V41 V116 5015.630202127108
L41_116 V41 V116 6.1578986741230115e-12
C41_116 V41 V116 1.3685194214024125e-19

R41_117 V41 V117 1786.2539603957173
L41_117 V41 V117 8.294448641833319e-12
C41_117 V41 V117 1.0110067532420945e-19

R41_118 V41 V118 -2055.946255163028
L41_118 V41 V118 1.0376023040416148e-10
C41_118 V41 V118 1.0806371904488256e-19

R41_119 V41 V119 -3782.1441119885158
L41_119 V41 V119 4.914308951174084e-11
C41_119 V41 V119 -1.984571441724148e-20

R41_120 V41 V120 -3378.258301632466
L41_120 V41 V120 5.828628613640826e-12
C41_120 V41 V120 2.7797982473441224e-20

R41_121 V41 V121 -4327.5717945903925
L41_121 V41 V121 1.2126975163964325e-11
C41_121 V41 V121 -8.034053499658293e-20

R41_122 V41 V122 237765.3798982527
L41_122 V41 V122 -1.5322959488559718e-11
C41_122 V41 V122 -4.993509086942312e-20

R41_123 V41 V123 -4222.114834330643
L41_123 V41 V123 -2.7998077238988084e-12
C41_123 V41 V123 -9.558845632823926e-20

R41_124 V41 V124 -7770.211800312859
L41_124 V41 V124 -1.965244201530447e-12
C41_124 V41 V124 -2.172927284332017e-19

R41_125 V41 V125 -2200.416766247924
L41_125 V41 V125 6.122401010758334e-12
C41_125 V41 V125 -3.23080191066158e-20

R41_126 V41 V126 11200.420450770953
L41_126 V41 V126 -3.203018660094095e-11
C41_126 V41 V126 -1.3965327238007056e-19

R41_127 V41 V127 3310.5760497669467
L41_127 V41 V127 6.484214573615438e-12
C41_127 V41 V127 -3.7903556787970275e-20

R41_128 V41 V128 2953.802121552923
L41_128 V41 V128 4.107701618850729e-12
C41_128 V41 V128 -3.755257780844568e-21

R41_129 V41 V129 1551.004850526163
L41_129 V41 V129 -1.9752685684450063e-12
C41_129 V41 V129 -2.589633348842419e-19

R41_130 V41 V130 6622.087684754415
L41_130 V41 V130 7.331984828802465e-12
C41_130 V41 V130 1.6044995054181746e-19

R41_131 V41 V131 -4506.310046229898
L41_131 V41 V131 2.10960628953798e-11
C41_131 V41 V131 1.0226692677882183e-19

R41_132 V41 V132 -3606.378052210817
L41_132 V41 V132 9.539009316620794e-12
C41_132 V41 V132 2.0253667895692118e-19

R41_133 V41 V133 2767.423007126694
L41_133 V41 V133 1.9513667571557466e-12
C41_133 V41 V133 3.831226299638749e-19

R41_134 V41 V134 -3756.6096323545967
L41_134 V41 V134 -4.150604785817891e-12
C41_134 V41 V134 -2.7320576925539566e-20

R41_135 V41 V135 -19355.227102806683
L41_135 V41 V135 -4.606676791034663e-12
C41_135 V41 V135 -2.07821623771545e-21

R41_136 V41 V136 -8349.985298281581
L41_136 V41 V136 -2.5738273889416274e-12
C41_136 V41 V136 -9.475038022052973e-20

R41_137 V41 V137 -1882.3625688764625
L41_137 V41 V137 -2.4647109564041653e-11
C41_137 V41 V137 1.249861311193212e-19

R41_138 V41 V138 4234.829037345762
L41_138 V41 V138 1.0354130998771374e-11
C41_138 V41 V138 -5.469729083430853e-20

R41_139 V41 V139 2638.932338214353
L41_139 V41 V139 2.4661712777195317e-12
C41_139 V41 V139 1.1995884642900245e-20

R41_140 V41 V140 5222.665435589003
L41_140 V41 V140 2.043358035299656e-12
C41_140 V41 V140 9.868665601232779e-20

R41_141 V41 V141 -2077.837874586754
L41_141 V41 V141 -1.6916103871994884e-12
C41_141 V41 V141 -3.9030776197316897e-19

R41_142 V41 V142 3807.737649667148
L41_142 V41 V142 3.3694571194720336e-12
C41_142 V41 V142 1.1367747044552038e-20

R41_143 V41 V143 -3125.8120716795
L41_143 V41 V143 -5.752459060132944e-12
C41_143 V41 V143 -1.9201725045469565e-20

R41_144 V41 V144 5192.151280780922
L41_144 V41 V144 -3.389140702169563e-11
C41_144 V41 V144 -7.516086936499883e-20

R41_145 V41 V145 1098.5770517702902
L41_145 V41 V145 2.8535438192632526e-12
C41_145 V41 V145 -5.898448867982098e-20

R41_146 V41 V146 -2511.474074712383
L41_146 V41 V146 -2.7690065346972432e-12
C41_146 V41 V146 5.918864824586979e-20

R41_147 V41 V147 3070.8705652578947
L41_147 V41 V147 -3.922447009609291e-12
C41_147 V41 V147 -1.115499007846857e-19

R41_148 V41 V148 -1523.9907264823028
L41_148 V41 V148 -2.3812496843033702e-12
C41_148 V41 V148 -1.1388510022714987e-19

R41_149 V41 V149 6439.858336160694
L41_149 V41 V149 1.7237161190537851e-12
C41_149 V41 V149 2.5428317336844646e-19

R41_150 V41 V150 -1948.3297575459012
L41_150 V41 V150 -1.2927702775922261e-11
C41_150 V41 V150 -1.7825446438780912e-19

R41_151 V41 V151 -1818.2545817749817
L41_151 V41 V151 1.2507571477289794e-11
C41_151 V41 V151 3.419783962554354e-20

R41_152 V41 V152 3104.1171859903366
L41_152 V41 V152 8.958426510077815e-12
C41_152 V41 V152 4.356776348838884e-20

R41_153 V41 V153 -2093.987115393908
L41_153 V41 V153 -2.9057621583017817e-12
C41_153 V41 V153 6.633863713487532e-20

R41_154 V41 V154 3878.4444416584574
L41_154 V41 V154 7.747755992667725e-12
C41_154 V41 V154 1.0087334581038828e-19

R41_155 V41 V155 779.7147270475269
L41_155 V41 V155 3.151539487108382e-12
C41_155 V41 V155 3.9161212675929907e-20

R41_156 V41 V156 -2325.8871377343526
L41_156 V41 V156 7.487788423602191e-12
C41_156 V41 V156 1.220463559047061e-19

R41_157 V41 V157 -9042.302016425714
L41_157 V41 V157 -1.5836375693393526e-12
C41_157 V41 V157 -1.2206531212556582e-19

R41_158 V41 V158 -9899.372140131027
L41_158 V41 V158 7.967243443871528e-12
C41_158 V41 V158 2.405482185148514e-20

R41_159 V41 V159 -1261.8399522985583
L41_159 V41 V159 -7.67869576626053e-12
C41_159 V41 V159 6.29908677653309e-20

R41_160 V41 V160 3312.7388018846377
L41_160 V41 V160 -2.5693122276071257e-10
C41_160 V41 V160 1.0922577864032886e-20

R41_161 V41 V161 3348.681067107163
L41_161 V41 V161 1.9764779979591994e-12
C41_161 V41 V161 -8.635776735719376e-20

R41_162 V41 V162 8907.468343523811
L41_162 V41 V162 7.852066565312347e-12
C41_162 V41 V162 9.242919444689913e-20

R41_163 V41 V163 -5501.826504839855
L41_163 V41 V163 -1.1842416703903235e-11
C41_163 V41 V163 2.564083305867796e-21

R41_164 V41 V164 -1600.0066610035044
L41_164 V41 V164 -1.081133522293443e-11
C41_164 V41 V164 1.4560229874436092e-20

R41_165 V41 V165 2094.3897561433914
L41_165 V41 V165 3.2691861233590077e-12
C41_165 V41 V165 -2.335083298862865e-21

R41_166 V41 V166 -2468.8310714612007
L41_166 V41 V166 -4.5330353185061884e-11
C41_166 V41 V166 -9.898486848557218e-20

R41_167 V41 V167 -3942.5322837943563
L41_167 V41 V167 6.5170019374974996e-12
C41_167 V41 V167 -6.425934561707822e-20

R41_168 V41 V168 1593.3880029411187
L41_168 V41 V168 3.5615019675377654e-12
C41_168 V41 V168 -1.4714298950470184e-19

R41_169 V41 V169 -1508.3804543469278
L41_169 V41 V169 -1.6499926203233165e-12
C41_169 V41 V169 1.1693512478564799e-20

R41_170 V41 V170 4431.162541462925
L41_170 V41 V170 1.124706642441592e-11
C41_170 V41 V170 1.6189937002442472e-20

R41_171 V41 V171 1471.8658544657947
L41_171 V41 V171 5.898489169052294e-12
C41_171 V41 V171 5.900754887922906e-21

R41_172 V41 V172 5081.400004173371
L41_172 V41 V172 -1.2342203322528033e-11
C41_172 V41 V172 4.458553739825864e-20

R41_173 V41 V173 55148.4553069438
L41_173 V41 V173 3.4946059435380504e-12
C41_173 V41 V173 1.5633827636665094e-19

R41_174 V41 V174 2271.585151296961
L41_174 V41 V174 -6.2949452261538136e-12
C41_174 V41 V174 2.6914835116696638e-20

R41_175 V41 V175 -2262.41210196723
L41_175 V41 V175 -5.305723605020728e-12
C41_175 V41 V175 1.648278788508411e-19

R41_176 V41 V176 -2382.7925169082473
L41_176 V41 V176 -7.076212514878513e-12
C41_176 V41 V176 2.277835108203415e-19

R41_177 V41 V177 3530.7700268779995
L41_177 V41 V177 -1.776079813848156e-11
C41_177 V41 V177 -1.2420790426986615e-19

R41_178 V41 V178 -1566.0110222093683
L41_178 V41 V178 -6.439930240773123e-12
C41_178 V41 V178 -1.8701348157110073e-20

R41_179 V41 V179 5955.263472106104
L41_179 V41 V179 -1.2125801730581301e-11
C41_179 V41 V179 -1.3468905357210386e-19

R41_180 V41 V180 -9107.2937994484
L41_180 V41 V180 -3.968357870214603e-11
C41_180 V41 V180 -1.5835143225285344e-19

R41_181 V41 V181 -9023.804690752237
L41_181 V41 V181 3.848595326767944e-12
C41_181 V41 V181 -1.5570859129316128e-19

R41_182 V41 V182 2207.238591589569
L41_182 V41 V182 2.7301953456568417e-12
C41_182 V41 V182 5.3056980061626125e-20

R41_183 V41 V183 -6435.912365507771
L41_183 V41 V183 -8.482355972946878e-12
C41_183 V41 V183 -5.600947912229407e-20

R41_184 V41 V184 7796.433144710178
L41_184 V41 V184 -9.879062297786155e-12
C41_184 V41 V184 -5.2582254108477806e-20

R41_185 V41 V185 -4837.051514034937
L41_185 V41 V185 -7.78304919684446e-12
C41_185 V41 V185 1.8738015963678177e-19

R41_186 V41 V186 2094.1871575964888
L41_186 V41 V186 -4.024304583833311e-11
C41_186 V41 V186 -1.4240049613365934e-19

R41_187 V41 V187 4677.770904182422
L41_187 V41 V187 4.261330267282109e-12
C41_187 V41 V187 1.0763776415862271e-19

R41_188 V41 V188 1564.6032453852188
L41_188 V41 V188 2.120123076118185e-12
C41_188 V41 V188 7.334235150752751e-20

R41_189 V41 V189 -2006.9016465113955
L41_189 V41 V189 -4.050585444628919e-12
C41_189 V41 V189 8.164793840842127e-20

R41_190 V41 V190 -1788.3725257560936
L41_190 V41 V190 -1.5360967412808784e-11
C41_190 V41 V190 -1.913565999087398e-20

R41_191 V41 V191 -7921.54081875683
L41_191 V41 V191 5.5023223843606505e-12
C41_191 V41 V191 6.394889950735487e-20

R41_192 V41 V192 -2383.023480356191
L41_192 V41 V192 -4.927479801730337e-12
C41_192 V41 V192 7.188180950248912e-20

R41_193 V41 V193 1040.5083601492872
L41_193 V41 V193 2.0774411483791044e-12
C41_193 V41 V193 -1.289630684793197e-20

R41_194 V41 V194 -1923.852253353318
L41_194 V41 V194 -2.5704005186829375e-12
C41_194 V41 V194 3.971522884546229e-21

R41_195 V41 V195 -2841.479293400623
L41_195 V41 V195 -2.3498554702944305e-12
C41_195 V41 V195 -1.5590973030827305e-19

R41_196 V41 V196 -1449.3014670074504
L41_196 V41 V196 -3.3160850668971874e-12
C41_196 V41 V196 -1.774734856139244e-20

R41_197 V41 V197 -10557.383434962967
L41_197 V41 V197 -3.761987577921276e-12
C41_197 V41 V197 -2.0587219885955192e-19

R41_198 V41 V198 2372.4793805922363
L41_198 V41 V198 1.517481715826793e-11
C41_198 V41 V198 -2.0758207162079286e-20

R41_199 V41 V199 2657.3397757097023
L41_199 V41 V199 2.8108295393689292e-11
C41_199 V41 V199 1.7653488574157405e-21

R41_200 V41 V200 915.0973804222872
L41_200 V41 V200 4.7237361012411005e-12
C41_200 V41 V200 -8.626357315190305e-20

R42_42 V42 0 -418.1586574815296
L42_42 V42 0 3.1275862374472126e-12
C42_42 V42 0 7.43021946437999e-20

R42_43 V42 V43 -12546.555644471142
L42_43 V42 V43 -2.1264555140653832e-12
C42_43 V42 V43 -3.235949521889993e-19

R42_44 V42 V44 -10793.408378365877
L42_44 V42 V44 -1.5495312305228336e-12
C42_44 V42 V44 -4.102719609640407e-19

R42_45 V42 V45 7419.546500907195
L42_45 V42 V45 8.12474178259688e-12
C42_45 V42 V45 1.6835416004172526e-20

R42_46 V42 V46 3065.972927965191
L42_46 V42 V46 1.2812224258036068e-12
C42_46 V42 V46 4.423782776912527e-19

R42_47 V42 V47 -6782.732426047699
L42_47 V42 V47 6.943381302700081e-12
C42_47 V42 V47 7.219580889601786e-20

R42_48 V42 V48 -6265.888294423157
L42_48 V42 V48 9.263576101819003e-12
C42_48 V42 V48 4.312891628092017e-20

R42_49 V42 V49 6803.352577571517
L42_49 V42 V49 3.5573377112372334e-12
C42_49 V42 V49 1.911702397660172e-19

R42_50 V42 V50 4205.724564206663
L42_50 V42 V50 8.817137119951373e-13
C42_50 V42 V50 7.327912809542081e-19

R42_51 V42 V51 -29654.710801271725
L42_51 V42 V51 2.5416521606231654e-12
C42_51 V42 V51 2.4760133053924504e-19

R42_52 V42 V52 4526789.492489627
L42_52 V42 V52 2.035721836310433e-12
C42_52 V42 V52 3.663842237480558e-19

R42_53 V42 V53 6436.815144152212
L42_53 V42 V53 -5.1598656459768696e-12
C42_53 V42 V53 -1.415548549718088e-19

R42_54 V42 V54 -12231.49078432914
L42_54 V42 V54 -9.544674157217883e-13
C42_54 V42 V54 -6.120923943666553e-19

R42_55 V42 V55 22772.235971829832
L42_55 V42 V55 -3.4862473518136497e-12
C42_55 V42 V55 -2.0312945272695387e-19

R42_56 V42 V56 12425.99934163203
L42_56 V42 V56 -3.532020084297587e-12
C42_56 V42 V56 -1.487281125989448e-19

R42_57 V42 V57 40602.246036392185
L42_57 V42 V57 -1.2376677289190425e-11
C42_57 V42 V57 -4.4180767497816456e-21

R42_58 V42 V58 -35013.5826342498
L42_58 V42 V58 -2.957138250607473e-11
C42_58 V42 V58 2.910220577348433e-20

R42_59 V42 V59 -72575.11899871788
L42_59 V42 V59 -4.9551519950648776e-12
C42_59 V42 V59 -1.8205779158453144e-19

R42_60 V42 V60 -39882.72654876256
L42_60 V42 V60 -3.7252692466075416e-12
C42_60 V42 V60 -1.9886765985397128e-19

R42_61 V42 V61 -11932.13003779844
L42_61 V42 V61 4.456573960662594e-12
C42_61 V42 V61 9.423808637152777e-20

R42_62 V42 V62 -4627.464975520346
L42_62 V42 V62 3.727522216854374e-12
C42_62 V42 V62 1.6144008570017712e-19

R42_63 V42 V63 -98056.34557602617
L42_63 V42 V63 3.689475274137325e-12
C42_63 V42 V63 2.167927191077248e-19

R42_64 V42 V64 -151254.39319203686
L42_64 V42 V64 2.6578674350369005e-12
C42_64 V42 V64 2.7744959886137587e-19

R42_65 V42 V65 16235.507553054025
L42_65 V42 V65 -3.733226178748972e-11
C42_65 V42 V65 -1.019084684727637e-19

R42_66 V42 V66 6188.096859849575
L42_66 V42 V66 9.595808708541021e-12
C42_66 V42 V66 -5.395661136847823e-20

R42_67 V42 V67 -31483.11291870645
L42_67 V42 V67 1.4869338583380958e-11
C42_67 V42 V67 -3.9283738901074236e-21

R42_68 V42 V68 -22225.421659764153
L42_68 V42 V68 4.018921204310025e-11
C42_68 V42 V68 -4.9781898415597115e-20

R42_69 V42 V69 13657.141888562704
L42_69 V42 V69 -5.211035726854384e-12
C42_69 V42 V69 -7.54001720884701e-20

R42_70 V42 V70 3580.3702978607917
L42_70 V42 V70 -1.0997889948963303e-11
C42_70 V42 V70 -3.1876699057423714e-20

R42_71 V42 V71 -12400.82977338441
L42_71 V42 V71 -1.2108987302793912e-11
C42_71 V42 V71 -6.733148907780822e-20

R42_72 V42 V72 -10254.039202815009
L42_72 V42 V72 -7.09932214303127e-12
C42_72 V42 V72 -9.626283435394139e-20

R42_73 V42 V73 5559.012194407652
L42_73 V42 V73 5.500219952078511e-12
C42_73 V42 V73 1.088757933517545e-19

R42_74 V42 V74 -4628.768543510043
L42_74 V42 V74 -3.979290270179181e-12
C42_74 V42 V74 1.5259335384105317e-21

R42_75 V42 V75 14826.590372292532
L42_75 V42 V75 -1.0285602874358838e-11
C42_75 V42 V75 -4.4578757738500445e-20

R42_76 V42 V76 7653.086682033207
L42_76 V42 V76 7.349202571623889e-11
C42_76 V42 V76 9.933949028091548e-20

R42_77 V42 V77 -28638.556000603894
L42_77 V42 V77 4.429767839535428e-10
C42_77 V42 V77 2.3954948713458167e-20

R42_78 V42 V78 -9743.331865492144
L42_78 V42 V78 1.441109614557904e-12
C42_78 V42 V78 1.8672063907440385e-19

R42_79 V42 V79 22604.92238199121
L42_79 V42 V79 1.0967914915674842e-11
C42_79 V42 V79 2.5491570520724967e-20

R42_80 V42 V80 165951.85088889778
L42_80 V42 V80 8.878676425007207e-12
C42_80 V42 V80 -1.2226385049312661e-20

R42_81 V42 V81 6419.409063237589
L42_81 V42 V81 1.1268974030189214e-11
C42_81 V42 V81 -7.765590483840036e-20

R42_82 V42 V82 4285.625200751893
L42_82 V42 V82 -2.690381385113654e-12
C42_82 V42 V82 -1.6530431865710666e-19

R42_83 V42 V83 -16306.90078186858
L42_83 V42 V83 8.034258974237574e-12
C42_83 V42 V83 6.967335568736913e-20

R42_84 V42 V84 -18429.222814678345
L42_84 V42 V84 1.4362608917883108e-11
C42_84 V42 V84 1.8097571681599475e-20

R42_85 V42 V85 -19986.789491126903
L42_85 V42 V85 -5.777762068651672e-11
C42_85 V42 V85 -1.888060587407039e-20

R42_86 V42 V86 4575.177216371713
L42_86 V42 V86 -1.8188237019368222e-12
C42_86 V42 V86 -1.9950068057393179e-19

R42_87 V42 V87 -5158.212607747956
L42_87 V42 V87 -6.713350698641733e-12
C42_87 V42 V87 -2.3782826842660606e-20

R42_88 V42 V88 -5147.069301126084
L42_88 V42 V88 -8.649181306754878e-12
C42_88 V42 V88 4.735287758561004e-20

R42_89 V42 V89 9850.21845791386
L42_89 V42 V89 -2.6369339026408547e-11
C42_89 V42 V89 9.063032108441172e-22

R42_90 V42 V90 -1855.0942617831327
L42_90 V42 V90 1.0158725257571714e-12
C42_90 V42 V90 4.527651780035803e-19

R42_91 V42 V91 34703.75834794837
L42_91 V42 V91 4.520764448558439e-11
C42_91 V42 V91 -1.3561576051655458e-19

R42_92 V42 V92 9941.11462936393
L42_92 V42 V92 -7.690084053746462e-12
C42_92 V42 V92 -1.706314880371892e-19

R42_93 V42 V93 45303.49897842776
L42_93 V42 V93 5.7310170894800936e-11
C42_93 V42 V93 4.8972712390952943e-20

R42_94 V42 V94 13811.074489608982
L42_94 V42 V94 -4.087715593191226e-12
C42_94 V42 V94 -2.3558953423434967e-19

R42_95 V42 V95 2883.845167319456
L42_95 V42 V95 9.280961511166032e-12
C42_95 V42 V95 5.3983254977913587e-20

R42_96 V42 V96 2562.707302970012
L42_96 V42 V96 5.462704974086888e-12
C42_96 V42 V96 5.158702948106616e-20

R42_97 V42 V97 9135.187159350993
L42_97 V42 V97 -2.500339338085477e-10
C42_97 V42 V97 -4.9542419717735993e-20

R42_98 V42 V98 2841.8286482632107
L42_98 V42 V98 -1.435156830978899e-12
C42_98 V42 V98 -2.812447822671712e-19

R42_99 V42 V99 -1687.3607997594693
L42_99 V42 V99 1.669448948717646e-11
C42_99 V42 V99 1.5106521901566756e-19

R42_100 V42 V100 -1448.038649920828
L42_100 V42 V100 6.572960312136566e-12
C42_100 V42 V100 2.7000366741117686e-19

R42_101 V42 V101 9589.890732913915
L42_101 V42 V101 3.886847678682241e-12
C42_101 V42 V101 6.905549844201056e-21

R42_102 V42 V102 -1686.7223905585608
L42_102 V42 V102 1.2852362719332244e-12
C42_102 V42 V102 5.264889956232893e-19

R42_103 V42 V103 12452.36975426793
L42_103 V42 V103 -2.8098074189087517e-12
C42_103 V42 V103 -2.0102726689059172e-19

R42_104 V42 V104 11999.911572865527
L42_104 V42 V104 -1.8560313687664437e-12
C42_104 V42 V104 -3.200373572670013e-19

R42_105 V42 V105 20487.383559963913
L42_105 V42 V105 -2.766192699124516e-12
C42_105 V42 V105 -4.441266423749475e-20

R42_106 V42 V106 1147.0448197357287
L42_106 V42 V106 -3.655045760911312e-12
C42_106 V42 V106 -1.7300419394907694e-19

R42_107 V42 V107 5229.631695657602
L42_107 V42 V107 3.8692119818836195e-12
C42_107 V42 V107 3.6539015733880034e-20

R42_108 V42 V108 3129.5478544997704
L42_108 V42 V108 3.854422419620549e-12
C42_108 V42 V108 7.409906248407093e-20

R42_109 V42 V109 -3292.817920513317
L42_109 V42 V109 7.175173260075216e-11
C42_109 V42 V109 -3.4275624468723584e-20

R42_110 V42 V110 -2314.272262651847
L42_110 V42 V110 -3.6136072545218434e-12
C42_110 V42 V110 -2.5435011551223455e-19

R42_111 V42 V111 -4813.014921626711
L42_111 V42 V111 4.046690703401891e-12
C42_111 V42 V111 1.1805586450153015e-19

R42_112 V42 V112 -3212.4748938302773
L42_112 V42 V112 4.571790684484549e-12
C42_112 V42 V112 7.197167975948278e-20

R42_113 V42 V113 2738.24092909737
L42_113 V42 V113 1.8022394922164608e-12
C42_113 V42 V113 1.033639429395333e-19

R42_114 V42 V114 -1526.2718549997685
L42_114 V42 V114 3.787720741604569e-12
C42_114 V42 V114 1.6110681852505114e-19

R42_115 V42 V115 23637.27412159503
L42_115 V42 V115 -2.782025082029917e-12
C42_115 V42 V115 -6.585801012876193e-20

R42_116 V42 V116 -46649.10986251635
L42_116 V42 V116 -3.5874722285836917e-12
C42_116 V42 V116 -5.674714850463975e-20

R42_117 V42 V117 2163.529569806223
L42_117 V42 V117 -4.5521972487744834e-12
C42_117 V42 V117 -5.085842247380649e-21

R42_118 V42 V118 983.3063746048352
L42_118 V42 V118 -2.7118306635344432e-12
C42_118 V42 V118 2.467543206818429e-19

R42_119 V42 V119 18448.065953409012
L42_119 V42 V119 -2.1171246938296338e-11
C42_119 V42 V119 2.919310682886331e-20

R42_120 V42 V120 -77632.35117422928
L42_120 V42 V120 1.8331100189045826e-10
C42_120 V42 V120 1.0264503969546316e-19

R42_121 V42 V121 -2365.923063184769
L42_121 V42 V121 -2.3930096993441382e-12
C42_121 V42 V121 -1.1674805574382536e-19

R42_122 V42 V122 -27121.787063715998
L42_122 V42 V122 5.379375931320148e-12
C42_122 V42 V122 -1.4632654412697565e-19

R42_123 V42 V123 32673.462750792904
L42_123 V42 V123 6.865349666754714e-12
C42_123 V42 V123 5.865984173378389e-21

R42_124 V42 V124 9792.32018132719
L42_124 V42 V124 5.979119149340485e-10
C42_124 V42 V124 -1.6646903583927043e-19

R42_125 V42 V125 -3940.03661508545
L42_125 V42 V125 3.449080407828428e-12
C42_125 V42 V125 7.190230347684026e-20

R42_126 V42 V126 -1278.0285753703647
L42_126 V42 V126 5.175444313330975e-12
C42_126 V42 V126 -3.0757227319506437e-19

R42_127 V42 V127 -4506.806166339821
L42_127 V42 V127 5.677500373219997e-12
C42_127 V42 V127 -1.701853336830947e-20

R42_128 V42 V128 -6428.739749766082
L42_128 V42 V128 3.64614009049379e-12
C42_128 V42 V128 4.770498084314486e-20

R42_129 V42 V129 1763.3760504704762
L42_129 V42 V129 3.0514485183763333e-12
C42_129 V42 V129 -3.182407808562954e-20

R42_130 V42 V130 1901.3509064488915
L42_130 V42 V130 -2.3322729559779654e-12
C42_130 V42 V130 2.8395309395504213e-19

R42_131 V42 V131 4021.2261269710416
L42_131 V42 V131 -2.7486691397507315e-12
C42_131 V42 V131 2.4740234975393678e-20

R42_132 V42 V132 3886.968803845196
L42_132 V42 V132 -1.7394080551748153e-12
C42_132 V42 V132 3.9146795270840996e-20

R42_133 V42 V133 6905.136905859499
L42_133 V42 V133 -2.6285105980972096e-12
C42_133 V42 V133 7.723604916201173e-21

R42_134 V42 V134 5017.84086331651
L42_134 V42 V134 3.4810103718107294e-12
C42_134 V42 V134 1.628264289635922e-19

R42_135 V42 V135 11209.253369340278
L42_135 V42 V135 -7.531496393872188e-12
C42_135 V42 V135 -4.238609793014697e-20

R42_136 V42 V136 5487.358927714171
L42_136 V42 V136 -3.3902241930460146e-12
C42_136 V42 V136 -1.7044818558204237e-19

R42_137 V42 V137 -3053.7646898253442
L42_137 V42 V137 -1.5697788990024843e-11
C42_137 V42 V137 9.394971258252781e-21

R42_138 V42 V138 -2690.6793870974598
L42_138 V42 V138 -9.532148020694803e-12
C42_138 V42 V138 -2.950460299849993e-19

R42_139 V42 V139 -3653.220301874372
L42_139 V42 V139 2.187549060061238e-12
C42_139 V42 V139 6.372549541487876e-20

R42_140 V42 V140 -1949.3115436842293
L42_140 V42 V140 1.1621728003459658e-12
C42_140 V42 V140 2.3910293996800975e-19

R42_141 V42 V141 -4105.919039430499
L42_141 V42 V141 1.2152884441937056e-10
C42_141 V42 V141 1.0023376900438944e-20

R42_142 V42 V142 -2331.4572380052696
L42_142 V42 V142 -2.7926246242112786e-12
C42_142 V42 V142 -1.267558875113597e-20

R42_143 V42 V143 6658.308163707282
L42_143 V42 V143 -5.21027455064835e-12
C42_143 V42 V143 2.0932138018651036e-20

R42_144 V42 V144 3414.125048827935
L42_144 V42 V144 -3.126982705911444e-12
C42_144 V42 V144 -4.7246116136000206e-20

R42_145 V42 V145 1153.9589248734262
L42_145 V42 V145 -1.4664661904723429e-10
C42_145 V42 V145 -1.8493694665528026e-20

R42_146 V42 V146 495.46853335582455
L42_146 V42 V146 4.434917379141248e-12
C42_146 V42 V146 1.3493687394725415e-19

R42_147 V42 V147 2384.2506087407214
L42_147 V42 V147 -3.904819430707413e-12
C42_147 V42 V147 -1.3284022426259695e-19

R42_148 V42 V148 3946.004704101489
L42_148 V42 V148 -3.6551047236022465e-12
C42_148 V42 V148 -1.5040319912344377e-19

R42_149 V42 V149 -4209.2914568724555
L42_149 V42 V149 3.2616886437562513e-12
C42_149 V42 V149 -7.406262790583028e-20

R42_150 V42 V150 -716.9041413836909
L42_150 V42 V150 3.6133639004840962e-12
C42_150 V42 V150 4.807821674501221e-20

R42_151 V42 V151 -1415.4720502392945
L42_151 V42 V151 3.7488374598157155e-11
C42_151 V42 V151 5.380777425551359e-21

R42_152 V42 V152 -1197.407799471843
L42_152 V42 V152 5.5128208724153704e-12
C42_152 V42 V152 4.953252032017225e-20

R42_153 V42 V153 -3186.029998077799
L42_153 V42 V153 -9.08545863296274e-12
C42_153 V42 V153 2.415311703425638e-20

R42_154 V42 V154 -1151.6826490484507
L42_154 V42 V154 -3.573081323566144e-12
C42_154 V42 V154 -1.2322256493773098e-19

R42_155 V42 V155 1333.212338443267
L42_155 V42 V155 8.976394348712266e-12
C42_155 V42 V155 1.8691836289292725e-20

R42_156 V42 V156 1512.1008313119635
L42_156 V42 V156 9.691993447166787e-12
C42_156 V42 V156 1.011160326751876e-19

R42_157 V42 V157 -3541.783727716478
L42_157 V42 V157 -2.6932912171372957e-12
C42_157 V42 V157 6.467834036688516e-20

R42_158 V42 V158 875.4619589190781
L42_158 V42 V158 -3.7119144986053325e-12
C42_158 V42 V158 3.3551695951906355e-20

R42_159 V42 V159 4782.32664911085
L42_159 V42 V159 -2.413845809725462e-11
C42_159 V42 V159 3.8673110432830616e-21

R42_160 V42 V160 2081.435508510103
L42_160 V42 V160 -6.5092301355232086e-12
C42_160 V42 V160 -5.03161922438122e-20

R42_161 V42 V161 7014.751191863591
L42_161 V42 V161 2.045750657364536e-12
C42_161 V42 V161 2.982241897216397e-20

R42_162 V42 V162 1034.7715499306237
L42_162 V42 V162 1.5212318155701778e-12
C42_162 V42 V162 7.042264200491369e-20

R42_163 V42 V163 -1690.0263642798561
L42_163 V42 V163 5.022875044666344e-12
C42_163 V42 V163 3.709517151550249e-20

R42_164 V42 V164 -1159.6791411112997
L42_164 V42 V164 4.997944020564434e-12
C42_164 V42 V164 3.083997929241734e-20

R42_165 V42 V165 1246.593433304078
L42_165 V42 V165 5.558969843574121e-12
C42_165 V42 V165 -1.3292878471178882e-19

R42_166 V42 V166 -565.0932471542465
L42_166 V42 V166 9.277510153943312e-12
C42_166 V42 V166 -9.205072836282996e-20

R42_167 V42 V167 2904.75059598422
L42_167 V42 V167 6.126153340681095e-12
C42_167 V42 V167 2.4077652477481096e-20

R42_168 V42 V168 1204.7395242151022
L42_168 V42 V168 3.2872676952711965e-12
C42_168 V42 V168 1.7759044106836622e-20

R42_169 V42 V169 -3342.3621010301804
L42_169 V42 V169 -1.3844731374560654e-12
C42_169 V42 V169 -7.318644878522927e-20

R42_170 V42 V170 3303.9268014622735
L42_170 V42 V170 -1.0614982749471122e-12
C42_170 V42 V170 -1.2297094006656473e-20

R42_171 V42 V171 2177.077383114038
L42_171 V42 V171 -2.9434188907004104e-12
C42_171 V42 V171 -1.2350493882768859e-19

R42_172 V42 V172 4608.014697463012
L42_172 V42 V172 -2.764593838628888e-12
C42_172 V42 V172 -7.818219700729683e-20

R42_173 V42 V173 -702267.7620350973
L42_173 V42 V173 2.562815836163598e-12
C42_173 V42 V173 1.85737669837447e-19

R42_174 V42 V174 778.50617228066
L42_174 V42 V174 3.3315144906194225e-12
C42_174 V42 V174 6.66730592908202e-20

R42_175 V42 V175 -1471.849952738814
L42_175 V42 V175 -7.1823777335173526e-12
C42_175 V42 V175 5.553841648269621e-20

R42_176 V42 V176 -1266.3336800058398
L42_176 V42 V176 -1.0707985438552702e-11
C42_176 V42 V176 1.0747780885737763e-19

R42_177 V42 V177 2601.931047859811
L42_177 V42 V177 2.8827868697573663e-12
C42_177 V42 V177 -7.049188338860034e-20

R42_178 V42 V178 -1601.6077315575665
L42_178 V42 V178 1.1144415709236967e-12
C42_178 V42 V178 -1.291686355702734e-21

R42_179 V42 V179 2823.7366155100735
L42_179 V42 V179 2.93235342757934e-12
C42_179 V42 V179 4.190993430504587e-20

R42_180 V42 V180 1924.723574063255
L42_180 V42 V180 2.927965824277233e-12
C42_180 V42 V180 -1.7537247793876637e-21

R42_181 V42 V181 -3618.9678883170645
L42_181 V42 V181 -3.5646694982342292e-12
C42_181 V42 V181 -7.662519927944586e-20

R42_182 V42 V182 -2752.624200622729
L42_182 V42 V182 -1.194226704282893e-12
C42_182 V42 V182 -4.571572616418486e-20

R42_183 V42 V183 6513.4572078460205
L42_183 V42 V183 1.0559163589572558e-11
C42_183 V42 V183 -1.6063353387062772e-20

R42_184 V42 V184 6094.021492210787
L42_184 V42 V184 1.873567724379288e-11
C42_184 V42 V184 -2.2497805433826503e-20

R42_185 V42 V185 -9863.17525541836
L42_185 V42 V185 -5.2228252883801246e-12
C42_185 V42 V185 9.047518236580481e-20

R42_186 V42 V186 5596.14580395849
L42_186 V42 V186 -1.6799466338190382e-12
C42_186 V42 V186 -3.446598347120189e-20

R42_187 V42 V187 -7482.135703841635
L42_187 V42 V187 -6.424768180907893e-12
C42_187 V42 V187 -5.071903858817664e-21

R42_188 V42 V188 -3680.892817881689
L42_188 V42 V188 -2.418739874958256e-11
C42_188 V42 V188 2.0847033893661465e-21

R42_189 V42 V189 35661.937867361405
L42_189 V42 V189 3.5700109582375894e-12
C42_189 V42 V189 -3.0446198240343994e-20

R42_190 V42 V190 2637.5570770821178
L42_190 V42 V190 1.0271634606035772e-12
C42_190 V42 V190 6.002307737032103e-20

R42_191 V42 V191 -9260.145624651166
L42_191 V42 V191 1.0326062445195262e-11
C42_191 V42 V191 -3.7601498972990477e-20

R42_192 V42 V192 62206.23340009716
L42_192 V42 V192 -2.894090783448696e-11
C42_192 V42 V192 -7.759613943509681e-20

R42_193 V42 V193 4435.545326922692
L42_193 V42 V193 3.29411556976704e-12
C42_193 V42 V193 1.1708344165789016e-20

R42_194 V42 V194 -2723.0780085455335
L42_194 V42 V194 -1.303083024703384e-12
C42_194 V42 V194 -1.0790445966740637e-19

R42_195 V42 V195 40482.457307701894
L42_195 V42 V195 1.2934384532343528e-11
C42_195 V42 V195 3.411753545363159e-20

R42_196 V42 V196 -7745.563695404423
L42_196 V42 V196 3.221978266239663e-12
C42_196 V42 V196 2.1033020308721413e-19

R42_197 V42 V197 -4679.280518821479
L42_197 V42 V197 -3.3848418964122283e-12
C42_197 V42 V197 2.3825798280866837e-21

R42_198 V42 V198 -1491.5471836224742
L42_198 V42 V198 -1.9735812147868075e-12
C42_198 V42 V198 2.8673843767666347e-21

R42_199 V42 V199 -82930.24069647696
L42_199 V42 V199 2.497064551473706e-11
C42_199 V42 V199 5.276882320560906e-20

R42_200 V42 V200 2758.219151301906
L42_200 V42 V200 3.637066177531221e-11
C42_200 V42 V200 -8.55915728242537e-21

R43_43 V43 0 -1356.77596584338
L43_43 V43 0 -9.005723734824024e-13
C43_43 V43 0 -3.5185440760562357e-19

R43_44 V43 V44 -6692.56673419647
L43_44 V43 V44 -1.4824310285516574e-12
C43_44 V43 V44 -4.630064725211972e-19

R43_45 V43 V45 5519.685140703304
L43_45 V43 V45 2.6230077985298097e-12
C43_45 V43 V45 1.4823021065420134e-19

R43_46 V43 V46 -319641.5975398505
L43_46 V43 V46 2.8097226140175535e-12
C43_46 V43 V46 2.1296287221668843e-19

R43_47 V43 V47 7766.424836168184
L43_47 V43 V47 7.485274196409033e-13
C43_47 V43 V47 8.025164502257319e-19

R43_48 V43 V48 -4072.4116454352315
L43_48 V43 V48 2.473939001972186e-12
C43_48 V43 V48 2.044025053429609e-19

R43_49 V43 V49 4112.5263809707085
L43_49 V43 V49 3.8149829650194924e-12
C43_49 V43 V49 1.85787003300764e-19

R43_50 V43 V50 25956.995347936772
L43_50 V43 V50 2.1409842906697554e-12
C43_50 V43 V50 3.1349359538015613e-19

R43_51 V43 V51 11660.666409487227
L43_51 V43 V51 2.372390486939469e-12
C43_51 V43 V51 1.9751456546285915e-19

R43_52 V43 V52 -206293.9451667294
L43_52 V43 V52 3.5196741489232973e-12
C43_52 V43 V52 1.67246347911215e-19

R43_53 V43 V53 5476.351807847627
L43_53 V43 V53 -3.830614273057572e-12
C43_53 V43 V53 -2.207883147279883e-19

R43_54 V43 V54 15533.297437702488
L43_54 V43 V54 -2.0433893800309915e-12
C43_54 V43 V54 -3.0679463485943503e-19

R43_55 V43 V55 10234.81421563918
L43_55 V43 V55 -9.793995457345079e-13
C43_55 V43 V55 -6.182140318556519e-19

R43_56 V43 V56 4913.470449504121
L43_56 V43 V56 -2.091046778730559e-12
C43_56 V43 V56 -2.767106197538883e-19

R43_57 V43 V57 29446.449932626227
L43_57 V43 V57 -7.803983375923482e-12
C43_57 V43 V57 5.1352828776597355e-20

R43_58 V43 V58 -8444.146849775561
L43_58 V43 V58 -1.241348225655528e-11
C43_58 V43 V58 -4.662788492129967e-20

R43_59 V43 V59 -5337.574488847762
L43_59 V43 V59 8.645475169959762e-12
C43_59 V43 V59 2.298280455863367e-19

R43_60 V43 V60 -22636.060032766243
L43_60 V43 V60 -7.752471213256392e-12
C43_60 V43 V60 4.135266845281296e-20

R43_61 V43 V61 -8550.511957942204
L43_61 V43 V61 3.7123365099813816e-12
C43_61 V43 V61 9.971973024620232e-20

R43_62 V43 V62 53214.97563165744
L43_62 V43 V62 3.4091066976074737e-12
C43_62 V43 V62 2.2622886177649024e-19

R43_63 V43 V63 -13441.85377932182
L43_63 V43 V63 6.304701998934266e-12
C43_63 V43 V63 4.896569816386448e-20

R43_64 V43 V64 -18968.11369090046
L43_64 V43 V64 3.5848281358659915e-12
C43_64 V43 V64 1.5329857647509713e-19

R43_65 V43 V65 10130.455953463575
L43_65 V43 V65 8.082792632453553e-12
C43_65 V43 V65 8.091785072911364e-21

R43_66 V43 V66 25852.622354018036
L43_66 V43 V66 4.572374308958596e-11
C43_66 V43 V66 -1.5581389068363752e-20

R43_67 V43 V67 10137.983201283867
L43_67 V43 V67 6.889394761759011e-12
C43_67 V43 V67 -3.440151089534742e-20

R43_68 V43 V68 -16213.77676392873
L43_68 V43 V68 1.1079973110130917e-11
C43_68 V43 V68 -7.052420954949493e-20

R43_69 V43 V69 5252.875878306673
L43_69 V43 V69 -4.601964072390665e-12
C43_69 V43 V69 -1.3232659020708826e-19

R43_70 V43 V70 -21885.01655588636
L43_70 V43 V70 -7.983044103297603e-12
C43_70 V43 V70 -8.431416247604257e-20

R43_71 V43 V71 23186.80307595427
L43_71 V43 V71 -3.9294508043122226e-10
C43_71 V43 V71 4.3246392271956027e-20

R43_72 V43 V72 -7282.682352675668
L43_72 V43 V72 2.1075941346037507e-10
C43_72 V43 V72 1.8156736466335175e-20

R43_73 V43 V73 11155.812806137486
L43_73 V43 V73 2.069934705382896e-11
C43_73 V43 V73 3.204205994656084e-20

R43_74 V43 V74 355095.1068013637
L43_74 V43 V74 -2.948102173248493e-11
C43_74 V43 V74 2.2889303445892915e-20

R43_75 V43 V75 -5620.446585962334
L43_75 V43 V75 -2.5198514960586904e-12
C43_75 V43 V75 -1.2143258792581725e-19

R43_76 V43 V76 5653.803147573389
L43_76 V43 V76 -3.701292446000419e-12
C43_76 V43 V76 -6.159355822532346e-20

R43_77 V43 V77 -15625.268502652494
L43_77 V43 V77 1.271269709351327e-10
C43_77 V43 V77 1.2275017265315848e-19

R43_78 V43 V78 -74961.80323807437
L43_78 V43 V78 1.4454301339746205e-11
C43_78 V43 V78 -3.999029420813208e-20

R43_79 V43 V79 9462.309978609548
L43_79 V43 V79 2.298045757733023e-12
C43_79 V43 V79 1.313019172792545e-19

R43_80 V43 V80 13227.51309377958
L43_80 V43 V80 8.208693452890106e-12
C43_80 V43 V80 1.5534284338237253e-20

R43_81 V43 V81 4452.772772449219
L43_81 V43 V81 4.502760697748805e-12
C43_81 V43 V81 -2.612751621645657e-20

R43_82 V43 V82 68235.98456826489
L43_82 V43 V82 1.0104921915225685e-11
C43_82 V43 V82 1.023866227439191e-19

R43_83 V43 V83 -129414.52065589145
L43_83 V43 V83 -4.4775695048803755e-11
C43_83 V43 V83 -9.894553670930591e-21

R43_84 V43 V84 -6943.084724676268
L43_84 V43 V84 3.763750131450559e-12
C43_84 V43 V84 1.3404872717864893e-19

R43_85 V43 V85 88069.76704333913
L43_85 V43 V85 1.7381942458960054e-10
C43_85 V43 V85 -3.14022843526329e-20

R43_86 V43 V86 -8357.875960515925
L43_86 V43 V86 -3.52317038668694e-11
C43_86 V43 V86 2.7008115018661374e-20

R43_87 V43 V87 -3264.378965843892
L43_87 V43 V87 -1.3437021171694483e-12
C43_87 V43 V87 -3.1198082374998378e-19

R43_88 V43 V88 -2813.8063090235373
L43_88 V43 V88 -3.1276679327574453e-12
C43_88 V43 V88 -1.3587030879803886e-19

R43_89 V43 V89 8386.129803656573
L43_89 V43 V89 -8.180347166821535e-12
C43_89 V43 V89 -8.823758930274935e-20

R43_90 V43 V90 -29914.655419615592
L43_90 V43 V90 -3.806891842513121e-12
C43_90 V43 V90 -2.1089232495294662e-19

R43_91 V43 V91 3616.0626847505177
L43_91 V43 V91 6.16202908419481e-13
C43_91 V43 V91 6.208308635255717e-19

R43_92 V43 V92 2976.0005242209863
L43_92 V43 V92 6.3507499884984625e-12
C43_92 V43 V92 -2.689237961000421e-20

R43_93 V43 V93 -32950.01978587771
L43_93 V43 V93 -9.00793499510866e-12
C43_93 V43 V93 -1.674640125203716e-21

R43_94 V43 V94 7311.016045801259
L43_94 V43 V94 -1.2549848629726022e-10
C43_94 V43 V94 4.0419121741827255e-20

R43_95 V43 V95 4580.526032104887
L43_95 V43 V95 -8.90838871999259e-12
C43_95 V43 V95 -6.136113200176988e-20

R43_96 V43 V96 2020.113415238941
L43_96 V43 V96 6.441060638609746e-12
C43_96 V43 V96 1.3092393868780475e-19

R43_97 V43 V97 2910.9460339577704
L43_97 V43 V97 3.0062631104530615e-12
C43_97 V43 V97 2.7769835076122317e-19

R43_98 V43 V98 -10857.789136975507
L43_98 V43 V98 2.8116211057941873e-12
C43_98 V43 V98 2.045691668433317e-19

R43_99 V43 V99 -2459.55745896477
L43_99 V43 V99 -5.661461908270716e-13
C43_99 V43 V99 -6.762402421794324e-19

R43_100 V43 V100 -1078.4176090692592
L43_100 V43 V100 -4.3450142532025605e-12
C43_100 V43 V100 1.4177977131920368e-20

R43_101 V43 V101 12074.820322374084
L43_101 V43 V101 6.392914237684127e-12
C43_101 V43 V101 -1.1186222774230621e-19

R43_102 V43 V102 -8186.88785373024
L43_102 V43 V102 -6.4075671223976065e-12
C43_102 V43 V102 -8.106984976678707e-20

R43_103 V43 V103 -3959.61336566824
L43_103 V43 V103 7.742992888164973e-13
C43_103 V43 V103 6.516073905267714e-19

R43_104 V43 V104 -367266.9285660041
L43_104 V43 V104 -1.587167706358659e-11
C43_104 V43 V104 -1.1106389494831046e-19

R43_105 V43 V105 -15099.104212926695
L43_105 V43 V105 -2.3099782931671897e-12
C43_105 V43 V105 -1.8286439010255355e-19

R43_106 V43 V106 -5875.664786263233
L43_106 V43 V106 -1.6438968328680938e-12
C43_106 V43 V106 -2.849300608833682e-19

R43_107 V43 V107 2612.4316995900276
L43_107 V43 V107 2.881374354175642e-12
C43_107 V43 V107 -8.229685150540614e-20

R43_108 V43 V108 2003.957282801151
L43_108 V43 V108 5.726705561011203e-12
C43_108 V43 V108 4.006418361089171e-20

R43_109 V43 V109 -18779.88619031002
L43_109 V43 V109 1.2431960009593868e-11
C43_109 V43 V109 1.5198651530492484e-19

R43_110 V43 V110 3543.098168556476
L43_110 V43 V110 2.508979047351018e-12
C43_110 V43 V110 1.6544724271620467e-19

R43_111 V43 V111 12072.206757193244
L43_111 V43 V111 -1.5325950814883711e-12
C43_111 V43 V111 -2.026158012632013e-19

R43_112 V43 V112 -2652.4448572050314
L43_112 V43 V112 -7.741063567766324e-11
C43_112 V43 V112 2.5538892644999585e-20

R43_113 V43 V113 1946.3669230512708
L43_113 V43 V113 1.7157218879407638e-12
C43_113 V43 V113 1.2512916453647778e-19

R43_114 V43 V114 14766.364134282487
L43_114 V43 V114 2.1777717629157674e-12
C43_114 V43 V114 2.307327557417589e-19

R43_115 V43 V115 -3474.865206882227
L43_115 V43 V115 -1.838934024415722e-12
C43_115 V43 V115 6.579740342948068e-20

R43_116 V43 V116 -81223.54233968443
L43_116 V43 V116 -5.1455042263092216e-12
C43_116 V43 V116 8.328801606524611e-21

R43_117 V43 V117 2737.787293115912
L43_117 V43 V117 -3.5254738081726972e-12
C43_117 V43 V117 -1.0075028728195168e-19

R43_118 V43 V118 -2635.4339419650496
L43_118 V43 V118 -1.4375994612835503e-12
C43_118 V43 V118 -2.693708733180296e-19

R43_119 V43 V119 4407.142691091924
L43_119 V43 V119 1.7285177764314741e-12
C43_119 V43 V119 -4.0313302198566645e-20

R43_120 V43 V120 -6956.254750305691
L43_120 V43 V120 2.67237483840281e-10
C43_120 V43 V120 -9.60235301184497e-20

R43_121 V43 V121 -2028.2916528402536
L43_121 V43 V121 -3.642891430831424e-12
C43_121 V43 V121 -9.367801175556144e-21

R43_122 V43 V122 11030.419325325483
L43_122 V43 V122 4.4767117583667083e-10
C43_122 V43 V122 -5.136164051656417e-21

R43_123 V43 V123 -12928.575760880898
L43_123 V43 V123 3.074699666530917e-12
C43_123 V43 V123 2.8474908922471215e-19

R43_124 V43 V124 16051.932657053112
L43_124 V43 V124 8.526422809208061e-12
C43_124 V43 V124 5.775582212588151e-20

R43_125 V43 V125 -3408.1918698254185
L43_125 V43 V125 3.5713211067292573e-12
C43_125 V43 V125 6.855790181860247e-23

R43_126 V43 V126 5514.809839644256
L43_126 V43 V126 1.2922705337863002e-12
C43_126 V43 V126 1.6023331284742427e-19

R43_127 V43 V127 64749.93897162774
L43_127 V43 V127 -1.4352765506532584e-12
C43_127 V43 V127 -3.2004228929677903e-19

R43_128 V43 V128 3490.1480720909735
L43_128 V43 V128 5.656460061283256e-12
C43_128 V43 V128 1.4006381730067205e-19

R43_129 V43 V129 1131.7375534637918
L43_129 V43 V129 4.908173274419618e-12
C43_129 V43 V129 4.823157742226743e-20

R43_130 V43 V130 -40378.64401612825
L43_130 V43 V130 -2.5133669830003605e-12
C43_130 V43 V130 -4.660484340172522e-20

R43_131 V43 V131 95672.20796990328
L43_131 V43 V131 6.329839353563973e-12
C43_131 V43 V131 6.468128314128705e-20

R43_132 V43 V132 -2666.5867667384837
L43_132 V43 V132 -2.0886455023615645e-12
C43_132 V43 V132 -2.9501377088868302e-19

R43_133 V43 V133 4948.876454795201
L43_133 V43 V133 -7.614694724002459e-12
C43_133 V43 V133 2.4932119955594868e-20

R43_134 V43 V134 -3636.8223913516745
L43_134 V43 V134 -8.899943526335264e-12
C43_134 V43 V134 -4.740080384852947e-20

R43_135 V43 V135 -2282.1055776054827
L43_135 V43 V135 2.4128477139319773e-12
C43_135 V43 V135 5.739169987039482e-19

R43_136 V43 V136 -4277.742166520935
L43_136 V43 V136 -8.786449382957402e-12
C43_136 V43 V136 1.3945886675335613e-21

R43_137 V43 V137 -1074.1330900876794
L43_137 V43 V137 -5.81394008515329e-12
C43_137 V43 V137 -3.577666536275696e-20

R43_138 V43 V138 4434.777752775744
L43_138 V43 V138 2.443867098498932e-12
C43_138 V43 V138 1.087226588069015e-19

R43_139 V43 V139 2168.041712228383
L43_139 V43 V139 -1.6603428496065997e-12
C43_139 V43 V139 -8.383259262370295e-19

R43_140 V43 V140 3455.602341291655
L43_140 V43 V140 1.98000000714722e-12
C43_140 V43 V140 1.0480137096462384e-19

R43_141 V43 V141 -4135.792133786596
L43_141 V43 V141 4.0971413739072704e-11
C43_141 V43 V141 8.507188234484555e-20

R43_142 V43 V142 3545.959336421478
L43_142 V43 V142 -2.7007086864846676e-11
C43_142 V43 V142 1.4637565165138932e-20

R43_143 V43 V143 1504.8059071911528
L43_143 V43 V143 1.0839512123572553e-11
C43_143 V43 V143 1.7174137297719782e-19

R43_144 V43 V144 1843.8168370201615
L43_144 V43 V144 -6.462261908040573e-12
C43_144 V43 V144 -5.932811310227454e-20

R43_145 V43 V145 656.016242788166
L43_145 V43 V145 3.07545222451496e-12
C43_145 V43 V145 6.700932578569458e-20

R43_146 V43 V146 4101.86417564026
L43_146 V43 V146 -2.895493448529318e-12
C43_146 V43 V146 -7.511704865924809e-20

R43_147 V43 V147 -1347.5492901001035
L43_147 V43 V147 3.846022957144603e-12
C43_147 V43 V147 5.219239802943622e-19

R43_148 V43 V148 -1265.4682089072953
L43_148 V43 V148 -7.161832122156188e-12
C43_148 V43 V148 9.683347334841348e-21

R43_149 V43 V149 -2180.51467116932
L43_149 V43 V149 -6.673202748293101e-12
C43_149 V43 V149 -2.6826669246919834e-19

R43_150 V43 V150 -1063.246466014525
L43_150 V43 V150 5.5611797047096495e-12
C43_150 V43 V150 9.176718476671404e-21

R43_151 V43 V151 -1290.272196701002
L43_151 V43 V151 -9.04247000807417e-11
C43_151 V43 V151 -2.6655157195601645e-19

R43_152 V43 V152 5394.411545950182
L43_152 V43 V152 9.917980037287284e-12
C43_152 V43 V152 3.578154117488414e-20

R43_153 V43 V153 -1589.5318979759097
L43_153 V43 V153 -9.627582745849649e-12
C43_153 V43 V153 7.314050601813956e-20

R43_154 V43 V154 -47586.61463052955
L43_154 V43 V154 6.106427303238262e-11
C43_154 V43 V154 3.443277116150899e-20

R43_155 V43 V155 4169.561424065474
L43_155 V43 V155 -1.3251857145676238e-12
C43_155 V43 V155 -3.144663810843479e-19

R43_156 V43 V156 -4545.357576533881
L43_156 V43 V156 8.183485301480351e-12
C43_156 V43 V156 2.6154567698310754e-20

R43_157 V43 V157 -5414.649664533919
L43_157 V43 V157 -8.694235688136603e-12
C43_157 V43 V157 1.7972273791495124e-19

R43_158 V43 V158 27903.843950302602
L43_158 V43 V158 -2.138189722182639e-11
C43_158 V43 V158 -4.3880687238913923e-20

R43_159 V43 V159 876.4532303506775
L43_159 V43 V159 2.0386742974005715e-12
C43_159 V43 V159 3.682619188915814e-19

R43_160 V43 V160 3682.4307933195805
L43_160 V43 V160 -4.751202623001603e-12
C43_160 V43 V160 -4.3629061639299573e-20

R43_161 V43 V161 2330.6476461705365
L43_161 V43 V161 4.754414961996889e-12
C43_161 V43 V161 -1.3242279205481988e-19

R43_162 V43 V162 3126.1079969847688
L43_162 V43 V162 -9.983097962603123e-12
C43_162 V43 V162 -7.815893664997985e-20

R43_163 V43 V163 -1895.5517986616308
L43_163 V43 V163 1.7575678607030167e-12
C43_163 V43 V163 -1.4132555806575037e-19

R43_164 V43 V164 -1366.2117574994716
L43_164 V43 V164 4.64968470389656e-12
C43_164 V43 V164 -4.4167427508979274e-20

R43_165 V43 V165 2183.182285750821
L43_165 V43 V165 1.9531827260875607e-12
C43_165 V43 V165 2.9025388064987656e-20

R43_166 V43 V166 -1760.890908939164
L43_166 V43 V166 4.3853668271483986e-12
C43_166 V43 V166 4.569260013805887e-20

R43_167 V43 V167 -931.1238182288087
L43_167 V43 V167 -1.7239932968089443e-12
C43_167 V43 V167 -1.0353440770459367e-19

R43_168 V43 V168 1058.6924745082251
L43_168 V43 V168 6.550107860505556e-12
C43_168 V43 V168 -2.8243099018326787e-20

R43_169 V43 V169 -2887.5635131524655
L43_169 V43 V169 -4.1020253122111e-12
C43_169 V43 V169 1.2825772087054428e-19

R43_170 V43 V170 3340.1400026847355
L43_170 V43 V170 -1.455200602426786e-11
C43_170 V43 V170 -3.236130913483061e-20

R43_171 V43 V171 1250.8522470455696
L43_171 V43 V171 -2.775744807253204e-12
C43_171 V43 V171 1.0429148683568451e-19

R43_172 V43 V172 7595.211857957266
L43_172 V43 V172 -1.086596350971618e-11
C43_172 V43 V172 3.2150942886360505e-20

R43_173 V43 V173 117600.46494986978
L43_173 V43 V173 -3.2786915319778256e-12
C43_173 V43 V173 -4.3647567127757663e-20

R43_174 V43 V174 5776.3340463343075
L43_174 V43 V174 -2.9937137923590467e-12
C43_174 V43 V174 5.28304357165433e-20

R43_175 V43 V175 7937.1530905202735
L43_175 V43 V175 4.786184282296869e-12
C43_175 V43 V175 -2.0617101450112317e-19

R43_176 V43 V176 -1417.512145941934
L43_176 V43 V176 -5.7400190295084064e-12
C43_176 V43 V176 5.441950331815554e-20

R43_177 V43 V177 5537.317944014191
L43_177 V43 V177 2.343156125865527e-12
C43_177 V43 V177 -2.5415961762062762e-20

R43_178 V43 V178 -3543.752324357353
L43_178 V43 V178 4.153899309617772e-12
C43_178 V43 V178 2.0346102287372015e-20

R43_179 V43 V179 -1965.11505397037
L43_179 V43 V179 1.7317822582767387e-12
C43_179 V43 V179 1.8024503746400332e-19

R43_180 V43 V180 3593.0664109220943
L43_180 V43 V180 5.864841292715555e-12
C43_180 V43 V180 2.363636018506739e-20

R43_181 V43 V181 -3057.693981489035
L43_181 V43 V181 -8.775936307380455e-12
C43_181 V43 V181 -1.9644641187236997e-20

R43_182 V43 V182 17646.775650928306
L43_182 V43 V182 -1.3948030585407015e-11
C43_182 V43 V182 -5.301782347197695e-20

R43_183 V43 V183 3097.7824150671036
L43_183 V43 V183 -3.74281189962864e-12
C43_183 V43 V183 -6.909987096483465e-21

R43_184 V43 V184 7201.499075583103
L43_184 V43 V184 4.322347165272986e-12
C43_184 V43 V184 1.6148159295268377e-20

R43_185 V43 V185 6060.587836264302
L43_185 V43 V185 -3.8323565488766205e-12
C43_185 V43 V185 1.840663276523288e-20

R43_186 V43 V186 5477.2115423508385
L43_186 V43 V186 -9.534530748473776e-11
C43_186 V43 V186 1.3348447458131388e-20

R43_187 V43 V187 34317.27468345332
L43_187 V43 V187 -2.529848148173852e-12
C43_187 V43 V187 -2.1229107817123042e-19

R43_188 V43 V188 4096.854835303255
L43_188 V43 V188 -3.782532880505152e-12
C43_188 V43 V188 -9.255054647634453e-20

R43_189 V43 V189 -5619.335841950491
L43_189 V43 V189 4.462834947346301e-12
C43_189 V43 V189 5.583274497431491e-20

R43_190 V43 V190 -4717.090405364888
L43_190 V43 V190 9.108733246098336e-12
C43_190 V43 V190 2.41857304110759e-20

R43_191 V43 V191 -8318.05950606018
L43_191 V43 V191 2.2421692128755714e-12
C43_191 V43 V191 2.0660340895807787e-19

R43_192 V43 V192 -5170.712725534283
L43_192 V43 V192 -9.22827194786746e-12
C43_192 V43 V192 3.611822970984222e-20

R43_193 V43 V193 3920.6726035979027
L43_193 V43 V193 4.680398725330487e-12
C43_193 V43 V193 1.7388323555996334e-20

R43_194 V43 V194 -2758.7849660398297
L43_194 V43 V194 -8.367354161832919e-12
C43_194 V43 V194 9.827398392167887e-20

R43_195 V43 V195 15138.242869774436
L43_195 V43 V195 -1.8463823936608168e-12
C43_195 V43 V195 -3.17078805650112e-19

R43_196 V43 V196 -4731.052632418326
L43_196 V43 V196 2.5259260098932332e-12
C43_196 V43 V196 1.7165270807465794e-19

R43_197 V43 V197 29700.789751355307
L43_197 V43 V197 -3.3672908296624915e-12
C43_197 V43 V197 -9.667460656832891e-20

R43_198 V43 V198 -87132.47935668871
L43_198 V43 V198 -7.942327558956502e-12
C43_198 V43 V198 -2.451858339676639e-20

R43_199 V43 V199 -2176.7283197064485
L43_199 V43 V199 -1.294580231478663e-11
C43_199 V43 V199 -1.32481813524047e-20

R43_200 V43 V200 1604.9742468455145
L43_200 V43 V200 -5.687992063794221e-12
C43_200 V43 V200 -1.5006879203215507e-19

R44_44 V44 0 -819.3280935649326
L44_44 V44 0 -4.99355911627445e-13
C44_44 V44 0 -1.297555188460528e-18

R44_45 V44 V45 4593.815766470957
L44_45 V44 V45 2.433247260027604e-12
C44_45 V44 V45 1.784389822311065e-19

R44_46 V44 V46 -32867.881002558664
L44_46 V44 V46 2.799411034388561e-12
C44_46 V44 V46 2.7082732782954256e-19

R44_47 V44 V47 -5712.173211755277
L44_47 V44 V47 1.6615295054656817e-12
C44_47 V44 V47 3.865332883005655e-19

R44_48 V44 V48 139170.72276120822
L44_48 V44 V48 6.191320687608832e-13
C44_48 V44 V48 1.0137178934299476e-18

R44_49 V44 V49 3346.490150474791
L44_49 V44 V49 2.39045032650009e-12
C44_49 V44 V49 2.9592462124426344e-19

R44_50 V44 V50 65876.13041773492
L44_50 V44 V50 1.3948913348323584e-12
C44_50 V44 V50 4.610175678886773e-19

R44_51 V44 V51 -98077.42938939757
L44_51 V44 V51 2.720108714724091e-12
C44_51 V44 V51 2.6681090876384584e-19

R44_52 V44 V52 45617.20866837687
L44_52 V44 V52 2.113346937589094e-12
C44_52 V44 V52 2.297953842686712e-19

R44_53 V44 V53 4373.4553725229725
L44_53 V44 V53 -3.2225918104182414e-12
C44_53 V44 V53 -2.9104021460232564e-19

R44_54 V44 V54 12724.856677112983
L44_54 V44 V54 -1.7222889747458467e-12
C44_54 V44 V54 -4.029564723671582e-19

R44_55 V44 V55 5678.456666253652
L44_55 V44 V55 -1.834231185682835e-12
C44_55 V44 V55 -3.7468036898783154e-19

R44_56 V44 V56 4129.106155109492
L44_56 V44 V56 -7.450210648167949e-13
C44_56 V44 V56 -9.197414499230537e-19

R44_57 V44 V57 15896.763113989768
L44_57 V44 V57 -5.93404393559816e-12
C44_57 V44 V57 1.1133494139716125e-19

R44_58 V44 V58 -5916.023344017794
L44_58 V44 V58 -7.534563519289372e-12
C44_58 V44 V58 -3.3629318289114125e-20

R44_59 V44 V59 -28336.214538873308
L44_59 V44 V59 -9.991404366582758e-12
C44_59 V44 V59 7.765287806222965e-20

R44_60 V44 V60 -4768.327985400373
L44_60 V44 V60 9.63816468739033e-12
C44_60 V44 V60 3.2058251340657103e-19

R44_61 V44 V61 -5989.5404792802465
L44_61 V44 V61 3.1480551494903673e-12
C44_61 V44 V61 1.0481848835158102e-19

R44_62 V44 V62 16443.424820246248
L44_62 V44 V62 2.6113302571628914e-12
C44_62 V44 V62 3.1654515035763594e-19

R44_63 V44 V63 -27858.460879999882
L44_63 V44 V63 5.048555482013243e-12
C44_63 V44 V63 1.4056539241442166e-19

R44_64 V44 V64 -7373.795183145412
L44_64 V44 V64 2.4713404213597483e-12
C44_64 V44 V64 8.232901064833713e-20

R44_65 V44 V65 9486.974276745008
L44_65 V44 V65 5.3468438706076856e-12
C44_65 V44 V65 4.2908067557649675e-20

R44_66 V44 V66 59055.545007901506
L44_66 V44 V66 1.2795653714173146e-11
C44_66 V44 V66 8.343825379026483e-21

R44_67 V44 V67 -29480.54165373768
L44_67 V44 V67 2.7026393416115047e-11
C44_67 V44 V67 -4.0465569274074686e-20

R44_68 V44 V68 68484.58819376338
L44_68 V44 V68 4.638396490677535e-12
C44_68 V44 V68 -6.723795011903153e-20

R44_69 V44 V69 4120.1569200058475
L44_69 V44 V69 -3.665805889434435e-12
C44_69 V44 V69 -2.1612883191425615e-19

R44_70 V44 V70 -10614.102361826324
L44_70 V44 V70 -5.535177072118003e-12
C44_70 V44 V70 -1.699540861833238e-19

R44_71 V44 V71 -7156.196068117922
L44_71 V44 V71 1.4181051187579268e-11
C44_71 V44 V71 1.1271942344609635e-20

R44_72 V44 V72 -12919.323435000304
L44_72 V44 V72 -1.3952961662820055e-11
C44_72 V44 V72 5.0910898780229915e-20

R44_73 V44 V73 12068.037650288605
L44_73 V44 V73 1.9470855098318756e-11
C44_73 V44 V73 8.141719634620326e-20

R44_74 V44 V74 33320.574603218134
L44_74 V44 V74 -1.994646091043503e-11
C44_74 V44 V74 6.303631272531796e-20

R44_75 V44 V75 22908.485965811058
L44_75 V44 V75 -5.459001747806241e-12
C44_75 V44 V75 -1.9901975390880954e-20

R44_76 V44 V76 24959.92541487336
L44_76 V44 V76 -1.5214500127564278e-12
C44_76 V44 V76 -2.9944902503316624e-19

R44_77 V44 V77 -22178.3632571255
L44_77 V44 V77 2.386384770738626e-11
C44_77 V44 V77 1.981605114133322e-19

R44_78 V44 V78 -159984.6440781471
L44_78 V44 V78 6.652015160594622e-12
C44_78 V44 V78 -5.720839085705368e-20

R44_79 V44 V79 4120.772070736581
L44_79 V44 V79 1.1003324820204283e-10
C44_79 V44 V79 -1.3621990697638296e-21

R44_80 V44 V80 6841.08789450108
L44_80 V44 V80 1.319710669167227e-12
C44_80 V44 V80 2.9386250409507315e-19

R44_81 V44 V81 3332.6126763131097
L44_81 V44 V81 3.317181675245026e-12
C44_81 V44 V81 -1.063932257836775e-20

R44_82 V44 V82 33351.75894679782
L44_82 V44 V82 1.4596390339936413e-11
C44_82 V44 V82 1.4015063573730626e-19

R44_83 V44 V83 -9627.798142508856
L44_83 V44 V83 7.317515388968184e-12
C44_83 V44 V83 1.6239055611264966e-19

R44_84 V44 V84 -10125.51885210367
L44_84 V44 V84 1.0284808462051649e-11
C44_84 V44 V84 2.501366809448973e-20

R44_85 V44 V85 94666.46117118934
L44_85 V44 V85 -1.9521616410826337e-11
C44_85 V44 V85 -6.358386258690377e-20

R44_86 V44 V86 -4480.923932974964
L44_86 V44 V86 -8.51677649152309e-12
C44_86 V44 V86 4.757167595494918e-20

R44_87 V44 V87 -2215.2247355496447
L44_87 V44 V87 -2.6472771463306575e-12
C44_87 V44 V87 -2.1000459635827942e-19

R44_88 V44 V88 -1997.9522982906337
L44_88 V44 V88 -9.939777447902253e-13
C44_88 V44 V88 -4.247376727509349e-19

R44_89 V44 V89 8522.016739914072
L44_89 V44 V89 -5.552927823879284e-12
C44_89 V44 V89 -1.3833214893970083e-19

R44_90 V44 V90 -30536.495091828
L44_90 V44 V90 -5.3574556071943246e-12
C44_90 V44 V90 -2.4317886919605473e-19

R44_91 V44 V91 2924.97337039983
L44_91 V44 V91 2.1340285927533166e-12
C44_91 V44 V91 1.847500478009309e-19

R44_92 V44 V92 2215.787261229771
L44_92 V44 V92 5.859542645453744e-13
C44_92 V44 V92 6.238778102710314e-19

R44_93 V44 V93 -28346.820375356976
L44_93 V44 V93 -8.111510159500057e-12
C44_93 V44 V93 4.293728589157584e-20

R44_94 V44 V94 3694.2175085679237
L44_94 V44 V94 -1.6251098079462397e-11
C44_94 V44 V94 7.994805048114569e-20

R44_95 V44 V95 2152.2908557278674
L44_95 V44 V95 6.516388696513076e-12
C44_95 V44 V95 1.2280445544664677e-19

R44_96 V44 V96 1723.8667644160946
L44_96 V44 V96 -5.515772556432892e-12
C44_96 V44 V96 -5.65855660491688e-20

R44_97 V44 V97 1979.4278760418931
L44_97 V44 V97 2.4682242605473984e-12
C44_97 V44 V97 4.420871767020003e-19

R44_98 V44 V98 -4886.345971862759
L44_98 V44 V98 2.2837582750063486e-12
C44_98 V44 V98 2.7777352410893194e-19

R44_99 V44 V99 -1338.9790956800848
L44_99 V44 V99 -1.4927739256339733e-12
C44_99 V44 V99 -1.8312641899042845e-19

R44_100 V44 V100 -1092.3106353485507
L44_100 V44 V100 -5.962980557782898e-13
C44_100 V44 V100 -7.075005414949119e-19

R44_101 V44 V101 10512.243334814315
L44_101 V44 V101 5.604169376016716e-12
C44_101 V44 V101 -1.857242392603652e-19

R44_102 V44 V102 -5891.90494493747
L44_102 V44 V102 -7.501049222121305e-12
C44_102 V44 V102 -9.099549581668044e-20

R44_103 V44 V103 -31953.021857094882
L44_103 V44 V103 2.7057820520536817e-11
C44_103 V44 V103 1.858927542410229e-20

R44_104 V44 V104 -3014.5914924277063
L44_104 V44 V104 8.336056957642143e-13
C44_104 V44 V104 6.697806147580783e-19

R44_105 V44 V105 -5848.739090929073
L44_105 V44 V105 -1.868859271666756e-12
C44_105 V44 V105 -2.3787395741314945e-19

R44_106 V44 V106 -4482.129633184602
L44_106 V44 V106 -1.456813407579533e-12
C44_106 V44 V106 -3.5124894482874757e-19

R44_107 V44 V107 2816.385937149016
L44_107 V44 V107 2.533710727107766e-12
C44_107 V44 V107 9.858883273635247e-20

R44_108 V44 V108 1415.7505468569661
L44_108 V44 V108 4.094682158461758e-12
C44_108 V44 V108 -2.0023069611728507e-19

R44_109 V44 V109 -14924.022807720865
L44_109 V44 V109 1.0701469625340784e-11
C44_109 V44 V109 2.6537931235319126e-19

R44_110 V44 V110 2840.3655857847098
L44_110 V44 V110 2.4417582118752683e-12
C44_110 V44 V110 1.2580806044296856e-19

R44_111 V44 V111 -2769.164700946768
L44_111 V44 V111 -1.1269287595941304e-11
C44_111 V44 V111 -2.806857095045852e-20

R44_112 V44 V112 -6377.326097314028
L44_112 V44 V112 -2.3411962532698102e-12
C44_112 V44 V112 1.013849694428289e-21

R44_113 V44 V113 1416.7745654831854
L44_113 V44 V113 1.2688920072607586e-12
C44_113 V44 V113 1.5301876671369785e-19

R44_114 V44 V114 6587.441833480261
L44_114 V44 V114 1.7875114845291606e-12
C44_114 V44 V114 3.2295668346891104e-19

R44_115 V44 V115 7719.019536643459
L44_115 V44 V115 -3.9634360939750116e-12
C44_115 V44 V115 -4.6800424078052004e-20

R44_116 V44 V116 -3668.219877187436
L44_116 V44 V116 -1.5394753321762132e-12
C44_116 V44 V116 1.0029486520270173e-19

R44_117 V44 V117 2024.710522374669
L44_117 V44 V117 -2.7527569789743326e-12
C44_117 V44 V117 -1.5516619981773827e-19

R44_118 V44 V118 -1697.8131215406536
L44_118 V44 V118 -1.2538052323973918e-12
C44_118 V44 V118 -2.959119404228313e-19

R44_119 V44 V119 -5631.518421378027
L44_119 V44 V119 -1.2995021408045773e-11
C44_119 V44 V119 -2.0368584848791805e-19

R44_120 V44 V120 -58704.787089437326
L44_120 V44 V120 1.7502180065502593e-12
C44_120 V44 V120 -4.1961962915509574e-19

R44_121 V44 V121 -1450.9525497067934
L44_121 V44 V121 -3.0430594387604837e-12
C44_121 V44 V121 -1.3161265942213931e-20

R44_122 V44 V122 10902.992828536799
L44_122 V44 V122 3.532034262080957e-11
C44_122 V44 V122 -9.753167542325408e-20

R44_123 V44 V123 -9881.465775724388
L44_123 V44 V123 4.672727983439329e-12
C44_123 V44 V123 2.0936638366698035e-19

R44_124 V44 V124 -558657.2623761299
L44_124 V44 V124 1.7707287271107672e-12
C44_124 V44 V124 6.761315259931059e-19

R44_125 V44 V125 -1902.5281957383668
L44_125 V44 V125 2.3297744825959328e-12
C44_125 V44 V125 1.6189702943046237e-20

R44_126 V44 V126 3691.4908335563096
L44_126 V44 V126 1.0167044594010571e-12
C44_126 V44 V126 1.6254018842746725e-19

R44_127 V44 V127 2548.982380536762
L44_127 V44 V127 1.7928632780077498e-12
C44_127 V44 V127 1.77651822867986e-19

R44_128 V44 V128 3011.888076010521
L44_128 V44 V128 -1.4280320759897758e-12
C44_128 V44 V128 -1.5081856472321333e-19

R44_129 V44 V129 768.5790483024701
L44_129 V44 V129 6.823752915706189e-12
C44_129 V44 V129 6.544781806595602e-20

R44_130 V44 V130 30649.087626433757
L44_130 V44 V130 -1.8480446936943745e-12
C44_130 V44 V130 -3.574115890198422e-20

R44_131 V44 V131 -2708.265134821782
L44_131 V44 V131 -1.3899434937419078e-12
C44_131 V44 V131 -3.196948022141484e-19

R44_132 V44 V132 -2940.7741788347066
L44_132 V44 V132 -1.592924946695585e-11
C44_132 V44 V132 -3.443935640422799e-19

R44_133 V44 V133 2672.0671439784683
L44_133 V44 V133 -8.411975093606352e-12
C44_133 V44 V133 -3.6625910343983977e-20

R44_134 V44 V134 -2216.358902818195
L44_134 V44 V134 -5.180717582069611e-12
C44_134 V44 V134 -2.322527413964475e-19

R44_135 V44 V135 -2609.8996930380035
L44_135 V44 V135 -8.747374782826891e-12
C44_135 V44 V135 3.4718285226894213e-20

R44_136 V44 V136 -1858.5647741603923
L44_136 V44 V136 2.9190410513354817e-12
C44_136 V44 V136 6.772668256876864e-19

R44_137 V44 V137 -695.6124335910415
L44_137 V44 V137 -1.208447566111092e-11
C44_137 V44 V137 6.822203215210441e-20

R44_138 V44 V138 2777.1252167525568
L44_138 V44 V138 1.9076894176314117e-12
C44_138 V44 V138 2.287240197817104e-19

R44_139 V44 V139 1440.0619093152493
L44_139 V44 V139 1.6468822270452136e-12
C44_139 V44 V139 2.4382920111400142e-20

R44_140 V44 V140 2240.690029836708
L44_140 V44 V140 -1.2865548395966521e-11
C44_140 V44 V140 -7.646525964104561e-19

R44_141 V44 V141 -2359.0890317809094
L44_141 V44 V141 -2.309580037161804e-11
C44_141 V44 V141 6.012693116365205e-20

R44_142 V44 V142 2063.587821623679
L44_142 V44 V142 1.2957336049989016e-11
C44_142 V44 V142 5.301820048056933e-20

R44_143 V44 V143 -17913.624168661107
L44_143 V44 V143 -1.3043957254768353e-11
C44_143 V44 V143 4.067404652402755e-20

R44_144 V44 V144 1016.1213569822868
L44_144 V44 V144 3.75095348600763e-11
C44_144 V44 V144 9.845173050642881e-20

R44_145 V44 V145 457.21075161930713
L44_145 V44 V145 3.50856283821327e-12
C44_145 V44 V145 -1.483523756745872e-20

R44_146 V44 V146 5123.8782505024965
L44_146 V44 V146 -1.946750988000456e-12
C44_146 V44 V146 -1.1152926755155224e-19

R44_147 V44 V147 2954.07589313628
L44_147 V44 V147 -7.248132001168726e-12
C44_147 V44 V147 1.4876900584532174e-19

R44_148 V44 V148 -1097.1151476530222
L44_148 V44 V148 4.468991365405401e-12
C44_148 V44 V148 5.08319827677092e-19

R44_149 V44 V149 -2023.514141045372
L44_149 V44 V149 8.237333764309395e-12
C44_149 V44 V149 -1.7057196799952152e-19

R44_150 V44 V150 -674.5546601266268
L44_150 V44 V150 4.5915799837698146e-12
C44_150 V44 V150 4.5942640433467365e-20

R44_151 V44 V151 -971.1402196441882
L44_151 V44 V151 -8.145735621715617e-12
C44_151 V44 V151 -6.58345038269805e-20

R44_152 V44 V152 -836.3989544622438
L44_152 V44 V152 -4.4105134894507645e-12
C44_152 V44 V152 -1.8173926289268276e-19

R44_153 V44 V153 -871.9548635201763
L44_153 V44 V153 -2.6422012221902e-12
C44_153 V44 V153 4.986432858424829e-20

R44_154 V44 V154 -4502.925878157082
L44_154 V44 V154 -5.8055035440354545e-12
C44_154 V44 V154 5.440618993915802e-20

R44_155 V44 V155 599.649995784244
L44_155 V44 V155 -6.1761328057815065e-12
C44_155 V44 V155 -1.1866796161243042e-19

R44_156 V44 V156 2736.238453041568
L44_156 V44 V156 -3.849461205727504e-12
C44_156 V44 V156 -3.5204771908555458e-19

R44_157 V44 V157 -7722.085819440539
L44_157 V44 V157 -6.046000317295839e-12
C44_157 V44 V157 3.0805841473008545e-19

R44_158 V44 V158 2983.0327597412615
L44_158 V44 V158 2.461909579021203e-11
C44_158 V44 V158 -4.389378271100433e-20

R44_159 V44 V159 -1134.456092269683
L44_159 V44 V159 -1.2802282540249007e-11
C44_159 V44 V159 8.256196270517023e-20

R44_160 V44 V160 536.0826072668189
L44_160 V44 V160 3.708236074000554e-12
C44_160 V44 V160 3.0226353482168866e-19

R44_161 V44 V161 2038.4745104555132
L44_161 V44 V161 9.588751886586038e-12
C44_161 V44 V161 -2.441364493894492e-19

R44_162 V44 V162 2222.5806219477427
L44_162 V44 V162 -1.7807295554272532e-11
C44_162 V44 V162 -5.12911680846719e-20

R44_163 V44 V163 -3306.2339663734933
L44_163 V44 V163 5.439414589842826e-12
C44_163 V44 V163 -1.9476007957992242e-21

R44_164 V44 V164 -852.0312500353759
L44_164 V44 V164 1.7707774589057779e-12
C44_164 V44 V164 -1.8848085734719373e-19

R44_165 V44 V165 1426.4526978448396
L44_165 V44 V165 1.474247087143477e-12
C44_165 V44 V165 5.921964356037233e-20

R44_166 V44 V166 -1121.604673087071
L44_166 V44 V166 4.149570626934842e-12
C44_166 V44 V166 1.0399355325926128e-19

R44_167 V44 V167 28220.850026423122
L44_167 V44 V167 -1.225481700020777e-09
C44_167 V44 V167 -7.329056928113554e-20

R44_168 V44 V168 -2396.972517782109
L44_168 V44 V168 -1.599437888351843e-12
C44_168 V44 V168 -1.269852459692619e-19

R44_169 V44 V169 -1545.8744424966521
L44_169 V44 V169 -2.574767080432456e-12
C44_169 V44 V169 2.3361478624969623e-19

R44_170 V44 V170 4146.675468327443
L44_170 V44 V170 -3.1543793758680915e-12
C44_170 V44 V170 -5.845381971510329e-20

R44_171 V44 V171 1386.4192858936112
L44_171 V44 V171 -3.322648062015693e-12
C44_171 V44 V171 -7.645903056213881e-21

R44_172 V44 V172 1160.1850571946682
L44_172 V44 V172 -7.797183020985135e-12
C44_172 V44 V172 1.3360456394996873e-19

R44_173 V44 V173 15811.146723516296
L44_173 V44 V173 -2.7708517332758894e-12
C44_173 V44 V173 -6.191994813282238e-20

R44_174 V44 V174 1919.4374896368047
L44_174 V44 V174 -6.2471413335896385e-12
C44_174 V44 V174 9.060862038141015e-20

R44_175 V44 V175 -1357.928895665208
L44_175 V44 V175 -2.003279193690594e-11
C44_175 V44 V175 3.365315736448497e-20

R44_176 V44 V176 -11495.475841469559
L44_176 V44 V176 1.2026322471499806e-11
C44_176 V44 V176 -2.596622636893031e-19

R44_177 V44 V177 3981.9157701027375
L44_177 V44 V177 2.089795961518875e-12
C44_177 V44 V177 -2.9581614270231834e-20

R44_178 V44 V178 -2322.7448079477886
L44_178 V44 V178 3.1244603320178577e-12
C44_178 V44 V178 7.820237098394495e-21

R44_179 V44 V179 1865.8907390800885
L44_179 V44 V179 4.120190301639143e-12
C44_179 V44 V179 8.637566155674328e-20

R44_180 V44 V180 -2976.9566167616285
L44_180 V44 V180 1.195305984235805e-12
C44_180 V44 V180 2.498773249058673e-19

R44_181 V44 V181 -2595.1359763042005
L44_181 V44 V181 -1.5367210954188088e-11
C44_181 V44 V181 -5.127716654238608e-20

R44_182 V44 V182 52784.33035838438
L44_182 V44 V182 -7.268446214030524e-12
C44_182 V44 V182 -3.2056717087082306e-21

R44_183 V44 V183 -6162.308803029956
L44_183 V44 V183 3.671120220843254e-12
C44_183 V44 V183 5.716552169333038e-20

R44_184 V44 V184 2402.378603753592
L44_184 V44 V184 -2.8753052828235497e-12
C44_184 V44 V184 -8.381944281100389e-20

R44_185 V44 V185 7066.599998347383
L44_185 V44 V185 -2.4346345109011316e-12
C44_185 V44 V185 4.1613795076660244e-20

R44_186 V44 V186 1981.9145737335655
L44_186 V44 V186 7.538936576559129e-11
C44_186 V44 V186 -7.22053647467622e-20

R44_187 V44 V187 8379.626760183153
L44_187 V44 V187 -1.6538976878899452e-11
C44_187 V44 V187 -1.732062691795132e-19

R44_188 V44 V188 21157.148857688117
L44_188 V44 V188 -1.2758135333694175e-12
C44_188 V44 V188 -1.740263817863974e-19

R44_189 V44 V189 -3521.8361506095343
L44_189 V44 V189 3.87755686161634e-12
C44_189 V44 V189 8.257044341331635e-20

R44_190 V44 V190 -2780.158129671967
L44_190 V44 V190 6.187810746325118e-12
C44_190 V44 V190 3.872880385375947e-20

R44_191 V44 V191 -5368.666683564311
L44_191 V44 V191 -2.3365418067250776e-12
C44_191 V44 V191 3.9951021668618354e-21

R44_192 V44 V192 -10602.130834996211
L44_192 V44 V192 1.0089796325416752e-12
C44_192 V44 V192 3.337570480951668e-19

R44_193 V44 V193 2553.7179210902004
L44_193 V44 V193 2.1796959072283636e-12
C44_193 V44 V193 7.48458406957896e-20

R44_194 V44 V194 -2356.029875743756
L44_194 V44 V194 -2.8527196275898407e-11
C44_194 V44 V194 2.684039728103522e-19

R44_195 V44 V195 -8506.476618399909
L44_195 V44 V195 1.883876395472986e-12
C44_195 V44 V195 2.1265953684212905e-19

R44_196 V44 V196 -2598.582297325014
L44_196 V44 V196 -9.680505097272768e-13
C44_196 V44 V196 -4.982711254601087e-19

R44_197 V44 V197 -24410.376376325054
L44_197 V44 V197 -2.378272060231545e-12
C44_197 V44 V197 -2.0144156396476513e-19

R44_198 V44 V198 145598.36543554597
L44_198 V44 V198 -6.58174800446463e-12
C44_198 V44 V198 3.820756850590997e-20

R44_199 V44 V199 9893.603196831842
L44_199 V44 V199 -8.592182735186725e-12
C44_199 V44 V199 -6.454004097032465e-20

R44_200 V44 V200 2067.3018936654103
L44_200 V44 V200 1.1682840641897464e-11
C44_200 V44 V200 1.0165250322097995e-20

R45_45 V45 0 144.4065596422565
L45_45 V45 0 1.729840960334153e-13
C45_45 V45 0 1.6048263344598741e-18

R45_46 V45 V46 -4912.989830550319
L45_46 V45 V46 -2.4655720014295494e-12
C45_46 V45 V46 -1.3895668434413323e-19

R45_47 V45 V47 -10973.889100957304
L45_47 V45 V47 -2.092478924449414e-12
C45_47 V45 V47 -2.1011254754403624e-19

R45_48 V45 V48 -3324.882672223139
L45_48 V45 V48 -1.354130335223129e-12
C45_48 V45 V48 -2.816945787015271e-19

R45_49 V45 V49 -1269.0910289146607
L45_49 V45 V49 2.8369625383028033e-12
C45_49 V45 V49 3.0904284387166984e-19

R45_50 V45 V50 16968.20102143802
L45_50 V45 V50 -6.6270407142794945e-12
C45_50 V45 V50 -1.2830974008748055e-19

R45_51 V45 V51 -125966.55031066935
L45_51 V45 V51 -5.3990893612008565e-12
C45_51 V45 V51 -3.9817573015787766e-20

R45_52 V45 V52 9661.59433396721
L45_52 V45 V52 -9.411226633151645e-12
C45_52 V45 V52 5.77715149749577e-21

R45_53 V45 V53 -2980.507977282525
L45_53 V45 V53 4.762241984787889e-12
C45_53 V45 V53 3.888660137310294e-19

R45_54 V45 V54 -95932.06133903461
L45_54 V45 V54 6.880495477499385e-12
C45_54 V45 V54 1.7168776914390358e-19

R45_55 V45 V55 -10935.338957647813
L45_55 V45 V55 1.5056159929613432e-11
C45_55 V45 V55 1.172254806304019e-19

R45_56 V45 V56 10991.900722340792
L45_56 V45 V56 3.223294481071e-12
C45_56 V45 V56 2.383960262226917e-19

R45_57 V45 V57 4573.165404848299
L45_57 V45 V57 8.678562059665242e-13
C45_57 V45 V57 2.194297987611137e-19

R45_58 V45 V58 4923.7790326473905
L45_58 V45 V58 1.822312394529711e-12
C45_58 V45 V58 1.6056620257366374e-19

R45_59 V45 V59 2862.2383742368675
L45_59 V45 V59 2.726720091065772e-12
C45_59 V45 V59 5.717423742313305e-21

R45_60 V45 V60 1925.1112953950876
L45_60 V45 V60 1.6278082184997388e-12
C45_60 V45 V60 7.462319129603444e-20

R45_61 V45 V61 3252.4615966427336
L45_61 V45 V61 -1.1041362751813447e-12
C45_61 V45 V61 -4.735927870296673e-19

R45_62 V45 V62 40906.80053131608
L45_62 V45 V62 -1.0398532202078219e-11
C45_62 V45 V62 -1.3098559400019358e-19

R45_63 V45 V63 422456.2432203227
L45_63 V45 V63 4.074601772018896e-12
C45_63 V45 V63 7.89769567553983e-20

R45_64 V45 V64 -7699.643793871826
L45_64 V45 V64 -6.313303016749348e-10
C45_64 V45 V64 -5.706647916875601e-22

R45_65 V45 V65 -999.4820568230383
L45_65 V45 V65 -1.0528968721487172e-12
C45_65 V45 V65 -4.0662567423647956e-19

R45_66 V45 V66 -35823.80009336553
L45_66 V45 V66 -3.0889392496736113e-12
C45_66 V45 V66 -1.8698443485176528e-19

R45_67 V45 V67 -78029.38976285778
L45_67 V45 V67 -2.597318167725085e-12
C45_67 V45 V67 -1.3483384104575219e-19

R45_68 V45 V68 -6030.531445034525
L45_68 V45 V68 -1.2007694571423035e-12
C45_68 V45 V68 -3.054210338594014e-19

R45_69 V45 V69 -1283.688075718071
L45_69 V45 V69 2.2190984237447583e-12
C45_69 V45 V69 5.499264723810678e-19

R45_70 V45 V70 5958.236827852131
L45_70 V45 V70 1.0599076614732637e-11
C45_70 V45 V70 9.848746314234643e-20

R45_71 V45 V71 6791.561189565886
L45_71 V45 V71 -3.097808893948042e-12
C45_71 V45 V71 -1.5471883528424813e-19

R45_72 V45 V72 4560.2268382787115
L45_72 V45 V72 -7.973864637235719e-12
C45_72 V45 V72 -4.840797400318578e-20

R45_73 V45 V73 3194.4628389756617
L45_73 V45 V73 -4.9608441373009165e-12
C45_73 V45 V73 -1.1885639217156383e-19

R45_74 V45 V74 13580.384843827223
L45_74 V45 V74 2.0579679060498386e-12
C45_74 V45 V74 2.507905858227979e-19

R45_75 V45 V75 -7124.5903217811065
L45_75 V45 V75 1.9280548678885833e-12
C45_75 V45 V75 2.3774531001913604e-19

R45_76 V45 V76 8120.493671408892
L45_76 V45 V76 9.370806541361743e-13
C45_76 V45 V76 4.7805303073514225e-19

R45_77 V45 V77 1325.5470495023715
L45_77 V45 V77 1.5974870088325582e-12
C45_77 V45 V77 2.6083360394553234e-20

R45_78 V45 V78 -2203.8479562136313
L45_78 V45 V78 -7.775137175808352e-12
C45_78 V45 V78 -7.934384849666049e-20

R45_79 V45 V79 -7802.89151532816
L45_79 V45 V79 5.6886272644914355e-12
C45_79 V45 V79 4.175736664738777e-20

R45_80 V45 V80 -3499.00621371226
L45_80 V45 V80 -4.810381086819966e-12
C45_80 V45 V80 -1.4729921004514204e-19

R45_81 V45 V81 -370.38596196104317
L45_81 V45 V81 -1.199724173050066e-12
C45_81 V45 V81 -2.5325656480558423e-19

R45_82 V45 V82 2726.813071969202
L45_82 V45 V82 -2.6475572554360094e-12
C45_82 V45 V82 -2.693443047515639e-19

R45_83 V45 V83 1476.5067430030151
L45_83 V45 V83 -4.1554801987055335e-12
C45_83 V45 V83 -1.574462076297296e-19

R45_84 V45 V84 2103.0408101839384
L45_84 V45 V84 -1.6016851651667267e-12
C45_84 V45 V84 -3.277934723295614e-19

R45_85 V45 V85 3312.5061890702605
L45_85 V45 V85 -3.1186271849692587e-12
C45_85 V45 V85 -2.1078478089568631e-19

R45_86 V45 V86 871.4161062850978
L45_86 V45 V86 -2.74477109871944e-11
C45_86 V45 V86 -5.1219507928746435e-20

R45_87 V45 V87 3754.602422383755
L45_87 V45 V87 3.4493290619568478e-12
C45_87 V45 V87 1.7345955815149522e-19

R45_88 V45 V88 2535.354680784873
L45_88 V45 V88 2.26453742043337e-12
C45_88 V45 V88 2.6687565825539785e-19

R45_89 V45 V89 1535.8083024709645
L45_89 V45 V89 -2.718183655796042e-12
C45_89 V45 V89 1.4311797617887347e-19

R45_90 V45 V90 -1046.9202371696615
L45_90 V45 V90 1.5402808241099602e-12
C45_90 V45 V90 4.559276526283198e-19

R45_91 V45 V91 -1029.181172036409
L45_91 V45 V91 -1.0906237928211467e-12
C45_91 V45 V91 -3.567804265592347e-19

R45_92 V45 V92 -1676.0645058305035
L45_92 V45 V92 -1.7488244599236967e-12
C45_92 V45 V92 -1.6344218666391938e-19

R45_93 V45 V93 -545.5019679006673
L45_93 V45 V93 1.5247343575453917e-12
C45_93 V45 V93 2.669280490958374e-19

R45_94 V45 V94 -2269.4820070300234
L45_94 V45 V94 -8.153437879870937e-12
C45_94 V45 V94 -8.862294225671856e-20

R45_95 V45 V95 28403.572404509534
L45_95 V45 V95 4.056959204760379e-12
C45_95 V45 V95 2.2564881371720193e-20

R45_96 V45 V96 -12549.627456405547
L45_96 V45 V96 2.960047273748534e-12
C45_96 V45 V96 -9.961570232098277e-21

R45_97 V45 V97 -3799.0737882069607
L45_97 V45 V97 -2.2442619250746137e-12
C45_97 V45 V97 -3.430854154185506e-19

R45_98 V45 V98 741.9724265034424
L45_98 V45 V98 -1.7623215440907475e-12
C45_98 V45 V98 -4.1103757294474365e-19

R45_99 V45 V99 678.9744822312846
L45_99 V45 V99 9.837174915028584e-13
C45_99 V45 V99 4.421943931108671e-19

R45_100 V45 V100 807.6683140449351
L45_100 V45 V100 1.7656750859262606e-12
C45_100 V45 V100 2.6595922916647694e-19

R45_101 V45 V101 960.3801075379594
L45_101 V45 V101 5.647803667873594e-11
C45_101 V45 V101 2.9323157769054164e-20

R45_102 V45 V102 18361.069271743636
L45_102 V45 V102 1.970849607923261e-12
C45_102 V45 V102 3.014085489899634e-19

R45_103 V45 V103 -4005.558386848492
L45_103 V45 V103 -2.8612250083492807e-12
C45_103 V45 V103 -1.2418480984458452e-19

R45_104 V45 V104 -11488.312432407285
L45_104 V45 V104 -2.5722321910011335e-12
C45_104 V45 V104 -1.4738127595799896e-19

R45_105 V45 V105 -324.7498114650683
L45_105 V45 V105 -3.2949558865116444e-12
C45_105 V45 V105 -4.55414894973942e-20

R45_106 V45 V106 -5989.4014506465055
L45_106 V45 V106 2.5713868025031303e-12
C45_106 V45 V106 1.8675473169231776e-19

R45_107 V45 V107 -3239.6458744937095
L45_107 V45 V107 -1.8513222707525555e-12
C45_107 V45 V107 -2.9832223010093013e-19

R45_108 V45 V108 -4020.935676677595
L45_108 V45 V108 -4.99076883613224e-12
C45_108 V45 V108 -8.84825183432061e-20

R45_109 V45 V109 2152.551947737529
L45_109 V45 V109 -1.2487227840655368e-12
C45_109 V45 V109 -2.9353124214706887e-19

R45_110 V45 V110 5978.854010517605
L45_110 V45 V110 -2.2734614528325103e-12
C45_110 V45 V110 -2.3867603231044835e-19

R45_111 V45 V111 24472.10099918395
L45_111 V45 V111 -9.281687050746691e-12
C45_111 V45 V111 3.35126973524387e-20

R45_112 V45 V112 10283.97165741719
L45_112 V45 V112 -1.0029959780581613e-11
C45_112 V45 V112 -1.4697466730926537e-21

R45_113 V45 V113 1527.0563440250505
L45_113 V45 V113 1.4829618738550379e-12
C45_113 V45 V113 3.7024529550993063e-19

R45_114 V45 V114 5340.542364968979
L45_114 V45 V114 -3.072409452144334e-12
C45_114 V45 V114 -1.4573529078078814e-19

R45_115 V45 V115 2422.1192427478136
L45_115 V45 V115 1.6309619148068125e-12
C45_115 V45 V115 2.33112293961311e-19

R45_116 V45 V116 3256.0327524909594
L45_116 V45 V116 1.9558575641784447e-12
C45_116 V45 V116 1.335922568466268e-19

R45_117 V45 V117 -751.3381080318586
L45_117 V45 V117 1.9445964106834306e-12
C45_117 V45 V117 7.504951662779745e-20

R45_118 V45 V118 -4416.519918685097
L45_118 V45 V118 1.9090926531905703e-12
C45_118 V45 V118 2.698611590763755e-19

R45_119 V45 V119 9178.278883158468
L45_119 V45 V119 -1.503760317538108e-11
C45_119 V45 V119 -1.2911650209378204e-21

R45_120 V45 V120 3916.12698831202
L45_120 V45 V120 -6.631687741247047e-11
C45_120 V45 V120 9.422983927635321e-20

R45_121 V45 V121 -3630.4757542532457
L45_121 V45 V121 -1.2082062792972019e-12
C45_121 V45 V121 -2.85544132225267e-19

R45_122 V45 V122 3447.334980078746
L45_122 V45 V122 -1.0883430904657196e-10
C45_122 V45 V122 -2.2770057136430568e-20

R45_123 V45 V123 -4307.513210279288
L45_123 V45 V123 -1.0482673664251363e-11
C45_123 V45 V123 -8.20743079400681e-20

R45_124 V45 V124 -2640.463961991108
L45_124 V45 V124 -2.894004555655159e-12
C45_124 V45 V124 -2.3898277852651957e-19

R45_125 V45 V125 -808.8139958603381
L45_125 V45 V125 -1.550013247326763e-12
C45_125 V45 V125 -1.2607997219725335e-19

R45_126 V45 V126 26719.518218797868
L45_126 V45 V126 -1.5280770138537426e-12
C45_126 V45 V126 -2.450229591938229e-19

R45_127 V45 V127 9411.551050832322
L45_127 V45 V127 -5.6420528991806916e-12
C45_127 V45 V127 -1.2599124829030377e-19

R45_128 V45 V128 -21431.47580967457
L45_128 V45 V128 -5.760144618944821e-12
C45_128 V45 V128 -1.1918571794955532e-19

R45_129 V45 V129 2138.676925532871
L45_129 V45 V129 8.07072098594278e-12
C45_129 V45 V129 -1.3734157784446156e-19

R45_130 V45 V130 22314.79157587527
L45_130 V45 V130 1.8121313830678181e-12
C45_130 V45 V130 2.0092719641753697e-19

R45_131 V45 V131 36410.23371742154
L45_131 V45 V131 9.98764747928702e-12
C45_131 V45 V131 1.5617438687498472e-19

R45_132 V45 V132 2082.7708742213003
L45_132 V45 V132 2.2377032112286596e-12
C45_132 V45 V132 3.5603671925608784e-19

R45_133 V45 V133 1072.4538036503952
L45_133 V45 V133 1.6924781351665092e-12
C45_133 V45 V133 5.018363191151822e-19

R45_134 V45 V134 3991.0132352990026
L45_134 V45 V134 -1.027510486575744e-11
C45_134 V45 V134 -2.6000818954067166e-20

R45_135 V45 V135 -3481.1763605397596
L45_135 V45 V135 1.1013037138919505e-11
C45_135 V45 V135 -1.4190766547257285e-20

R45_136 V45 V136 -1867.6129535561256
L45_136 V45 V136 -2.133596574787544e-11
C45_136 V45 V136 -1.3510797747933931e-19

R45_137 V45 V137 -580.351514744077
L45_137 V45 V137 1.8098611445730762e-12
C45_137 V45 V137 1.7293035202134892e-19

R45_138 V45 V138 -1386.6437195463168
L45_138 V45 V138 -4.935449541245512e-12
C45_138 V45 V138 -4.0970084430532875e-20

R45_139 V45 V139 1744.5038549283554
L45_139 V45 V139 5.385984438721628e-11
C45_139 V45 V139 1.4233600616629743e-19

R45_140 V45 V140 1997.790292935011
L45_140 V45 V140 5.897899951589314e-12
C45_140 V45 V140 2.599592503322741e-19

R45_141 V45 V141 2035.3192673754102
L45_141 V45 V141 -7.518776805494231e-13
C45_141 V45 V141 -8.044136857703417e-19

R45_142 V45 V142 968.290050576084
L45_142 V45 V142 1.2132867719706572e-11
C45_142 V45 V142 -5.290828772353037e-20

R45_143 V45 V143 5648.228586738471
L45_143 V45 V143 -3.55959227632414e-11
C45_143 V45 V143 -1.121093553595473e-19

R45_144 V45 V144 1421.7554363218344
L45_144 V45 V144 -7.540517897102072e-12
C45_144 V45 V144 -2.067065703996678e-19

R45_145 V45 V145 -1004.4321243200343
L45_145 V45 V145 -1.3245097510436711e-12
C45_145 V45 V145 -9.561114410026481e-20

R45_146 V45 V146 3403.4773538443796
L45_146 V45 V146 3.868637518370459e-12
C45_146 V45 V146 8.368658157181141e-20

R45_147 V45 V147 -4556.795590678202
L45_147 V45 V147 -3.831430101651787e-12
C45_147 V45 V147 -2.786801638830067e-19

R45_148 V45 V148 -768.446818694748
L45_148 V45 V148 -1.5251338998476215e-12
C45_148 V45 V148 -2.5469251655745998e-19

R45_149 V45 V149 341.6497886821553
L45_149 V45 V149 6.295451632743783e-13
C45_149 V45 V149 6.069289942555585e-19

R45_150 V45 V150 -723.6903820598914
L45_150 V45 V150 -1.9306363402543865e-12
C45_150 V45 V150 -3.2085366268316257e-19

R45_151 V45 V151 -1252.0706706101864
L45_151 V45 V151 -2.5976108305956353e-12
C45_151 V45 V151 9.784071285644203e-20

R45_152 V45 V152 1619.5145088184256
L45_152 V45 V152 5.004338455294693e-12
C45_152 V45 V152 1.2485491386031802e-19

R45_153 V45 V153 -421.8131270167914
L45_153 V45 V153 2.213901698917815e-12
C45_153 V45 V153 2.1738305298438775e-19

R45_154 V45 V154 3169.909030145657
L45_154 V45 V154 5.2766311420476526e-12
C45_154 V45 V154 2.3675850772351574e-19

R45_155 V45 V155 627.0199684790994
L45_155 V45 V155 1.6912637812747219e-12
C45_155 V45 V155 1.7099049555395092e-19

R45_156 V45 V156 -3143.955466240136
L45_156 V45 V156 7.732233637076363e-12
C45_156 V45 V156 2.5238128764401533e-19

R45_157 V45 V157 -558.0241923335203
L45_157 V45 V157 -7.570003355935869e-13
C45_157 V45 V157 -4.2237927212358987e-19

R45_158 V45 V158 1977.091202324195
L45_158 V45 V158 2.3813048880184766e-12
C45_158 V45 V158 6.050517576720482e-20

R45_159 V45 V159 -1779.6574262543074
L45_159 V45 V159 2.443016394541632e-12
C45_159 V45 V159 7.279143973515048e-20

R45_160 V45 V160 1798.9081660733384
L45_160 V45 V160 1.631198168025739e-12
C45_160 V45 V160 -1.0736400654832935e-20

R45_161 V45 V161 -2672.9868387061492
L45_161 V45 V161 4.8740447853579456e-12
C45_161 V45 V161 -1.8463029343418472e-19

R45_162 V45 V162 3106.8659834059117
L45_162 V45 V162 2.111004614816166e-12
C45_162 V45 V162 1.3639359453384843e-19

R45_163 V45 V163 1219.0992401552985
L45_163 V45 V163 4.616208931014469e-12
C45_163 V45 V163 1.2934849808924115e-20

R45_164 V45 V164 26658.635007602366
L45_164 V45 V164 -1.1210933311167993e-11
C45_164 V45 V164 2.789758420763054e-20

R45_165 V45 V165 -979.6486165798772
L45_165 V45 V165 -8.600077216550622e-13
C45_165 V45 V165 -8.711262129140383e-20

R45_166 V45 V166 5022.9247928766
L45_166 V45 V166 -9.788767215981275e-13
C45_166 V45 V166 -2.6899555707491807e-19

R45_167 V45 V167 -4682.715385144182
L45_167 V45 V167 -1.8166293676372358e-12
C45_167 V45 V167 -1.1113225118728261e-19

R45_168 V45 V168 974.2996161699896
L45_168 V45 V168 -1.84384610191515e-12
C45_168 V45 V168 -2.6015042317279635e-19

R45_169 V45 V169 -5334.3742190019475
L45_169 V45 V169 9.895602989608895e-13
C45_169 V45 V169 3.0695997386764868e-19

R45_170 V45 V170 -928.7214782912354
L45_170 V45 V170 3.4133862324011817e-12
C45_170 V45 V170 1.4006113116360224e-19

R45_171 V45 V171 -1259.3263328976489
L45_171 V45 V171 8.786366291619188e-12
C45_171 V45 V171 4.996295633911248e-20

R45_172 V45 V172 -1332.2648885947124
L45_172 V45 V172 1.882399877934347e-11
C45_172 V45 V172 1.3490496891996414e-19

R45_173 V45 V173 -1064.9158539483851
L45_173 V45 V173 1.2065639064259555e-12
C45_173 V45 V173 3.4549734513577726e-20

R45_174 V45 V174 838.5348345837142
L45_174 V45 V174 9.373056064823641e-13
C45_174 V45 V174 1.2368537966345344e-19

R45_175 V45 V175 1125.7794615551882
L45_175 V45 V175 1.2358442687775962e-12
C45_175 V45 V175 2.7793117144853146e-19

R45_176 V45 V176 1651.1329690455232
L45_176 V45 V176 9.112623756828776e-13
C45_176 V45 V176 3.7136935866723876e-19

R45_177 V45 V177 2880.673449958834
L45_177 V45 V177 -7.27553634978197e-13
C45_177 V45 V177 -1.823483640555552e-19

R45_178 V45 V178 -1874.1672873313178
L45_178 V45 V178 -2.189351844657033e-12
C45_178 V45 V178 -1.0642749446601413e-19

R45_179 V45 V179 7143.472760112281
L45_179 V45 V179 -2.1295429076418894e-12
C45_179 V45 V179 -2.4361411853806317e-19

R45_180 V45 V180 -3106.188082796024
L45_180 V45 V180 -1.5177888954366244e-12
C45_180 V45 V180 -3.1556237080417365e-19

R45_181 V45 V181 1287.2395603098273
L45_181 V45 V181 4.8568340501665205e-12
C45_181 V45 V181 -2.710561040100627e-19

R45_182 V45 V182 -2956.23192148968
L45_182 V45 V182 -7.187903835441969e-12
C45_182 V45 V182 7.122823427578482e-20

R45_183 V45 V183 -1871.8153894890231
L45_183 V45 V183 -2.9794210201220913e-12
C45_183 V45 V183 -4.960678566584264e-20

R45_184 V45 V184 -3493.73118085774
L45_184 V45 V184 -1.8208001552923995e-12
C45_184 V45 V184 -3.487381278055423e-20

R45_185 V45 V185 -409.17388329571656
L45_185 V45 V185 2.369177186677355e-12
C45_185 V45 V185 2.9396624177475654e-19

R45_186 V45 V186 791.4519683064835
L45_186 V45 V186 -1.3794250791840489e-12
C45_186 V45 V186 -1.9552502508176466e-19

R45_187 V45 V187 2643.815258370754
L45_187 V45 V187 1.0593470382639178e-11
C45_187 V45 V187 1.6613485493346774e-19

R45_188 V45 V188 1691.3264964773828
L45_188 V45 V188 2.3165877639012507e-12
C45_188 V45 V188 7.81649047196147e-20

R45_189 V45 V189 395.79078932259034
L45_189 V45 V189 2.2502118970680574e-12
C45_189 V45 V189 8.731387766986105e-20

R45_190 V45 V190 -2468.33992628836
L45_190 V45 V190 2.9347073962412253e-12
C45_190 V45 V190 -7.370055813897506e-20

R45_191 V45 V191 -1204.457960791496
L45_191 V45 V191 1.9305448552565825e-12
C45_191 V45 V191 3.1740469706243647e-20

R45_192 V45 V192 -1345.1265199884015
L45_192 V45 V192 2.160778838323442e-12
C45_192 V45 V192 1.1141664861892225e-19

R45_193 V45 V193 1280.2197642244578
L45_193 V45 V193 -7.047102888233721e-12
C45_193 V45 V193 2.3887523446726308e-20

R45_194 V45 V194 -864.331279155844
L45_194 V45 V194 9.193486093712684e-13
C45_194 V45 V194 1.3693228989107268e-19

R45_195 V45 V195 -7085.696002380766
L45_195 V45 V195 -2.942774458316195e-12
C45_195 V45 V195 -1.5542873062240958e-19

R45_196 V45 V196 -2605.368420122345
L45_196 V45 V196 5.635734458715048e-12
C45_196 V45 V196 2.5195482410425918e-20

R45_197 V45 V197 -487.3957451247916
L45_197 V45 V197 -2.0110782995625957e-12
C45_197 V45 V197 -2.375098744965572e-19

R45_198 V45 V198 1136.5018464133432
L45_198 V45 V198 -1.4905920277274465e-12
C45_198 V45 V198 -3.4475321396022145e-20

R45_199 V45 V199 737.3794411049861
L45_199 V45 V199 -2.004507580937076e-12
C45_199 V45 V199 5.627099116777505e-20

R45_200 V45 V200 671.7365879970248
L45_200 V45 V200 -1.1344080731667954e-12
C45_200 V45 V200 -1.2905079394945085e-19

R46_46 V46 0 211.2407632145545
L46_46 V46 0 2.6956515589562814e-13
C46_46 V46 0 2.8939678643804514e-18

R46_47 V46 V47 -4742.536669091243
L46_47 V46 V47 -2.244437288484958e-12
C46_47 V46 V47 -1.3995773956195827e-19

R46_48 V46 V48 -2610.6064331736047
L46_48 V46 V48 -1.5197983124624962e-12
C46_48 V46 V48 -2.1294128356299276e-19

R46_49 V46 V49 9912.171522527153
L46_49 V46 V49 2.3770512494791813e-11
C46_49 V46 V49 -7.284280950410291e-20

R46_50 V46 V50 -4241.903271211827
L46_50 V46 V50 3.1904655985520475e-12
C46_50 V46 V50 1.3047767809513178e-19

R46_51 V46 V51 -28262.503250462356
L46_51 V46 V51 -1.2222802896325594e-11
C46_51 V46 V51 -7.097208734082008e-20

R46_52 V46 V52 20648.339361276423
L46_52 V46 V52 -9.468115932987173e-12
C46_52 V46 V52 -4.414875392890132e-20

R46_53 V46 V53 15161.536499503489
L46_53 V46 V53 7.345900791366052e-12
C46_53 V46 V53 6.187677486735324e-20

R46_54 V46 V54 1823.1780369701382
L46_54 V46 V54 3.355250439199947e-13
C46_54 V46 V54 1.6548425002890606e-18

R46_55 V46 V55 5660.767121949929
L46_55 V46 V55 2.4472419737549703e-12
C46_55 V46 V55 2.1764453227210997e-19

R46_56 V46 V56 2263.500493525987
L46_56 V46 V56 1.291386672206886e-12
C46_56 V46 V56 4.296860058713097e-19

R46_57 V46 V57 14033.812449508026
L46_57 V46 V57 2.67583256857541e-12
C46_57 V46 V57 1.0399370363420059e-19

R46_58 V46 V58 -3204.338916920895
L46_58 V46 V58 -8.788024934462867e-13
C46_58 V46 V58 -7.335195204699469e-19

R46_59 V46 V59 -35029.64328068238
L46_59 V46 V59 -6.038122441163245e-12
C46_59 V46 V59 -1.4886676574208427e-19

R46_60 V46 V60 68388.41246604639
L46_60 V46 V60 -5.181048264670449e-12
C46_60 V46 V60 -1.4354312304641046e-19

R46_61 V46 V61 -6375.645200266278
L46_61 V46 V61 -2.390607950330174e-12
C46_61 V46 V61 -2.1426660167726456e-19

R46_62 V46 V62 2954.4825585496806
L46_62 V46 V62 -6.83402118500661e-13
C46_62 V46 V62 -9.116945795707374e-19

R46_63 V46 V63 -25555.93049873349
L46_63 V46 V63 3.2764099499248387e-11
C46_63 V46 V63 -1.5036873852053282e-20

R46_64 V46 V64 -4893.779626594538
L46_64 V46 V64 -3.213340238463389e-12
C46_64 V46 V64 -1.5611134666432786e-19

R46_65 V46 V65 -7752.941342918614
L46_65 V46 V65 -3.175726082006989e-12
C46_65 V46 V65 -1.891797035243718e-19

R46_66 V46 V66 -2663.2292397507617
L46_66 V46 V66 1.6283299695456138e-12
C46_66 V46 V66 3.399733848976908e-19

R46_67 V46 V67 25447.143851105917
L46_67 V46 V67 3.940686149228244e-12
C46_67 V46 V67 1.8127033351514382e-19

R46_68 V46 V68 -10861.020147919457
L46_68 V46 V68 -6.034371614545532e-11
C46_68 V46 V68 8.062111526265646e-20

R46_69 V46 V69 3325.0860945287895
L46_69 V46 V69 1.4280848375541842e-12
C46_69 V46 V69 4.116564848873302e-19

R46_70 V46 V70 -2142.979613375549
L46_70 V46 V70 1.29245328682221e-12
C46_70 V46 V70 5.171729673798333e-19

R46_71 V46 V71 -8037.4339135300725
L46_71 V46 V71 -2.4691760838336144e-12
C46_71 V46 V71 -1.9846375589971886e-19

R46_72 V46 V72 -13024.20685533349
L46_72 V46 V72 -1.4852051028629904e-11
C46_72 V46 V72 -1.3995660950629223e-20

R46_73 V46 V73 -3423.9315776681124
L46_73 V46 V73 -5.375313992773307e-12
C46_73 V46 V73 -1.650122772267782e-19

R46_74 V46 V74 1996.0431412724174
L46_74 V46 V74 -7.744511647888155e-11
C46_74 V46 V74 -2.1641678463358153e-19

R46_75 V46 V75 -9116.133278839347
L46_75 V46 V75 1.5917743909444834e-11
C46_75 V46 V75 -2.3753894698291394e-20

R46_76 V46 V76 3788.5333201567287
L46_76 V46 V76 1.5332692711715763e-12
C46_76 V46 V76 2.475280942891249e-19

R46_77 V46 V77 25622.92836860006
L46_77 V46 V77 4.005054463585115e-11
C46_77 V46 V77 -1.0792529807090346e-19

R46_78 V46 V78 3339.510597608755
L46_78 V46 V78 -1.646113525286254e-12
C46_78 V46 V78 -1.5403200382311566e-19

R46_79 V46 V79 3054.409418056419
L46_79 V46 V79 4.3326863217861635e-12
C46_79 V46 V79 9.654606466128022e-20

R46_80 V46 V80 8401.232831777483
L46_80 V46 V80 -2.4960970540725165e-12
C46_80 V46 V80 -1.8213109178150235e-19

R46_81 V46 V81 -26830.280656120976
L46_81 V46 V81 -3.4646508670137617e-12
C46_81 V46 V81 -1.1615778688733663e-19

R46_82 V46 V82 -2150.1367127680874
L46_82 V46 V82 -1.1223176568588433e-11
C46_82 V46 V82 -2.0230378936278374e-19

R46_83 V46 V83 -12680.899326006649
L46_83 V46 V83 -9.760891046319967e-12
C46_83 V46 V83 -2.9971301938864056e-20

R46_84 V46 V84 -4451.121902154452
L46_84 V46 V84 -1.617191755946695e-12
C46_84 V46 V84 -2.0595512652129698e-19

R46_85 V46 V85 18674.766244887163
L46_85 V46 V85 -3.6266779460679247e-12
C46_85 V46 V85 -1.453021082679105e-19

R46_86 V46 V86 -817.8482064447819
L46_86 V46 V86 5.934688294553131e-12
C46_86 V46 V86 7.170732107552845e-20

R46_87 V46 V87 -31482.356192409734
L46_87 V46 V87 3.5125159486917898e-12
C46_87 V46 V87 1.9772820849156057e-19

R46_88 V46 V88 26387.03894762001
L46_88 V46 V88 1.5208921306025506e-12
C46_88 V46 V88 3.6148143348583224e-19

R46_89 V46 V89 17689.700706733773
L46_89 V46 V89 1.3345877374129455e-12
C46_89 V46 V89 4.223006652449379e-19

R46_90 V46 V90 622.8678862675253
L46_90 V46 V90 9.034701167989893e-13
C46_90 V46 V90 6.11072905328132e-19

R46_91 V46 V91 -5915.122601669461
L46_91 V46 V91 -1.1310759574269483e-12
C46_91 V46 V91 -4.1091035747503745e-19

R46_92 V46 V92 -7478.16334160392
L46_92 V46 V92 -1.834666007191122e-12
C46_92 V46 V92 -1.806034650236565e-19

R46_93 V46 V93 -21611.423411299926
L46_93 V46 V93 8.909813220587852e-11
C46_93 V46 V93 -4.160043090654418e-20

R46_94 V46 V94 4016.448588504326
L46_94 V46 V94 -1.3794286992738032e-12
C46_94 V46 V94 -4.303259295859897e-19

R46_95 V46 V95 37693.54429488098
L46_95 V46 V95 -1.7871524417374266e-11
C46_95 V46 V95 -1.482626262065812e-19

R46_96 V46 V96 5018.109192629546
L46_96 V46 V96 -2.003610900543433e-11
C46_96 V46 V96 -2.344710676347584e-19

R46_97 V46 V97 5744.030098634774
L46_97 V46 V97 -1.142528821209565e-12
C46_97 V46 V97 -6.433187349769216e-19

R46_98 V46 V98 -760.0654689389172
L46_98 V46 V98 -2.1222530944003168e-12
C46_98 V46 V98 -2.6819497729196985e-19

R46_99 V46 V99 1472.759733211756
L46_99 V46 V99 8.694451125782997e-13
C46_99 V46 V99 6.19127404644373e-19

R46_100 V46 V100 2108.440202053254
L46_100 V46 V100 3.790047279828982e-12
C46_100 V46 V100 3.311891955853786e-19

R46_101 V46 V101 -132225.56585776634
L46_101 V46 V101 1.9034456548175514e-12
C46_101 V46 V101 3.478990277294265e-19

R46_102 V46 V102 1069.9850528258096
L46_102 V46 V102 1.3428013729097252e-12
C46_102 V46 V102 3.307931968390986e-19

R46_103 V46 V103 -1620.1223873599824
L46_103 V46 V103 -1.1609367286159288e-11
C46_103 V46 V103 2.938352703565601e-20

R46_104 V46 V104 -1280.6312356100714
L46_104 V46 V104 -1.0887256315015206e-11
C46_104 V46 V104 5.41008262195346e-20

R46_105 V46 V105 -4151.927834220409
L46_105 V46 V105 1.5242034610754854e-12
C46_105 V46 V105 3.132928628191456e-19

R46_106 V46 V106 -628.2853818026456
L46_106 V46 V106 -1.1152311395917435e-10
C46_106 V46 V106 1.7221675361630666e-19

R46_107 V46 V107 -6666.872719353489
L46_107 V46 V107 -1.0853970886989003e-12
C46_107 V46 V107 -5.343953190754791e-19

R46_108 V46 V108 19331.267205133005
L46_108 V46 V108 1.0567278874223663e-11
C46_108 V46 V108 -1.0329843993726259e-19

R46_109 V46 V109 3201.0239324278396
L46_109 V46 V109 -1.5629694990037012e-12
C46_109 V46 V109 -4.93410753327158e-19

R46_110 V46 V110 736.2501172334867
L46_110 V46 V110 -4.689672788746621e-12
C46_110 V46 V110 -1.7385568724355656e-19

R46_111 V46 V111 5264.343901277517
L46_111 V46 V111 -2.834610821792832e-12
C46_111 V46 V111 -5.805282938197591e-20

R46_112 V46 V112 3270.9476211963492
L46_112 V46 V112 -1.5794232528596747e-12
C46_112 V46 V112 -2.0010817474176697e-19

R46_113 V46 V113 12433.878922576212
L46_113 V46 V113 -1.5664952617185812e-12
C46_113 V46 V113 -2.402139314765068e-19

R46_114 V46 V114 835.7170933383768
L46_114 V46 V114 -2.4346191283033667e-12
C46_114 V46 V114 -3.298921888156936e-19

R46_115 V46 V115 2640.5711145712125
L46_115 V46 V115 8.145248550713783e-13
C46_115 V46 V115 4.76442388827411e-19

R46_116 V46 V116 4140.7359885136975
L46_116 V46 V116 1.7878246643087324e-12
C46_116 V46 V116 1.6203620008796005e-19

R46_117 V46 V117 7118.641038616476
L46_117 V46 V117 1.4720050023112632e-12
C46_117 V46 V117 3.5374073997931927e-19

R46_118 V46 V118 -334.41650309867714
L46_118 V46 V118 1.2838954747468793e-12
C46_118 V46 V118 4.751356890724453e-19

R46_119 V46 V119 -1499.9512353928312
L46_119 V46 V119 2.7688685384217908e-11
C46_119 V46 V119 5.728438468745856e-20

R46_120 V46 V120 -1481.7453322971676
L46_120 V46 V120 2.2647880554732293e-12
C46_120 V46 V120 3.0242276236189377e-19

R46_121 V46 V121 -3869.0371410723014
L46_121 V46 V121 1.6117472747919963e-12
C46_121 V46 V121 1.2421042432693514e-19

R46_122 V46 V122 2273.6354548783615
L46_122 V46 V122 -1.5658489051497234e-12
C46_122 V46 V122 -2.430402061537987e-19

R46_123 V46 V123 -5695.061238359589
L46_123 V46 V123 -1.1458279285838458e-12
C46_123 V46 V123 -3.2928186951876764e-19

R46_124 V46 V124 -11626.352311274388
L46_124 V46 V124 -9.015326253233954e-13
C46_124 V46 V124 -4.853037082862326e-19

R46_125 V46 V125 -1439.2871965582133
L46_125 V46 V125 -2.1330269648105074e-12
C46_125 V46 V125 -1.334163019399879e-19

R46_126 V46 V126 446.3609340864333
L46_126 V46 V126 -1.4475449325614273e-12
C46_126 V46 V126 -1.7338216013778977e-19

R46_127 V46 V127 856.7302652196357
L46_127 V46 V127 -1.1631332987325412e-11
C46_127 V46 V127 -1.0033225490811716e-19

R46_128 V46 V128 826.8480513251552
L46_128 V46 V128 -2.00645437038204e-11
C46_128 V46 V128 -1.1650765559528063e-19

R46_129 V46 V129 901.2566692259554
L46_129 V46 V129 -9.596880683923936e-13
C46_129 V46 V129 -5.715387032921219e-19

R46_130 V46 V130 -993.6555263943454
L46_130 V46 V130 9.05860666087302e-13
C46_130 V46 V130 4.39442533956017e-19

R46_131 V46 V131 -804.9758708788908
L46_131 V46 V131 2.0848867733189608e-12
C46_131 V46 V131 2.66422766426179e-19

R46_132 V46 V132 -619.8721318469046
L46_132 V46 V132 9.816393945708444e-13
C46_132 V46 V132 5.515169657537777e-19

R46_133 V46 V133 3095.4350802482063
L46_133 V46 V133 9.11802552761778e-13
C46_133 V46 V133 5.75127976614629e-19

R46_134 V46 V134 -601.1779238806307
L46_134 V46 V134 -1.4957592843229114e-12
C46_134 V46 V134 -5.174988078265592e-19

R46_135 V46 V135 -1868.5748516636797
L46_135 V46 V135 -2.1873110491124375e-11
C46_135 V46 V135 -4.8800194605234483e-20

R46_136 V46 V136 -961.123021536637
L46_136 V46 V136 -2.6333619786954338e-12
C46_136 V46 V136 -3.22430486166855e-19

R46_137 V46 V137 -666.5586033629916
L46_137 V46 V137 1.3805851235526035e-12
C46_137 V46 V137 4.0395310823607386e-19

R46_138 V46 V138 634.6889065945519
L46_138 V46 V138 -6.757574636303093e-12
C46_138 V46 V138 1.4986206061437828e-19

R46_139 V46 V139 629.303467481229
L46_139 V46 V139 3.5592966462906e-12
C46_139 V46 V139 1.9685123495745132e-19

R46_140 V46 V140 492.70313754181626
L46_140 V46 V140 -2.5469280694910712e-11
C46_140 V46 V140 2.583658751577359e-19

R46_141 V46 V141 -2163.087580167536
L46_141 V46 V141 -6.358332022166558e-13
C46_141 V46 V141 -9.801669179000693e-19

R46_142 V46 V142 429.78908687603194
L46_142 V46 V142 1.862473628374623e-12
C46_142 V46 V142 2.1329672926789414e-19

R46_143 V46 V143 -1334.0766503626023
L46_143 V46 V143 -1.7589330200638241e-12
C46_143 V46 V143 -3.1990893717233715e-19

R46_144 V46 V144 7681.118589254473
L46_144 V46 V144 9.411280819500942e-12
C46_144 V46 V144 -1.413266123077926e-19

R46_145 V46 V145 645.1397740031052
L46_145 V46 V145 -1.348696406334882e-12
C46_145 V46 V145 -3.257354284872692e-19

R46_146 V46 V146 -274.8316231829866
L46_146 V46 V146 -1.2339403983488725e-12
C46_146 V46 V146 -3.395666912274429e-20

R46_147 V46 V147 4442.106203992963
L46_147 V46 V147 -2.3909708085378383e-12
C46_147 V46 V147 -1.9571619467196447e-19

R46_148 V46 V148 -577.7940440882096
L46_148 V46 V148 -9.758192884424142e-13
C46_148 V46 V148 -2.5270951170866654e-19

R46_149 V46 V149 2422.4192784421434
L46_149 V46 V149 3.5772681263516775e-13
C46_149 V46 V149 1.4256039442579355e-18

R46_150 V46 V150 -587.0953150899418
L46_150 V46 V150 1.8762886875753146e-12
C46_150 V46 V150 -8.147239383086569e-19

R46_151 V46 V151 -33341.10773284244
L46_151 V46 V151 7.256233672524627e-12
C46_151 V46 V151 2.660182489826048e-19

R46_152 V46 V152 465.08116056430015
L46_152 V46 V152 8.367222366647225e-12
C46_152 V46 V152 4.8308198235549404e-20

R46_153 V46 V153 -724.3488719922289
L46_153 V46 V153 2.2378603305462005e-12
C46_153 V46 V153 1.19683537367423e-19

R46_154 V46 V154 519.8286114660174
L46_154 V46 V154 1.6355678011850542e-12
C46_154 V46 V154 5.876904295544115e-19

R46_155 V46 V155 688.3668992194008
L46_155 V46 V155 9.31317543916937e-13
C46_155 V46 V155 3.1507446604095344e-19

R46_156 V46 V156 -398.55876580564313
L46_156 V46 V156 2.5963645019425915e-12
C46_156 V46 V156 3.125794390767909e-19

R46_157 V46 V157 -1854.5214194777882
L46_157 V46 V157 -4.324199246278184e-13
C46_157 V46 V157 -1.3380087375314574e-18

R46_158 V46 V158 2223.7503112570503
L46_158 V46 V158 -1.6133927002582128e-12
C46_158 V46 V158 4.412305370397856e-20

R46_159 V46 V159 -408.51775492091195
L46_159 V46 V159 -2.3698718529695768e-11
C46_159 V46 V159 -3.6529378915877045e-20

R46_160 V46 V160 -2559.473938445863
L46_160 V46 V160 1.3977721049201713e-12
C46_160 V46 V160 4.098493914519525e-20

R46_161 V46 V161 674.9737924081651
L46_161 V46 V161 -3.400128712792131e-12
C46_161 V46 V161 -2.80881154390934e-20

R46_162 V46 V162 -1398.2858560123855
L46_162 V46 V162 -5.7373029233128834e-12
C46_162 V46 V162 1.0401409405936556e-19

R46_163 V46 V163 770.4717923619871
L46_163 V46 V163 -1.2912718144131777e-12
C46_163 V46 V163 -2.166773148388763e-19

R46_164 V46 V164 841.8239582198765
L46_164 V46 V164 -1.1696591673526563e-12
C46_164 V46 V164 2.226312644616427e-20

R46_165 V46 V165 -1501.5329231367268
L46_165 V46 V165 9.40568506689074e-13
C46_165 V46 V165 6.345818158663474e-19

R46_166 V46 V166 -706.104555345553
L46_166 V46 V166 8.573042066825086e-13
C46_166 V46 V166 -1.8619420711485458e-19

R46_167 V46 V167 -2792.4421106250434
L46_167 V46 V167 -1.722073155451489e-12
C46_167 V46 V167 -6.097719783438838e-20

R46_168 V46 V168 1552.166257685115
L46_168 V46 V168 -1.6636408244677037e-12
C46_168 V46 V168 -2.612712344191503e-19

R46_169 V46 V169 -610.4883307414777
L46_169 V46 V169 1.5565923154181977e-12
C46_169 V46 V169 -1.0364232944399195e-19

R46_170 V46 V170 904.4956594278442
L46_170 V46 V170 3.2731901612061593e-12
C46_170 V46 V170 3.269982130262871e-19

R46_171 V46 V171 -5250.832990741387
L46_171 V46 V171 6.020321613667364e-13
C46_171 V46 V171 4.845740030289834e-19

R46_172 V46 V172 -1076.9246506669335
L46_172 V46 V172 1.1311262065015625e-12
C46_172 V46 V172 3.1744966059786347e-19

R46_173 V46 V173 952.2285749503488
L46_173 V46 V173 -1.0953544415982265e-12
C46_173 V46 V173 -1.9234658987475297e-19

R46_174 V46 V174 953.003047234747
L46_174 V46 V174 -7.798573523883435e-13
C46_174 V46 V174 -3.0232636904672516e-19

R46_175 V46 V175 -20825.963253746875
L46_175 V46 V175 2.1246877591213216e-12
C46_175 V46 V175 1.7765041836943126e-19

R46_176 V46 V176 4585.582746151397
L46_176 V46 V176 1.4191108370294745e-12
C46_176 V46 V176 2.5797790117849754e-19

R46_177 V46 V177 18682.59412848607
L46_177 V46 V177 -2.8503413069993153e-12
C46_177 V46 V177 8.453133794203837e-20

R46_178 V46 V178 -832.125289355288
L46_178 V46 V178 -2.6096701304003805e-12
C46_178 V46 V178 -1.901545521235573e-19

R46_179 V46 V179 2901.8548027602815
L46_179 V46 V179 -6.761956837714538e-13
C46_179 V46 V179 -6.548116562976068e-19

R46_180 V46 V180 -4709.473931255028
L46_180 V46 V180 -6.823305642804889e-13
C46_180 V46 V180 -5.776423578831344e-19

R46_181 V46 V181 -1700.4625773142861
L46_181 V46 V181 2.0722029228025366e-12
C46_181 V46 V181 -1.5906171785247552e-19

R46_182 V46 V182 -48571.37277785298
L46_182 V46 V182 4.831885776408475e-13
C46_182 V46 V182 3.8106160522794717e-19

R46_183 V46 V183 -1387.9210784065692
L46_183 V46 V183 -1.840071240144804e-12
C46_183 V46 V183 -9.706787546518821e-20

R46_184 V46 V184 -3864.9616695004474
L46_184 V46 V184 -3.2632408171802212e-12
C46_184 V46 V184 5.008701384238192e-20

R46_185 V46 V185 1217595.1182806413
L46_185 V46 V185 3.341587483568439e-11
C46_185 V46 V185 7.035242694472263e-20

R46_186 V46 V186 3447.4777362765412
L46_186 V46 V186 -5.8080554161141935e-11
C46_186 V46 V186 -9.112633572749766e-20

R46_187 V46 V187 2054.8251736468824
L46_187 V46 V187 8.671931505481077e-13
C46_187 V46 V187 5.118905354099938e-19

R46_188 V46 V188 646.3018658671115
L46_188 V46 V188 6.087669899014578e-13
C46_188 V46 V188 3.848471374361403e-19

R46_189 V46 V189 89937.83102100564
L46_189 V46 V189 4.406349685554421e-12
C46_189 V46 V189 3.0844924288222675e-19

R46_190 V46 V190 -1856.9797460160714
L46_190 V46 V190 -8.531849503536773e-13
C46_190 V46 V190 -3.7815372655429507e-19

R46_191 V46 V191 2439.9092439771466
L46_191 V46 V191 1.0358845011672338e-12
C46_191 V46 V191 2.4673351521989353e-19

R46_192 V46 V192 -3164.571815519416
L46_192 V46 V192 1.2088867916280992e-11
C46_192 V46 V192 1.1620122344830782e-19

R46_193 V46 V193 1722.6319476296906
L46_193 V46 V193 -4.2644272003553175e-12
C46_193 V46 V193 -2.2318845324983586e-19

R46_194 V46 V194 -4819.144237880401
L46_194 V46 V194 8.217321802740595e-12
C46_194 V46 V194 -6.469108160938952e-20

R46_195 V46 V195 -1146.1566078143019
L46_195 V46 V195 -6.52174962698805e-13
C46_195 V46 V195 -6.031724466763407e-19

R46_196 V46 V196 -863.3133330411874
L46_196 V46 V196 -8.605345088217067e-13
C46_196 V46 V196 -3.893145465249034e-19

R46_197 V46 V197 13770.976851654765
L46_197 V46 V197 -2.2952084250151907e-12
C46_197 V46 V197 -2.481095934038848e-19

R46_198 V46 V198 6623.424103884716
L46_198 V46 V198 9.94651581934899e-13
C46_198 V46 V198 4.2850807471457133e-20

R46_199 V46 V199 -5482.604516276516
L46_199 V46 V199 -3.0181218190282696e-12
C46_199 V46 V199 -2.0970455990465264e-19

R46_200 V46 V200 941.6788515453927
L46_200 V46 V200 -4.989911352063395e-12
C46_200 V46 V200 -7.958854430451441e-20

R47_47 V47 0 394.1930784294639
L47_47 V47 0 4.1182461317019577e-13
C47_47 V47 0 1.4895370462975722e-18

R47_48 V47 V48 -2090.2912844502357
L47_48 V47 V48 -1.7312155844123032e-12
C47_48 V47 V48 -2.112645296167943e-19

R47_49 V47 V49 7509.338328913925
L47_49 V47 V49 -9.644011143856898e-12
C47_49 V47 V49 -9.815564844025912e-20

R47_50 V47 V50 -229858.47224351246
L47_50 V47 V50 -4.6739355094916435e-12
C47_50 V47 V50 -2.4952347608975027e-19

R47_51 V47 V51 -4677.37054989032
L47_51 V47 V51 9.549313668436424e-13
C47_51 V47 V51 8.882594467614408e-19

R47_52 V47 V52 13884.433886229956
L47_52 V47 V52 -1.5191832183629665e-11
C47_52 V47 V52 3.02027992166925e-22

R47_53 V47 V53 -25623.06775864622
L47_53 V47 V53 2.1235774026343207e-11
C47_53 V47 V53 3.898827292842591e-20

R47_54 V47 V54 15281.685105836248
L47_54 V47 V54 4.754417199508877e-12
C47_54 V47 V54 1.0498590927987702e-19

R47_55 V47 V55 2527.7886189867563
L47_55 V47 V55 5.204622342266604e-13
C47_55 V47 V55 9.937738224468129e-19

R47_56 V47 V56 2921.2258022319243
L47_56 V47 V56 2.3387623242117875e-12
C47_56 V47 V56 2.0906670554461157e-19

R47_57 V47 V57 7816.428421955226
L47_57 V47 V57 3.157197778349427e-12
C47_57 V47 V57 9.534652833278421e-20

R47_58 V47 V58 -3642.4194783410667
L47_58 V47 V58 3.54909886912932e-12
C47_58 V47 V58 1.6517397496558175e-19

R47_59 V47 V59 3193.122435685885
L47_59 V47 V59 -6.06997452937192e-13
C47_59 V47 V59 -1.221647138919686e-18

R47_60 V47 V60 5627.335190695361
L47_60 V47 V60 -3.983335730376393e-11
C47_60 V47 V60 -7.865457577271184e-20

R47_61 V47 V61 -7066.012021213717
L47_61 V47 V61 -5.121873991956877e-12
C47_61 V47 V61 -7.536702107122525e-20

R47_62 V47 V62 6067.06962196358
L47_62 V47 V62 -3.661011662395645e-12
C47_62 V47 V62 -2.1193566444221894e-19

R47_63 V47 V63 9030.378613379968
L47_63 V47 V63 7.87466058392009e-12
C47_63 V47 V63 2.4932267814900975e-19

R47_64 V47 V64 -6298.431395014797
L47_64 V47 V64 -5.263969306347789e-11
C47_64 V47 V64 3.972166625710944e-20

R47_65 V47 V65 -15475.691318245666
L47_65 V47 V65 -3.849773216936119e-12
C47_65 V47 V65 -1.5728546748739383e-19

R47_66 V47 V66 -14605.61644852728
L47_66 V47 V66 -4.8969944797315465e-12
C47_66 V47 V66 -1.4126424681817503e-19

R47_67 V47 V67 -2449.2955720563245
L47_67 V47 V67 1.4105449078351135e-12
C47_67 V47 V67 5.006310331759964e-19

R47_68 V47 V68 -3966.904728613168
L47_68 V47 V68 -5.808972949292211e-12
C47_68 V47 V68 -3.297962473052791e-20

R47_69 V47 V69 6000.349467464537
L47_69 V47 V69 4.209201724988152e-12
C47_69 V47 V69 1.3148626959502048e-19

R47_70 V47 V70 -26065.401271172286
L47_70 V47 V70 2.645366550696911e-12
C47_70 V47 V70 2.272020027774899e-19

R47_71 V47 V71 -1563.8023067250367
L47_71 V47 V71 -1.3128378265186792e-12
C47_71 V47 V71 -5.484197551103291e-19

R47_72 V47 V72 -4847.364723349766
L47_72 V47 V72 -1.374315182706361e-11
C47_72 V47 V72 -1.8071545837900615e-20

R47_73 V47 V73 -3824.4027746806905
L47_73 V47 V73 -9.620735434042446e-12
C47_73 V47 V73 -3.6333338959671437e-20

R47_74 V47 V74 11271.995790380342
L47_74 V47 V74 2.5253511626359407e-11
C47_74 V47 V74 -3.0146342071967614e-20

R47_75 V47 V75 1904.4657509959907
L47_75 V47 V75 5.127133374737586e-12
C47_75 V47 V75 2.761485090118514e-20

R47_76 V47 V76 2299.0249193570735
L47_76 V47 V76 2.0589496784210506e-12
C47_76 V47 V76 1.618950192982015e-19

R47_77 V47 V77 8271.149173829
L47_77 V47 V77 6.7204194389897255e-12
C47_77 V47 V77 -3.330273870574167e-20

R47_78 V47 V78 -6749.620357347533
L47_78 V47 V78 5.17807408543612e-11
C47_78 V47 V78 2.3826679148739353e-20

R47_79 V47 V79 1041.937933197791
L47_79 V47 V79 -1.3461041804831407e-11
C47_79 V47 V79 1.6299819954366895e-19

R47_80 V47 V80 3568.0561743939897
L47_80 V47 V80 -3.9341988842887585e-12
C47_80 V47 V80 -9.333460420309211e-20

R47_81 V47 V81 5332.140660939684
L47_81 V47 V81 -4.994167188825965e-12
C47_81 V47 V81 -5.0268454731490656e-20

R47_82 V47 V82 13005.219880177168
L47_82 V47 V82 -3.116162179295006e-12
C47_82 V47 V82 -1.827827403653828e-19

R47_83 V47 V83 -1790.1770536572217
L47_83 V47 V83 2.4071334089964643e-11
C47_83 V47 V83 -2.5610718226453602e-20

R47_84 V47 V84 -3213.821921192672
L47_84 V47 V84 -2.681243709727985e-12
C47_84 V47 V84 -1.0445055890376248e-19

R47_85 V47 V85 -24430.068743327178
L47_85 V47 V85 -3.849980213272936e-12
C47_85 V47 V85 -9.429443341579475e-20

R47_86 V47 V86 -2394.922981159552
L47_86 V47 V86 -7.459421728156359e-12
C47_86 V47 V86 -8.073588441802507e-20

R47_87 V47 V87 -732.1931669274512
L47_87 V47 V87 1.0043953894739129e-12
C47_87 V47 V87 2.3687311379307624e-19

R47_88 V47 V88 -4525.0350923881
L47_88 V47 V88 1.90466737721177e-12
C47_88 V47 V88 2.137191281704316e-19

R47_89 V47 V89 -3941.5802352062246
L47_89 V47 V89 3.604802764221632e-12
C47_89 V47 V89 1.40610690522637e-19

R47_90 V47 V90 28819.8641324173
L47_90 V47 V90 1.117255230067729e-12
C47_90 V47 V90 4.341429757379527e-19

R47_91 V47 V91 765.0421826380436
L47_91 V47 V91 -4.872813112317267e-13
C47_91 V47 V91 -6.582457271919337e-19

R47_92 V47 V92 20603.705331117195
L47_92 V47 V92 -1.6837879860559213e-12
C47_92 V47 V92 -1.693007512782781e-19

R47_93 V47 V93 11376.393600242685
L47_93 V47 V93 2.990016154028188e-12
C47_93 V47 V93 9.521029380834388e-20

R47_94 V47 V94 3217.681118743186
L47_94 V47 V94 -3.128078571597796e-12
C47_94 V47 V94 -2.0843274812662465e-19

R47_95 V47 V95 659.4973254945052
L47_95 V47 V95 -6.79705964476734e-12
C47_95 V47 V95 2.1213902429052135e-20

R47_96 V47 V96 1492.1608368123932
L47_96 V47 V96 -6.611773971308506e-11
C47_96 V47 V96 -9.821898018166411e-20

R47_97 V47 V97 1904.61218056584
L47_97 V47 V97 -1.4651813693692683e-12
C47_97 V47 V97 -3.5358407111292417e-19

R47_98 V47 V98 -2925.5950687457016
L47_98 V47 V98 -1.6162608717675213e-12
C47_98 V47 V98 -2.7686610937741555e-19

R47_99 V47 V99 -374.2583264856022
L47_99 V47 V99 3.9920354033382963e-13
C47_99 V47 V99 8.013071549278294e-19

R47_100 V47 V100 -2827.491403432764
L47_100 V47 V100 2.0951980295291223e-12
C47_100 V47 V100 2.423642879484083e-19

R47_101 V47 V101 -5194.986729877414
L47_101 V47 V101 2.4840724764456876e-11
C47_101 V47 V101 1.1550053270497393e-19

R47_102 V47 V102 436703.3372107776
L47_102 V47 V102 1.6641940652760851e-12
C47_102 V47 V102 3.1985957443553553e-19

R47_103 V47 V103 1386.8925984330729
L47_103 V47 V103 -8.874805291068968e-13
C47_103 V47 V103 -5.824989426995506e-19

R47_104 V47 V104 -2853.609530179283
L47_104 V47 V104 -4.682925852372785e-12
C47_104 V47 V104 -4.8003655800595275e-20

R47_105 V47 V105 -2654.841117306424
L47_105 V47 V105 1.5448064770183632e-12
C47_105 V47 V105 1.5908655777637827e-19

R47_106 V47 V106 -1785.7684943373952
L47_106 V47 V106 1.9065157744959294e-12
C47_106 V47 V106 1.2631391423012135e-19

R47_107 V47 V107 990.605230031091
L47_107 V47 V107 -7.597983711977321e-13
C47_107 V47 V107 -1.5166708858631492e-19

R47_108 V47 V108 6786.9719899981765
L47_108 V47 V108 -1.36445305395881e-11
C47_108 V47 V108 -8.597420478387268e-20

R47_109 V47 V109 101205.51843630002
L47_109 V47 V109 -3.536782224393683e-12
C47_109 V47 V109 -2.4930880009551604e-19

R47_110 V47 V110 2392.4930030078103
L47_110 V47 V110 -1.548952157327552e-12
C47_110 V47 V110 -1.9686497113714105e-19

R47_111 V47 V111 -405.472044160907
L47_111 V47 V111 1.2709601383115617e-12
C47_111 V47 V111 2.6729398160159847e-19

R47_112 V47 V112 -1819.3609256029918
L47_112 V47 V112 -4.8363805579965714e-12
C47_112 V47 V112 -8.839425488921374e-20

R47_113 V47 V113 1593.4806371976867
L47_113 V47 V113 -1.3041368198999643e-12
C47_113 V47 V113 -4.051076106456184e-20

R47_114 V47 V114 1607.9896927834418
L47_114 V47 V114 -1.9372582444435475e-12
C47_114 V47 V114 -1.6465805326917434e-19

R47_115 V47 V115 708.4737502533488
L47_115 V47 V115 9.127225534359389e-13
C47_115 V47 V115 2.7070100718669736e-20

R47_116 V47 V116 1294.0099363224222
L47_116 V47 V116 2.4248149695044936e-12
C47_116 V47 V116 1.1688578573388956e-19

R47_117 V47 V117 2414.166046528514
L47_117 V47 V117 2.6309750959159877e-12
C47_117 V47 V117 1.6761627601790366e-19

R47_118 V47 V118 -1164.0453292381144
L47_118 V47 V118 1.0430518532841622e-12
C47_118 V47 V118 3.691761528558123e-19

R47_119 V47 V119 84101.70965116977
L47_119 V47 V119 -8.144811264614704e-13
C47_119 V47 V119 1.4337078841734704e-20

R47_120 V47 V120 -2638.864435939412
L47_120 V47 V120 6.871548243374728e-12
C47_120 V47 V120 1.7810992525352446e-19

R47_121 V47 V121 -1933.7561939063742
L47_121 V47 V121 1.8218366403602503e-12
C47_121 V47 V121 -6.299012722456219e-20

R47_122 V47 V122 -6130.354555812298
L47_122 V47 V122 -5.715242989586395e-12
C47_122 V47 V122 -1.2182718157799768e-19

R47_123 V47 V123 -679.8332870326705
L47_123 V47 V123 1.1904496818298129e-11
C47_123 V47 V123 -1.5101068768809223e-19

R47_124 V47 V124 -1366.1303699395626
L47_124 V47 V124 -1.5729880233998306e-12
C47_124 V47 V124 -3.413818110416385e-19

R47_125 V47 V125 -1168.220859444539
L47_125 V47 V125 -5.481632685798545e-12
C47_125 V47 V125 -3.7112063185746015e-20

R47_126 V47 V126 5720.4813039188775
L47_126 V47 V126 -1.072081002991468e-12
C47_126 V47 V126 -2.490859417183111e-19

R47_127 V47 V127 807.082877641047
L47_127 V47 V127 1.214863029944753e-12
C47_127 V47 V127 5.127165774277093e-20

R47_128 V47 V128 1464.42921200564
L47_128 V47 V128 1.728498105508271e-11
C47_128 V47 V128 -7.011995779750505e-20

R47_129 V47 V129 838.4889605513353
L47_129 V47 V129 -1.2588182616442868e-12
C47_129 V47 V129 -2.191017275952439e-19

R47_130 V47 V130 1522.208762929895
L47_130 V47 V130 1.326736317801498e-12
C47_130 V47 V130 2.790190570474712e-19

R47_131 V47 V131 -1627.2195793099213
L47_131 V47 V131 -1.329086149609861e-12
C47_131 V47 V131 8.301797834991752e-20

R47_132 V47 V132 -4493.031711240586
L47_132 V47 V132 2.4193919585551944e-12
C47_132 V47 V132 3.9178016154908186e-19

R47_133 V47 V133 1327.6295466369904
L47_133 V47 V133 2.838489298913375e-12
C47_133 V47 V133 2.7143165560127747e-19

R47_134 V47 V134 -5209.3371238036525
L47_134 V47 V134 -3.64308263862817e-12
C47_134 V47 V134 -8.841285106440131e-20

R47_135 V47 V135 -905.2638827780979
L47_135 V47 V135 2.7044328528947077e-12
C47_135 V47 V135 -2.5767052136445363e-19

R47_136 V47 V136 -1861.0370765397256
L47_136 V47 V136 -3.606497313476552e-12
C47_136 V47 V136 -2.197699438855556e-19

R47_137 V47 V137 -820.3873224281542
L47_137 V47 V137 1.1549237734951972e-12
C47_137 V47 V137 1.5943276441455078e-19

R47_138 V47 V138 13872.993412675401
L47_138 V47 V138 -5.436618615788318e-12
C47_138 V47 V138 -7.392751612180983e-20

R47_139 V47 V139 465.8834642436077
L47_139 V47 V139 1.8136403472568775e-11
C47_139 V47 V139 4.2205677615345984e-19

R47_140 V47 V140 1025.1179874481113
L47_140 V47 V140 7.946630894568423e-12
C47_140 V47 V140 1.8952528869758917e-19

R47_141 V47 V141 -891.9505903628448
L47_141 V47 V141 -1.4127337899527979e-12
C47_141 V47 V141 -4.921172943514351e-19

R47_142 V47 V142 7672.749531051621
L47_142 V47 V142 3.4254779197401096e-12
C47_142 V47 V142 8.479958016207273e-21

R47_143 V47 V143 -978.0464678799628
L47_143 V47 V143 -8.839055348235441e-13
C47_143 V47 V143 -1.7238224216651048e-19

R47_144 V47 V144 -4202.652169132992
L47_144 V47 V144 -1.015504010738801e-11
C47_144 V47 V144 -7.994451082162543e-20

R47_145 V47 V145 615.5429439937633
L47_145 V47 V145 -9.203576608249687e-13
C47_145 V47 V145 -1.5465628966718348e-19

R47_146 V47 V146 -7952.877323191766
L47_146 V47 V146 -3.0810176933083843e-12
C47_146 V47 V146 8.901732997768265e-20

R47_147 V47 V147 1048.2044034736032
L47_147 V47 V147 1.4924688941459555e-12
C47_147 V47 V147 -3.3855800914382505e-19

R47_148 V47 V148 -9869.681677076227
L47_148 V47 V148 -1.335746841030811e-12
C47_148 V47 V148 -1.8256069489153173e-19

R47_149 V47 V149 2794.6625905470096
L47_149 V47 V149 6.515016449216606e-13
C47_149 V47 V149 6.5519218561627e-19

R47_150 V47 V150 -810.7728720348096
L47_150 V47 V150 -8.594221603342233e-12
C47_150 V47 V150 -2.8533885780353896e-19

R47_151 V47 V151 -262.31557311666467
L47_151 V47 V151 9.182636616312385e-13
C47_151 V47 V151 1.4039151808297555e-19

R47_152 V47 V152 -2700.1902957701964
L47_152 V47 V152 5.05792515709376e-12
C47_152 V47 V152 3.4956759635517406e-20

R47_153 V47 V153 -2677.055121700467
L47_153 V47 V153 1.935182855197459e-12
C47_153 V47 V153 8.060640272748822e-20

R47_154 V47 V154 5887.58677244416
L47_154 V47 V154 1.8054410803408627e-12
C47_154 V47 V154 1.7861656080699914e-19

R47_155 V47 V155 118.3850218796986
L47_155 V47 V155 4.057272473930124e-12
C47_155 V47 V155 3.723917099311313e-19

R47_156 V47 V156 -2296.773502548753
L47_156 V47 V156 2.975359839087627e-12
C47_156 V47 V156 1.7684393436332625e-19

R47_157 V47 V157 -1771.975309388877
L47_157 V47 V157 -1.4154198034714383e-12
C47_157 V47 V157 -5.569641377220176e-19

R47_158 V47 V158 -7268.571602322918
L47_158 V47 V158 4.583094529927332e-12
C47_158 V47 V158 3.0726106669944844e-20

R47_159 V47 V159 -327.9108536199082
L47_159 V47 V159 -5.806653076640679e-13
C47_159 V47 V159 -1.9037671776683204e-19

R47_160 V47 V160 1572.6842712814307
L47_160 V47 V160 2.533652256858537e-12
C47_160 V47 V160 3.906908511747845e-21

R47_161 V47 V161 3736.8406235698535
L47_161 V47 V161 -6.2768943438373344e-12
C47_161 V47 V161 -7.110533539962945e-21

R47_162 V47 V162 19866.137103348236
L47_162 V47 V162 7.937304591801185e-12
C47_162 V47 V162 9.968088184751622e-20

R47_163 V47 V163 -525.1719609731185
L47_163 V47 V163 5.3940311848430245e-12
C47_163 V47 V163 2.4664091016681276e-20

R47_164 V47 V164 -840.8271005774991
L47_164 V47 V164 -1.9397163340282475e-12
C47_164 V47 V164 4.0939578580745774e-20

R47_165 V47 V165 48948.85432179149
L47_165 V47 V165 -7.009373476246753e-12
C47_165 V47 V165 1.5584722929489427e-19

R47_166 V47 V166 -1636.5118392374554
L47_166 V47 V166 -2.3551583480198194e-12
C47_166 V47 V166 -1.5772426455433087e-19

R47_167 V47 V167 3899.939870220435
L47_167 V47 V167 1.0939322212051058e-12
C47_167 V47 V167 8.067914664260623e-21

R47_168 V47 V168 973.4016561414355
L47_168 V47 V168 -7.011959615926185e-12
C47_168 V47 V168 -1.0847032249944726e-19

R47_169 V47 V169 -1383.7431492586104
L47_169 V47 V169 8.608438703267116e-12
C47_169 V47 V169 -5.963799261917349e-20

R47_170 V47 V170 -5421.569348148988
L47_170 V47 V170 7.035663254899856e-12
C47_170 V47 V170 1.668267915634553e-19

R47_171 V47 V171 380.93771317156546
L47_171 V47 V171 2.8578035178434464e-12
C47_171 V47 V171 7.875232071276127e-20

R47_172 V47 V172 2396.3970897343224
L47_172 V47 V172 5.816669010124337e-12
C47_172 V47 V172 8.74056488664334e-20

R47_173 V47 V173 2420.372826960417
L47_173 V47 V173 2.8029206521775395e-12
C47_173 V47 V173 2.771931161362203e-20

R47_174 V47 V174 800.3855198498917
L47_174 V47 V174 2.0274400479792976e-12
C47_174 V47 V174 -7.928763503805392e-20

R47_175 V47 V175 -451.25052281240806
L47_175 V47 V175 -2.7269237132547094e-12
C47_175 V47 V175 1.6057111988584639e-19

R47_176 V47 V176 -7971.406255340011
L47_176 V47 V176 2.901188903770846e-12
C47_176 V47 V176 1.739948054283238e-19

R47_177 V47 V177 -2251.6328592297227
L47_177 V47 V177 -2.6574332772465056e-12
C47_177 V47 V177 -2.8106297502278147e-20

R47_178 V47 V178 -1101.9221647625359
L47_178 V47 V178 -2.9301033522474583e-12
C47_178 V47 V178 -1.0314010082903987e-19

R47_179 V47 V179 466.4540416430404
L47_179 V47 V179 -1.3196249192305812e-12
C47_179 V47 V179 -2.258563301388205e-19

R47_180 V47 V180 -1971.6576249784355
L47_180 V47 V180 -2.102647343310459e-12
C47_180 V47 V180 -2.653922818595241e-19

R47_181 V47 V181 7178.800339072723
L47_181 V47 V181 8.031389592678983e-12
C47_181 V47 V181 -1.0959011847504517e-19

R47_182 V47 V182 1615.9287783586392
L47_182 V47 V182 3.095225577895022e-12
C47_182 V47 V182 1.2746443002568039e-19

R47_183 V47 V183 -579.81596728909
L47_183 V47 V183 3.239411448220489e-12
C47_183 V47 V183 -5.560626241277819e-20

R47_184 V47 V184 -40905.91687635772
L47_184 V47 V184 -2.9843050299213395e-12
C47_184 V47 V184 1.0572243171660466e-20

R47_185 V47 V185 5998.115699306751
L47_185 V47 V185 8.558782666350366e-12
C47_185 V47 V185 9.743750391133615e-20

R47_186 V47 V186 2398.8664668791384
L47_186 V47 V186 -3.7379679382968965e-12
C47_186 V47 V186 -6.917926495886455e-20

R47_187 V47 V187 -7117.373153982104
L47_187 V47 V187 1.2721268275374255e-12
C47_187 V47 V187 2.3461625013501337e-19

R47_188 V47 V188 705.7330945781713
L47_188 V47 V188 1.1313017660380676e-12
C47_188 V47 V188 1.9970250334965918e-19

R47_189 V47 V189 -1869.5880398547906
L47_189 V47 V189 -6.82886356075659e-11
C47_189 V47 V189 8.515100845054445e-20

R47_190 V47 V190 -1555.4331855231344
L47_190 V47 V190 2.6682756282234484e-11
C47_190 V47 V190 -1.1111904345226407e-19

R47_191 V47 V191 1040.561423045188
L47_191 V47 V191 -4.6188676777213264e-12
C47_191 V47 V191 -1.5755446527829222e-20

R47_192 V47 V192 -3721.614037443522
L47_192 V47 V192 2.3326273805170925e-11
C47_192 V47 V192 -1.7790120557207455e-20

R47_193 V47 V193 2738.376351659823
L47_193 V47 V193 -8.326113658571859e-11
C47_193 V47 V193 -7.82636399420087e-20

R47_194 V47 V194 7078.2819509221345
L47_194 V47 V194 -2.9241630701890876e-10
C47_194 V47 V194 -8.666311720802033e-20

R47_195 V47 V195 -1135.383839121224
L47_195 V47 V195 -3.807761546121916e-12
C47_195 V47 V195 -7.723787592714249e-20

R47_196 V47 V196 -549.0441555632881
L47_196 V47 V196 -1.6336463334635235e-12
C47_196 V47 V196 -1.1922449454239038e-19

R47_197 V47 V197 -6821.989381296605
L47_197 V47 V197 -8.894641217303995e-12
C47_197 V47 V197 -9.011747302148123e-20

R47_198 V47 V198 -2293.48999596569
L47_198 V47 V198 -1.3272098340348694e-11
C47_198 V47 V198 1.8423259250251758e-20

R47_199 V47 V199 -8578.766643050147
L47_199 V47 V199 2.8507364399630187e-12
C47_199 V47 V199 -1.7367656041026932e-20

R47_200 V47 V200 1207.428629001166
L47_200 V47 V200 7.2902626097085e-12
C47_200 V47 V200 2.348843127364256e-20

R48_48 V48 0 132.68995547501856
L48_48 V48 0 1.8603132039842346e-13
C48_48 V48 0 2.9891627716026827e-18

R48_49 V48 V49 7868.557809620061
L48_49 V48 V49 -1.1089333449185006e-11
C48_49 V48 V49 -9.630096339417959e-20

R48_50 V48 V50 27488.60541848
L48_50 V48 V50 -7.522486701879751e-12
C48_50 V48 V50 -2.314868636663932e-19

R48_51 V48 V51 -7971.421176913037
L48_51 V48 V51 -2.563072266632671e-12
C48_51 V48 V51 -2.528729517967512e-19

R48_52 V48 V52 7288.807236652612
L48_52 V48 V52 8.932379870868644e-13
C48_52 V48 V52 9.04969418219179e-19

R48_53 V48 V53 -19539.517719079922
L48_53 V48 V53 1.9306789242879867e-11
C48_53 V48 V53 7.456111186330557e-20

R48_54 V48 V54 4988.899798899357
L48_54 V48 V54 2.584064572306343e-12
C48_54 V48 V54 2.001876323490758e-19

R48_55 V48 V55 12800.668331113078
L48_55 V48 V55 6.761031492307092e-12
C48_55 V48 V55 7.063482825142291e-20

R48_56 V48 V56 920.0957432746782
L48_56 V48 V56 3.830798099621521e-13
C48_56 V48 V56 1.3853373085027124e-18

R48_57 V48 V57 5070.900213120788
L48_57 V48 V57 1.9479948081306135e-12
C48_57 V48 V57 1.502028616787247e-19

R48_58 V48 V58 -2409.1275940261357
L48_58 V48 V58 4.763782805304146e-12
C48_58 V48 V58 1.285473266918851e-19

R48_59 V48 V59 7932.394289195384
L48_59 V48 V59 1.5946510322105577e-11
C48_59 V48 V59 -2.9239763607724423e-20

R48_60 V48 V60 1879.3700057501742
L48_60 V48 V60 -6.209744497577186e-13
C48_60 V48 V60 -1.2634920041284958e-18

R48_61 V48 V61 -5093.937869082993
L48_61 V48 V61 -2.682857477751746e-12
C48_61 V48 V61 -1.66196770245264e-19

R48_62 V48 V62 4432.1517770455475
L48_62 V48 V62 -2.4392916626237357e-12
C48_62 V48 V62 -3.038288777260865e-19

R48_63 V48 V63 -10838.365454867344
L48_63 V48 V63 4.175896469409764e-12
C48_63 V48 V63 8.963326674988782e-20

R48_64 V48 V64 -5413.470257120452
L48_64 V48 V64 -3.5631394643482884e-12
C48_64 V48 V64 1.2285014657079635e-19

R48_65 V48 V65 -4760.18948028553
L48_65 V48 V65 -2.2394781350471104e-12
C48_65 V48 V65 -2.6462296737075223e-19

R48_66 V48 V66 -16668.213773663796
L48_66 V48 V66 -5.202605485622756e-12
C48_66 V48 V66 -1.669577759214334e-19

R48_67 V48 V67 68921.86741969711
L48_67 V48 V67 -1.5199315734228484e-11
C48_67 V48 V67 -3.753971318084862e-20

R48_68 V48 V68 -1452.0004906899828
L48_68 V48 V68 2.240454693774114e-12
C48_68 V48 V68 3.9947427223083426e-19

R48_69 V48 V69 4281.597373504269
L48_69 V48 V69 2.4513116035731518e-12
C48_69 V48 V69 2.561600757941225e-19

R48_70 V48 V70 -13733.897671418874
L48_70 V48 V70 1.907920545815554e-12
C48_70 V48 V70 3.3085491539854016e-19

R48_71 V48 V71 -5534.308098546015
L48_71 V48 V71 -2.7255164915343596e-12
C48_71 V48 V71 -1.0537016582795113e-19

R48_72 V48 V72 -1135.2806949288617
L48_72 V48 V72 -1.916705746367263e-12
C48_72 V48 V72 -4.264798954249679e-19

R48_73 V48 V73 -3407.260927849045
L48_73 V48 V73 -6.727444154894191e-12
C48_73 V48 V73 -6.652039541931492e-20

R48_74 V48 V74 5566.14726279686
L48_74 V48 V74 1.3516445129262576e-11
C48_74 V48 V74 -2.0704871301949455e-20

R48_75 V48 V75 -5839.712061504607
L48_75 V48 V75 1.7646284866881016e-11
C48_75 V48 V75 -5.651140186341745e-20

R48_76 V48 V76 651.5535537022173
L48_76 V48 V76 1.00078447609455e-12
C48_76 V48 V76 3.6246524733742363e-19

R48_77 V48 V77 6281.614662775922
L48_77 V48 V77 4.209898377797315e-12
C48_77 V48 V77 -2.504165642850983e-20

R48_78 V48 V78 -3151.114122965867
L48_78 V48 V78 -1.5985785039835833e-11
C48_78 V48 V78 2.1151741825728055e-21

R48_79 V48 V79 2070.719737139591
L48_79 V48 V79 5.072947259168252e-12
C48_79 V48 V79 6.330921849870351e-20

R48_80 V48 V80 1736.9384837854454
L48_80 V48 V80 -1.2215926801750372e-12
C48_80 V48 V80 -1.3486367642138012e-19

R48_81 V48 V81 -6741.480793874996
L48_81 V48 V81 -2.04522768424622e-12
C48_81 V48 V81 -1.6957266255718607e-19

R48_82 V48 V82 12267.051400307178
L48_82 V48 V82 -2.3925115977929395e-12
C48_82 V48 V82 -2.56592322175967e-19

R48_83 V48 V83 -4608.785177828381
L48_83 V48 V83 -1.1944084119865713e-11
C48_83 V48 V83 -2.2427149724310883e-20

R48_84 V48 V84 -1286.412426019363
L48_84 V48 V84 -2.5003328520955548e-12
C48_84 V48 V84 -1.2245217710064887e-19

R48_85 V48 V85 36548.844366043086
L48_85 V48 V85 -2.7980372943293034e-12
C48_85 V48 V85 -1.3433822553775032e-19

R48_86 V48 V86 -2822.4020333272
L48_86 V48 V86 -6.302216642456769e-12
C48_86 V48 V86 -9.405389843145113e-20

R48_87 V48 V87 -3966.9876138969444
L48_87 V48 V87 2.8488484494969916e-12
C48_87 V48 V87 1.367848060565575e-19

R48_88 V48 V88 -633.207032019592
L48_88 V48 V88 6.950907019848561e-13
C48_88 V48 V88 4.080833743939859e-19

R48_89 V48 V89 -5437.031525267322
L48_89 V48 V89 2.092946111811428e-12
C48_89 V48 V89 2.3539429723157513e-19

R48_90 V48 V90 14581.727661515491
L48_90 V48 V90 8.331272570229631e-13
C48_90 V48 V90 5.701044389190416e-19

R48_91 V48 V91 -2126.7843505543724
L48_91 V48 V91 -9.372038659483886e-13
C48_91 V48 V91 -3.8963769328587135e-19

R48_92 V48 V92 503.87424172339433
L48_92 V48 V92 -4.935195491095047e-13
C48_92 V48 V92 -5.64207514158277e-19

R48_93 V48 V93 -4017.6905866408724
L48_93 V48 V93 2.5444385736506535e-12
C48_93 V48 V93 1.0712781482672615e-19

R48_94 V48 V94 6931.712443627501
L48_94 V48 V94 -2.354971141206045e-12
C48_94 V48 V94 -2.9042980518908037e-19

R48_95 V48 V95 1660.3538032101337
L48_95 V48 V95 4.3363939382422365e-11
C48_95 V48 V95 -6.867654903449896e-20

R48_96 V48 V96 438.3856017813874
L48_96 V48 V96 1.6036822304545746e-11
C48_96 V48 V96 -4.2518792133766636e-20

R48_97 V48 V97 1481.292095101905
L48_97 V48 V97 -1.0620174594169768e-12
C48_97 V48 V97 -4.898646553557842e-19

R48_98 V48 V98 -4211.391293109732
L48_98 V48 V98 -1.1172969532355549e-12
C48_98 V48 V98 -3.915948101607616e-19

R48_99 V48 V99 58622.144225022304
L48_99 V48 V99 8.590661498874264e-13
C48_99 V48 V99 4.3035951694316326e-19

R48_100 V48 V100 -244.5337237754671
L48_100 V48 V100 4.60157304451921e-13
C48_100 V48 V100 8.681802450805164e-19

R48_101 V48 V101 -4259.018353070506
L48_101 V48 V101 8.753851976059835e-12
C48_101 V48 V101 1.2412244146432866e-19

R48_102 V48 V102 7248.35937301686
L48_102 V48 V102 1.2426905689772529e-12
C48_102 V48 V102 4.1573519415301405e-19

R48_103 V48 V103 -1757.9863754984758
L48_103 V48 V103 -4.520871638315447e-12
C48_103 V48 V103 -8.015823519581401e-21

R48_104 V48 V104 1753.3873115695458
L48_104 V48 V104 -8.119790711829328e-13
C48_104 V48 V104 -6.565934704829066e-19

R48_105 V48 V105 -1281.8156390692936
L48_105 V48 V105 1.4201404674718538e-12
C48_105 V48 V105 1.9199276194027377e-19

R48_106 V48 V106 -945.4717195551381
L48_106 V48 V106 1.68639101866093e-12
C48_106 V48 V106 1.6537219386677369e-19

R48_107 V48 V107 -8647.590534743167
L48_107 V48 V107 -1.2238340646546005e-12
C48_107 V48 V107 -3.879604541381857e-19

R48_108 V48 V108 435.83371409889116
L48_108 V48 V108 -1.3288275456532954e-12
C48_108 V48 V108 -1.353191142009773e-21

R48_109 V48 V109 2017.5071733203883
L48_109 V48 V109 -1.8874808128344298e-12
C48_109 V48 V109 -3.592153894551765e-19

R48_110 V48 V110 946.7129085509023
L48_110 V48 V110 -1.434620285491094e-12
C48_110 V48 V110 -2.286715858507496e-19

R48_111 V48 V111 -2053.3936999777156
L48_111 V48 V111 -7.932305866041856e-12
C48_111 V48 V111 7.284041459693768e-22

R48_112 V48 V112 -365.2945687179777
L48_112 V48 V112 4.2304280647233725e-12
C48_112 V48 V112 1.1125877737158301e-19

R48_113 V48 V113 1944.4848021507676
L48_113 V48 V113 -1.3372032846233636e-12
C48_113 V48 V113 -1.8074579377776803e-20

R48_114 V48 V114 1277.060244428878
L48_114 V48 V114 -1.6352651668092428e-12
C48_114 V48 V114 -2.124426036029009e-19

R48_115 V48 V115 661.0517098816431
L48_115 V48 V115 1.0781629005590683e-12
C48_115 V48 V115 3.4501309546803953e-19

R48_116 V48 V116 1339.254688924819
L48_116 V48 V116 8.86731700083682e-13
C48_116 V48 V116 -1.5989680003824986e-20

R48_117 V48 V117 2713.8447708570197
L48_117 V48 V117 1.5061280592743685e-12
C48_117 V48 V117 2.3918203602790676e-19

R48_118 V48 V118 -596.294083080282
L48_118 V48 V118 8.762308265594529e-13
C48_118 V48 V118 4.469601860998063e-19

R48_119 V48 V119 -1503.2753620068652
L48_119 V48 V119 4.7789403268852295e-12
C48_119 V48 V119 1.016022914073972e-19

R48_120 V48 V120 13144.071857779316
L48_120 V48 V120 -1.3426346703797184e-12
C48_120 V48 V120 3.4495688085377736e-19

R48_121 V48 V121 -3162.7759497107145
L48_121 V48 V121 3.4765557984550446e-12
C48_121 V48 V121 -1.2838447249145497e-19

R48_122 V48 V122 3336.448808578002
L48_122 V48 V122 -3.439101567421228e-12
C48_122 V48 V122 -1.1780624051423322e-19

R48_123 V48 V123 -1204.3912133664192
L48_123 V48 V123 -1.2140327945618964e-12
C48_123 V48 V123 -2.5601417679683715e-19

R48_124 V48 V124 -915.1519147901714
L48_124 V48 V124 -1.206852205958864e-12
C48_124 V48 V124 -6.101853730623674e-19

R48_125 V48 V125 -801.415652390076
L48_125 V48 V125 -2.2186704298908998e-12
C48_125 V48 V125 -5.768066053643218e-20

R48_126 V48 V126 1908.6724700457999
L48_126 V48 V126 -8.343502777776991e-13
C48_126 V48 V126 -2.973513187749161e-19

R48_127 V48 V127 739.5839804925048
L48_127 V48 V127 -2.099423741514114e-12
C48_127 V48 V127 -1.6264708288522339e-19

R48_128 V48 V128 717.6554332221781
L48_128 V48 V128 1.070948211389035e-12
C48_128 V48 V128 2.7021141405548424e-20

R48_129 V48 V129 610.2044910637147
L48_129 V48 V129 -1.4038464293456114e-12
C48_129 V48 V129 -3.1216273554314255e-19

R48_130 V48 V130 2145.4621595705325
L48_130 V48 V130 8.602598463336144e-13
C48_130 V48 V130 3.8436147616731525e-19

R48_131 V48 V131 -913.2768934044161
L48_131 V48 V131 1.1722467060924949e-12
C48_131 V48 V131 3.159968289991508e-19

R48_132 V48 V132 -801.6480971101553
L48_132 V48 V132 -5.434963867776904e-12
C48_132 V48 V132 4.592094977189709e-19

R48_133 V48 V133 1203.6158424703733
L48_133 V48 V133 1.5018502366922982e-12
C48_133 V48 V133 4.52101075430066e-19

R48_134 V48 V134 -1686.94300171836
L48_134 V48 V134 -4.220840393565589e-12
C48_134 V48 V134 -7.895153458718137e-20

R48_135 V48 V135 -9447.366727832425
L48_135 V48 V135 -1.4464082050259627e-10
C48_135 V48 V135 1.8262812407052535e-20

R48_136 V48 V136 -663.6399591698774
L48_136 V48 V136 -3.685314154060029e-12
C48_136 V48 V136 -5.533348783699626e-19

R48_137 V48 V137 -587.7521597608106
L48_137 V48 V137 1.0549303909525116e-12
C48_137 V48 V137 2.1135934006843247e-19

R48_138 V48 V138 2217.0714346435643
L48_138 V48 V138 -2.2466859505576725e-12
C48_138 V48 V138 -1.1239910937435932e-19

R48_139 V48 V139 630.6872543340413
L48_139 V48 V139 3.106638496261524e-11
C48_139 V48 V139 3.891472841160638e-20

R48_140 V48 V140 494.9422946110516
L48_140 V48 V140 2.1935907658683467e-12
C48_140 V48 V140 6.216116299149323e-19

R48_141 V48 V141 -943.3982524644777
L48_141 V48 V141 -7.79415204592266e-13
C48_141 V48 V141 -7.245667096384415e-19

R48_142 V48 V142 1149.9388934341055
L48_142 V48 V142 3.496718208208325e-12
C48_142 V48 V142 3.344112412791502e-20

R48_143 V48 V143 -866.5956116426022
L48_143 V48 V143 -2.7865268384599544e-12
C48_143 V48 V143 -1.533554063578073e-19

R48_144 V48 V144 475.5246183727053
L48_144 V48 V144 -9.815499480172602e-13
C48_144 V48 V144 -1.597008171037592e-19

R48_145 V48 V145 462.6886812120634
L48_145 V48 V145 -8.227294251983084e-13
C48_145 V48 V145 -1.927635490978935e-19

R48_146 V48 V146 -2281.332948906108
L48_146 V48 V146 -3.2598732297450923e-12
C48_146 V48 V146 1.0296225900797999e-19

R48_147 V48 V147 1170.469937445765
L48_147 V48 V147 -1.7732399498397556e-12
C48_147 V48 V147 -2.1123484126995405e-19

R48_148 V48 V148 -178.8659046211096
L48_148 V48 V148 -3.907277890795291e-11
C48_148 V48 V148 -4.5817409280174035e-19

R48_149 V48 V149 3124.505722873259
L48_149 V48 V149 4.686499986753962e-13
C48_149 V48 V149 8.254157799132308e-19

R48_150 V48 V150 -435.3929513871677
L48_150 V48 V150 -8.869344464013522e-12
C48_150 V48 V150 -4.847622758488168e-19

R48_151 V48 V151 -1071.6998346956784
L48_151 V48 V151 1.1112213401962441e-11
C48_151 V48 V151 1.1625183854521116e-19

R48_152 V48 V152 855.4125308991172
L48_152 V48 V152 7.538904894730545e-13
C48_152 V48 V152 1.3095760710515548e-19

R48_153 V48 V153 -2402.4240672445217
L48_153 V48 V153 1.090945788603441e-12
C48_153 V48 V153 1.9220403437104125e-19

R48_154 V48 V154 694.9681496991404
L48_154 V48 V154 1.4388831434491468e-12
C48_154 V48 V154 2.9164944912494876e-19

R48_155 V48 V155 368.81941481260054
L48_155 V48 V155 8.988925264946057e-13
C48_155 V48 V155 2.1722600188615873e-19

R48_156 V48 V156 -17127.586338591394
L48_156 V48 V156 -1.8361300623097498e-10
C48_156 V48 V156 3.945214329133861e-19

R48_157 V48 V157 -679.866672215978
L48_157 V48 V157 -6.746877723271921e-13
C48_157 V48 V157 -8.17252569470826e-19

R48_158 V48 V158 -1208.8467294588552
L48_158 V48 V158 4.0446548348954996e-12
C48_158 V48 V158 3.1549664334986095e-20

R48_159 V48 V159 -405.4065696659019
L48_159 V48 V159 3.4415803741377024e-12
C48_159 V48 V159 1.4303938855865198e-21

R48_160 V48 V160 358.08970353214124
L48_160 V48 V160 -6.613648670763946e-13
C48_160 V48 V160 -8.069406407539056e-20

R48_161 V48 V161 1169.2247173635901
L48_161 V48 V161 -2.69909419983766e-11
C48_161 V48 V161 -7.188242736634352e-20

R48_162 V48 V162 6539.566767303633
L48_162 V48 V162 3.927382529262308e-12
C48_162 V48 V162 1.1901458826941535e-19

R48_163 V48 V163 -64257.65397989791
L48_163 V48 V163 -1.665134468354139e-12
C48_163 V48 V163 -9.704524962949762e-20

R48_164 V48 V164 -184.6367802744405
L48_164 V48 V164 5.186841091610924e-12
C48_164 V48 V164 7.707445100475327e-20

R48_165 V48 V165 -1182.3462811871152
L48_165 V48 V165 -4.284934102777188e-11
C48_165 V48 V165 2.1248225977511263e-19

R48_166 V48 V166 -798.7743329530892
L48_166 V48 V166 -1.603199668337163e-12
C48_166 V48 V166 -2.637759347464842e-19

R48_167 V48 V167 -590.1718535933738
L48_167 V48 V167 -3.2941452151386433e-12
C48_167 V48 V167 -7.762294694013258e-20

R48_168 V48 V168 206.93108444456843
L48_168 V48 V168 9.054964279984232e-13
C48_168 V48 V168 -1.5091516552612055e-19

R48_169 V48 V169 -1258.250243185288
L48_169 V48 V169 4.938163708280082e-12
C48_169 V48 V169 -6.937828484911004e-20

R48_170 V48 V170 7422.103903974069
L48_170 V48 V170 2.49177908672015e-12
C48_170 V48 V170 2.1109460159759146e-19

R48_171 V48 V171 662.4724360284171
L48_171 V48 V171 1.1226057523913113e-12
C48_171 V48 V171 1.8823000284729736e-19

R48_172 V48 V172 2017.637831736546
L48_172 V48 V172 -4.35758891733651e-12
C48_172 V48 V172 1.1761821954292923e-19

R48_173 V48 V173 1662.592535668292
L48_173 V48 V173 2.447470105382516e-12
C48_173 V48 V173 6.208144210657329e-20

R48_174 V48 V174 526.8974577368972
L48_174 V48 V174 2.0172777824349574e-12
C48_174 V48 V174 -7.58654278192174e-20

R48_175 V48 V175 222136.45562751533
L48_175 V48 V175 2.293315793439711e-12
C48_175 V48 V175 2.006442395969555e-19

R48_176 V48 V176 -396.24620022519076
L48_176 V48 V176 9.158432131563938e-12
C48_176 V48 V176 3.7998991321671966e-19

R48_177 V48 V177 -1374.3986598994893
L48_177 V48 V177 -2.21615088557481e-12
C48_177 V48 V177 -7.434905725297184e-20

R48_178 V48 V178 -668.7032711023996
L48_178 V48 V178 -1.5798037704159682e-12
C48_178 V48 V178 -1.2859208910603415e-19

R48_179 V48 V179 -3460.5899936824376
L48_179 V48 V179 -1.15211760960037e-12
C48_179 V48 V179 -3.7811312860344957e-19

R48_180 V48 V180 799.3897772226879
L48_180 V48 V180 -7.429197930473111e-13
C48_180 V48 V180 -4.129264737721609e-19

R48_181 V48 V181 3432.300424923711
L48_181 V48 V181 8.403127543456364e-12
C48_181 V48 V181 -1.9292119589402204e-19

R48_182 V48 V182 1213.840801189969
L48_182 V48 V182 1.4708589262119778e-12
C48_182 V48 V182 1.595589226502521e-19

R48_183 V48 V183 -2141.3928404031494
L48_183 V48 V183 -1.4564708394113565e-12
C48_183 V48 V183 -8.55925347048935e-20

R48_184 V48 V184 -1367.3959666307467
L48_184 V48 V184 7.992560053119687e-12
C48_184 V48 V184 5.452597675568018e-20

R48_185 V48 V185 -12231.258037566884
L48_185 V48 V185 1.634246877119925e-11
C48_185 V48 V185 1.7035139987045813e-19

R48_186 V48 V186 2347.713360409938
L48_186 V48 V186 -2.2454531677930343e-12
C48_186 V48 V186 -9.601342181800941e-20

R48_187 V48 V187 1177.5536917298323
L48_187 V48 V187 1.924190063563298e-12
C48_187 V48 V187 3.415718556412293e-19

R48_188 V48 V188 542.25656588771
L48_188 V48 V188 4.919101354079812e-13
C48_188 V48 V188 1.8637840531133783e-19

R48_189 V48 V189 -3551.571910630254
L48_189 V48 V189 6.912216932434683e-12
C48_189 V48 V189 1.3650537380661555e-19

R48_190 V48 V190 -953.5737040939721
L48_190 V48 V190 -4.882599414921778e-11
C48_190 V48 V190 -1.8719920211275497e-19

R48_191 V48 V191 4154.677988979914
L48_191 V48 V191 8.766030633939536e-13
C48_191 V48 V191 9.660540126891498e-20

R48_192 V48 V192 6157.915279655938
L48_192 V48 V192 -1.0192935404936226e-12
C48_192 V48 V192 -3.197777655336707e-20

R48_193 V48 V193 979.8619001956166
L48_193 V48 V193 -1.9243691561692534e-11
C48_193 V48 V193 -9.068614996847553e-20

R48_194 V48 V194 -3738.6005100622656
L48_194 V48 V194 -3.727476942478415e-11
C48_194 V48 V194 -1.217391212034414e-19

R48_195 V48 V195 -876.1888352313739
L48_195 V48 V195 -7.143066526796291e-13
C48_195 V48 V195 -4.246763242164148e-19

R48_196 V48 V196 -422.2082759798269
L48_196 V48 V196 6.151036451371967e-12
C48_196 V48 V196 1.2271405275645507e-19

R48_197 V48 V197 505496.6845586712
L48_197 V48 V197 -2.6678976936254726e-12
C48_197 V48 V197 -1.5067259946248356e-19

R48_198 V48 V198 -1449.924764285921
L48_198 V48 V198 -3.2664526860464824e-11
C48_198 V48 V198 -2.636020339249597e-20

R48_199 V48 V199 -479.1359651616581
L48_199 V48 V199 -5.155554330698334e-12
C48_199 V48 V199 -6.721100163052742e-20

R48_200 V48 V200 372.58901533089823
L48_200 V48 V200 3.2184422286284466e-12
C48_200 V48 V200 -8.549045150346539e-20

R49_49 V49 0 164.96341349858753
L49_49 V49 0 9.416537183139408e-13
C49_49 V49 0 2.2944477691907665e-19

R49_50 V49 V50 9194.483330445586
L49_50 V49 V50 -2.5810937160763998e-12
C49_50 V49 V50 -1.6731456669129022e-19

R49_51 V49 V51 11966.46973674054
L49_51 V49 V51 -4.1192336408228395e-12
C49_51 V49 V51 -1.2220752346587433e-19

R49_52 V49 V52 7276.872768420831
L49_52 V49 V52 -3.4457926121393782e-12
C49_52 V49 V52 -1.4656553154276926e-19

R49_53 V49 V53 -2815.9170222784655
L49_53 V49 V53 4.068100916546549e-12
C49_53 V49 V53 2.366463556131159e-19

R49_54 V49 V54 -4588.387482852648
L49_54 V49 V54 2.587520815734022e-11
C49_54 V49 V54 1.203492126482099e-19

R49_55 V49 V55 -4163.863074143404
L49_55 V49 V55 9.878202070958364e-12
C49_55 V49 V55 1.374341006630839e-19

R49_56 V49 V56 -3504.9205952767998
L49_56 V49 V56 1.1111819189985277e-11
C49_56 V49 V56 1.554725764257973e-19

R49_57 V49 V57 5064.318109692499
L49_57 V49 V57 4.951336455385927e-12
C49_57 V49 V57 -4.2224303635413476e-20

R49_58 V49 V58 3559.4915521949524
L49_58 V49 V58 7.191627557381284e-12
C49_58 V49 V58 4.412890930830788e-21

R49_59 V49 V59 3972.8012128315218
L49_59 V49 V59 6.555353050351073e-12
C49_59 V49 V59 -2.408245132933832e-20

R49_60 V49 V60 2809.1990423253237
L49_60 V49 V60 4.355673710485669e-12
C49_60 V49 V60 -7.12133056402996e-21

R49_61 V49 V61 16919.704782885503
L49_61 V49 V61 -5.787919613357948e-12
C49_61 V49 V61 2.4883880647509452e-20

R49_62 V49 V62 -20529.090292289766
L49_62 V49 V62 -1.7699800224974578e-11
C49_62 V49 V62 -7.624685630778643e-20

R49_63 V49 V63 11876.946571658797
L49_63 V49 V63 -3.0224413666993334e-11
C49_63 V49 V63 -2.6300837788163304e-20

R49_64 V49 V64 15235.519289832951
L49_64 V49 V64 -2.8615751453014394e-11
C49_64 V49 V64 -4.220952424136419e-20

R49_65 V49 V65 -1108.5049880203876
L49_65 V49 V65 9.709216848233223e-12
C49_65 V49 V65 1.319938116168803e-19

R49_66 V49 V66 5239.933443835454
L49_66 V49 V66 -2.7830547356578335e-11
C49_66 V49 V66 2.595632910135403e-20

R49_67 V49 V67 6258.2367367963825
L49_67 V49 V67 -1.206577499198838e-11
C49_67 V49 V67 1.259014361525352e-20

R49_68 V49 V68 5157.826661874634
L49_68 V49 V68 -1.8809755898875537e-11
C49_68 V49 V68 4.176339838786573e-20

R49_69 V49 V69 -6693.603920351412
L49_69 V49 V69 -5.114542791525242e-12
C49_69 V49 V69 -1.929388040377232e-19

R49_70 V49 V70 22303.7525148186
L49_70 V49 V70 4.848995182374307e-11
C49_70 V49 V70 5.648407924349636e-20

R49_71 V49 V71 -18697.480200182345
L49_71 V49 V71 -4.4140284825657673e-10
C49_71 V49 V71 2.1401572191339336e-20

R49_72 V49 V72 -42970.87884403791
L49_72 V49 V72 -1.4921105285453535e-11
C49_72 V49 V72 1.7768466196343426e-22

R49_73 V49 V73 -1895.1900475791076
L49_73 V49 V73 3.427325982513888e-12
C49_73 V49 V73 1.6444868438011799e-19

R49_74 V49 V74 -3126.2070729071384
L49_74 V49 V74 -1.1680944643824526e-10
C49_74 V49 V74 -6.449780767267257e-20

R49_75 V49 V75 -8433.496784073848
L49_75 V49 V75 6.478051256775472e-12
C49_75 V49 V75 1.707845318154771e-20

R49_76 V49 V76 -5384.914933234738
L49_76 V49 V76 8.737636951770834e-12
C49_76 V49 V76 2.005160192234548e-20

R49_77 V49 V77 -5945.220871167088
L49_77 V49 V77 -4.208302343160034e-12
C49_77 V49 V77 -1.3276369673567354e-19

R49_78 V49 V78 3588.9292818498566
L49_78 V49 V78 2.3816811321517665e-11
C49_78 V49 V78 6.455072528415539e-20

R49_79 V49 V79 5649.997453296013
L49_79 V49 V79 -8.70696968793903e-12
C49_79 V49 V79 -7.382668106021102e-20

R49_80 V49 V80 3335.750356460013
L49_80 V49 V80 -2.1983671862047976e-11
C49_80 V49 V80 -7.057708181584746e-20

R49_81 V49 V81 -1801.1066451872264
L49_81 V49 V81 -4.4742236444707966e-11
C49_81 V49 V81 1.650591891407699e-20

R49_82 V49 V82 10385.526387538554
L49_82 V49 V82 -1.5420265336846578e-11
C49_82 V49 V82 -4.930046442259658e-20

R49_83 V49 V83 5607.907315488237
L49_83 V49 V83 -1.0905412458717993e-11
C49_83 V49 V83 -1.323300264847707e-20

R49_84 V49 V84 3886.981526426282
L49_84 V49 V84 -5.551848470257687e-11
C49_84 V49 V84 2.918422970545687e-21

R49_85 V49 V85 -3167.5098755210925
L49_85 V49 V85 4.098283505076464e-12
C49_85 V49 V85 2.060606748862452e-19

R49_86 V49 V86 10758.756262629708
L49_86 V49 V86 -2.0544090483572497e-11
C49_86 V49 V86 -1.2807711545057376e-20

R49_87 V49 V87 6186.793378192281
L49_87 V49 V87 1.3324445365046585e-11
C49_87 V49 V87 4.65597816607598e-20

R49_88 V49 V88 6762.6181482286265
L49_88 V49 V88 2.887664118794037e-11
C49_88 V49 V88 7.537674966813095e-20

R49_89 V49 V89 -1315.230164842875
L49_89 V49 V89 -8.387888400916208e-12
C49_89 V49 V89 -1.3984017676949215e-21

R49_90 V49 V90 7420.34497768177
L49_90 V49 V90 1.0488428824999095e-11
C49_90 V49 V90 9.830566838617841e-20

R49_91 V49 V91 4952.635905419364
L49_91 V49 V91 7.37887001547794e-12
C49_91 V49 V91 3.5797075187518905e-20

R49_92 V49 V92 7209.32804358987
L49_92 V49 V92 1.747747259332007e-11
C49_92 V49 V92 -3.7143510736608165e-20

R49_93 V49 V93 6289.297188150023
L49_93 V49 V93 -5.080775733578506e-12
C49_93 V49 V93 -2.5193746078277313e-19

R49_94 V49 V94 -4927.09427689528
L49_94 V49 V94 2.908216071482575e-11
C49_94 V49 V94 -7.445286108256739e-20

R49_95 V49 V95 -2697.52433561419
L49_95 V49 V95 -9.586663567666588e-12
C49_95 V49 V95 -6.45768613349264e-20

R49_96 V49 V96 -2019.6504869202993
L49_96 V49 V96 -7.764438781710344e-12
C49_96 V49 V96 -8.012576751590987e-20

R49_97 V49 V97 -1130.9056572102832
L49_97 V49 V97 1.7763085871154742e-12
C49_97 V49 V97 1.690032277220795e-19

R49_98 V49 V98 3238.327205842999
L49_98 V49 V98 -7.581363715811528e-12
C49_98 V49 V98 1.6478995613659924e-21

R49_99 V49 V99 1713.047551197107
L49_99 V49 V99 -8.384035210992994e-12
C49_99 V49 V99 -3.997778228199558e-20

R49_100 V49 V100 1048.3632513787436
L49_100 V49 V100 1.3931030465774867e-11
C49_100 V49 V100 5.749444176319068e-20

R49_101 V49 V101 -2538.15830813522
L49_101 V49 V101 -2.0478035143753705e-12
C49_101 V49 V101 -1.65702383518692e-20

R49_102 V49 V102 20254.36591791752
L49_102 V49 V102 -1.4003724002075716e-11
C49_102 V49 V102 -1.8034431331256815e-20

R49_103 V49 V103 7832.767740649663
L49_103 V49 V103 1.4926004474764265e-11
C49_103 V49 V103 1.0856363910933149e-20

R49_104 V49 V104 7367.979510976533
L49_104 V49 V104 1.3944064382401527e-11
C49_104 V49 V104 -1.0633065507371149e-20

R49_105 V49 V105 -1224.5414779228306
L49_105 V49 V105 -1.7473211917583293e-11
C49_105 V49 V105 5.605362591499316e-20

R49_106 V49 V106 1320.4848664685057
L49_106 V49 V106 5.3353684527971545e-12
C49_106 V49 V106 6.8227327043736e-20

R49_107 V49 V107 -23567.257952942033
L49_107 V49 V107 1.7189516696180965e-11
C49_107 V49 V107 6.732266855279065e-20

R49_108 V49 V108 -3072.4560067571138
L49_108 V49 V108 -8.851525341146108e-12
C49_108 V49 V108 5.875496604064893e-20

R49_109 V49 V109 1864.9817068535829
L49_109 V49 V109 1.7691507947207938e-12
C49_109 V49 V109 5.4179602570900107e-20

R49_110 V49 V110 -1682.0725407690447
L49_110 V49 V110 -7.43201844038272e-12
C49_110 V49 V110 1.1776971874573128e-20

R49_111 V49 V111 3221.664820512558
L49_111 V49 V111 6.245184666778796e-11
C49_111 V49 V111 -2.2059252815358622e-20

R49_112 V49 V112 2282.4528102993645
L49_112 V49 V112 2.0521117268060133e-11
C49_112 V49 V112 -9.20344173717077e-20

R49_113 V49 V113 -884.0616327656086
L49_113 V49 V113 -1.7921300737564505e-12
C49_113 V49 V113 -2.3713601056078463e-19

R49_114 V49 V114 -8433.888745212147
L49_114 V49 V114 5.669885820565324e-11
C49_114 V49 V114 -4.872529420622026e-20

R49_115 V49 V115 -5472.084353242996
L49_115 V49 V115 -2.1458898652759538e-11
C49_115 V49 V115 -2.914002479684881e-20

R49_116 V49 V116 -5427.622840950333
L49_116 V49 V116 2.111949504575264e-10
C49_116 V49 V116 -2.2456677621939485e-20

R49_117 V49 V117 -1816.6518899834775
L49_117 V49 V117 5.365751909293125e-12
C49_117 V49 V117 1.722432374288076e-19

R49_118 V49 V118 2011.8488765313218
L49_118 V49 V118 2.7006702366318593e-11
C49_118 V49 V118 2.0492043024417365e-21

R49_119 V49 V119 4186.8804642300975
L49_119 V49 V119 -2.37690894400923e-10
C49_119 V49 V119 6.06743280917284e-20

R49_120 V49 V120 2397.373705958573
L49_120 V49 V120 -1.7476515349681885e-11
C49_120 V49 V120 1.2186416112730706e-19

R49_121 V49 V121 1523.4100159725026
L49_121 V49 V121 -1.6971456362500305e-10
C49_121 V49 V121 -8.928205015512773e-20

R49_122 V49 V122 5505.06846955054
L49_122 V49 V122 1.2804106447843847e-10
C49_122 V49 V122 1.6078714381145812e-20

R49_123 V49 V123 5837.23943866393
L49_123 V49 V123 1.8838798509138893e-11
C49_123 V49 V123 -6.258847685314699e-20

R49_124 V49 V124 26773.857743201017
L49_124 V49 V124 1.7392855417386317e-11
C49_124 V49 V124 -1.5370599538737193e-19

R49_125 V49 V125 -856.0327062053474
L49_125 V49 V125 -4.86771620974915e-12
C49_125 V49 V125 1.9416369516838988e-20

R49_126 V49 V126 -5364.325953719643
L49_126 V49 V126 -9.383871165732875e-12
C49_126 V49 V126 2.8099718040578985e-20

R49_127 V49 V127 -2990.899125203636
L49_127 V49 V127 -1.4486760146253591e-11
C49_127 V49 V127 4.424703456698684e-20

R49_128 V49 V128 -1979.9029791496462
L49_128 V49 V128 -2.829056399425058e-11
C49_128 V49 V128 7.970536916746588e-20

R49_129 V49 V129 -2983.615595603792
L49_129 V49 V129 2.8394945069742855e-12
C49_129 V49 V129 2.1281651602563603e-19

R49_130 V49 V130 -4064.588705969549
L49_130 V49 V130 6.492988381932934e-11
C49_130 V49 V130 -8.444605657155639e-21

R49_131 V49 V131 4434.378269795702
L49_131 V49 V131 1.3004174715024466e-11
C49_131 V49 V131 -2.2387376792409035e-21

R49_132 V49 V132 1771.670871126461
L49_132 V49 V132 2.1988920314511272e-11
C49_132 V49 V132 -1.856879175840955e-20

R49_133 V49 V133 1378.0154748441676
L49_133 V49 V133 -3.094860278211411e-12
C49_133 V49 V133 -3.119747460761052e-19

R49_134 V49 V134 1109.0568405818728
L49_134 V49 V134 4.205894833785513e-12
C49_134 V49 V134 1.9249862450717783e-20

R49_135 V49 V135 4548.751491210919
L49_135 V49 V135 1.6458772090753626e-11
C49_135 V49 V135 -5.465438196408744e-20

R49_136 V49 V136 6294.221469156451
L49_136 V49 V136 1.0664538279349402e-11
C49_136 V49 V136 -1.3454963382698708e-19

R49_137 V49 V137 -1784.8029933351715
L49_137 V49 V137 -8.375158490216568e-12
C49_137 V49 V137 -3.237272661397477e-20

R49_138 V49 V138 -1020.1103835029182
L49_138 V49 V138 -3.351906044046423e-12
C49_138 V49 V138 -4.873363183831212e-20

R49_139 V49 V139 -3197.434863011166
L49_139 V49 V139 -3.552094552166581e-12
C49_139 V49 V139 2.110705455764778e-20

R49_140 V49 V140 -4662.137745612085
L49_140 V49 V140 -2.8302251376831395e-12
C49_140 V49 V140 8.399922819505961e-20

R49_141 V49 V141 1119.4335901083748
L49_141 V49 V141 1.660335785517981e-12
C49_141 V49 V141 2.800531165490835e-19

R49_142 V49 V142 24110.593517607787
L49_142 V49 V142 -1.6225064398661618e-11
C49_142 V49 V142 4.491165744055193e-20

R49_143 V49 V143 3055.7817562586242
L49_143 V49 V143 8.876364529204315e-12
C49_143 V49 V143 8.129490677110685e-21

R49_144 V49 V144 -24681.310806915706
L49_144 V49 V144 1.135401593621819e-11
C49_144 V49 V144 5.671955557582168e-20

R49_145 V49 V145 -559.6501623763212
L49_145 V49 V145 -3.5252748300867677e-12
C49_145 V49 V145 -1.167331678967525e-19

R49_146 V49 V146 1428.629598341176
L49_146 V49 V146 3.393078505963626e-12
C49_146 V49 V146 -4.239760981378362e-21

R49_147 V49 V147 -2271.0850702708976
L49_147 V49 V147 7.923442988673599e-12
C49_147 V49 V147 7.965905851990722e-21

R49_148 V49 V148 3190.422323031681
L49_148 V49 V148 4.277417005591077e-12
C49_148 V49 V148 -1.406863169794787e-20

R49_149 V49 V149 722.0597284404951
L49_149 V49 V149 -1.4446199463118356e-12
C49_149 V49 V149 1.3055053379047739e-20

R49_150 V49 V150 27706.382686005687
L49_150 V49 V150 -7.725868634342915e-11
C49_150 V49 V150 3.224592202277448e-20

R49_151 V49 V151 2677.7421851139566
L49_151 V49 V151 1.278452311043602e-11
C49_151 V49 V151 1.393370057123487e-20

R49_152 V49 V152 10703.396613864019
L49_152 V49 V152 -5.0460508161382636e-11
C49_152 V49 V152 -2.7072648055393134e-20

R49_153 V49 V153 -1479.47073391801
L49_153 V49 V153 2.1611911723371516e-12
C49_153 V49 V153 3.549998654498846e-20

R49_154 V49 V154 -51708.67601241712
L49_154 V49 V154 6.62765308325768e-11
C49_154 V49 V154 -2.886225403676016e-20

R49_155 V49 V155 -1604.2356903442608
L49_155 V49 V155 -1.024654436772638e-11
C49_155 V49 V155 5.670919008948053e-21

R49_156 V49 V156 2912.0526318176403
L49_156 V49 V156 -3.0261116384929175e-11
C49_156 V49 V156 1.9927950038439496e-20

R49_157 V49 V157 -1943.222348980189
L49_157 V49 V157 1.4267639959009882e-12
C49_157 V49 V157 -7.55873971786808e-20

R49_158 V49 V158 5980.0466120927495
L49_158 V49 V158 -1.1258223938751417e-11
C49_158 V49 V158 -1.371151470665481e-20

R49_159 V49 V159 1955.672229290055
L49_159 V49 V159 -1.7495356364959707e-11
C49_159 V49 V159 -5.421296045720829e-20

R49_160 V49 V160 -2824.149934909393
L49_160 V49 V160 -1.0808243273164707e-11
C49_160 V49 V160 -4.1517823182265626e-20

R49_161 V49 V161 -916.3086677958639
L49_161 V49 V161 -1.2593838122467002e-12
C49_161 V49 V161 -6.139819494813763e-20

R49_162 V49 V162 -9746.070566643424
L49_162 V49 V162 -5.35726598409839e-12
C49_162 V49 V162 -1.806742560013733e-20

R49_163 V49 V163 1853.2074190714254
L49_163 V49 V163 -1.0056700315751876e-11
C49_163 V49 V163 -1.6964972690364674e-20

R49_164 V49 V164 1195.9259831771897
L49_164 V49 V164 -1.218075818422362e-11
C49_164 V49 V164 1.3002479825642423e-20

R49_165 V49 V165 -2152.098677461639
L49_165 V49 V165 9.288039643420522e-12
C49_165 V49 V165 2.0092689552123914e-19

R49_166 V49 V166 921.0394634473878
L49_166 V49 V166 5.788105140769546e-12
C49_166 V49 V166 2.2274479306227525e-20

R49_167 V49 V167 3906.026176775949
L49_167 V49 V167 1.6294154091655547e-11
C49_167 V49 V167 2.6865080999628314e-20

R49_168 V49 V168 -5208.856218663089
L49_168 V49 V168 -2.69835903706905e-10
C49_168 V49 V168 7.101247018828263e-20

R49_169 V49 V169 1881.9417827508817
L49_169 V49 V169 3.244801418382662e-12
C49_169 V49 V169 -1.9222477863004484e-19

R49_170 V49 V170 -779.4553680959542
L49_170 V49 V170 -7.217064407038642e-12
C49_170 V49 V170 6.673397575354623e-21

R49_171 V49 V171 -788.8595593646697
L49_171 V49 V171 -1.1876469588435478e-11
C49_171 V49 V171 8.020700723668626e-21

R49_172 V49 V172 -1390.7739284921952
L49_172 V49 V172 -1.1373816193944736e-09
C49_172 V49 V172 -2.6452901212804816e-20

R49_173 V49 V173 -664.0360878594477
L49_173 V49 V173 -2.3826250884102108e-12
C49_173 V49 V173 2.0470761768928442e-20

R49_174 V49 V174 4078.7916795658493
L49_174 V49 V174 9.123694489799293e-12
C49_174 V49 V174 -2.000301447103033e-21

R49_175 V49 V175 798.5621972218825
L49_175 V49 V175 4.8887081216847686e-12
C49_175 V49 V175 -3.1764305280327146e-20

R49_176 V49 V176 853.9674566240813
L49_176 V49 V176 5.821297424365906e-12
C49_176 V49 V176 -3.26756819794716e-20

R49_177 V49 V177 1062.1689669392379
L49_177 V49 V177 3.385577519457842e-12
C49_177 V49 V177 6.327289880036041e-20

R49_178 V49 V178 2340.7444568169913
L49_178 V49 V178 1.5502182679360174e-11
C49_178 V49 V178 -3.0470448152637746e-20

R49_179 V49 V179 -2579.0301175470713
L49_179 V49 V179 -3.2243473207560106e-11
C49_179 V49 V179 -1.526794430330904e-21

R49_180 V49 V180 -2683.556259535741
L49_180 V49 V180 -7.613398861881635e-11
C49_180 V49 V180 -1.3456357065269107e-20

R49_181 V49 V181 4011.1151101463406
L49_181 V49 V181 -2.3184790075889332e-12
C49_181 V49 V181 3.7493131275684086e-20

R49_182 V49 V182 -1594.4433823428321
L49_182 V49 V182 -6.757111983001025e-12
C49_182 V49 V182 7.147000357451767e-22

R49_183 V49 V183 -20309.150619610115
L49_183 V49 V183 -1.0592627755602391e-10
C49_183 V49 V183 1.3865060494834027e-20

R49_184 V49 V184 -3961.412168962068
L49_184 V49 V184 -3.501048851804169e-11
C49_184 V49 V184 3.494474289442881e-20

R49_185 V49 V185 -471.24778897066113
L49_185 V49 V185 1.0952597942345378e-11
C49_185 V49 V185 -7.442496526245273e-20

R49_186 V49 V186 1469.7543818764743
L49_186 V49 V186 2.064392269300831e-11
C49_186 V49 V186 6.509166855659364e-20

R49_187 V49 V187 5157.514540295464
L49_187 V49 V187 6.933428836254843e-11
C49_187 V49 V187 -1.3603009942666582e-20

R49_188 V49 V188 -3635.6265774789595
L49_188 V49 V188 -1.2342352749736135e-11
C49_188 V49 V188 2.3805712352593596e-20

R49_189 V49 V189 362.9198498696859
L49_189 V49 V189 2.9129906968030238e-12
C49_189 V49 V189 -8.197914224718395e-20

R49_190 V49 V190 7148.291257932753
L49_190 V49 V190 -2.8000923114762237e-11
C49_190 V49 V190 -4.905161983159854e-21

R49_191 V49 V191 -1434.531543896077
L49_191 V49 V191 -2.986878555336317e-11
C49_191 V49 V191 -3.704603398816584e-20

R49_192 V49 V192 -3814.3643264112916
L49_192 V49 V192 1.0664156275861888e-11
C49_192 V49 V192 -1.1079723636029712e-19

R49_193 V49 V193 -1658.1631815373416
L49_193 V49 V193 -1.8630831827822125e-12
C49_193 V49 V193 1.1903861182797537e-20

R49_194 V49 V194 -1630.8138309445985
L49_194 V49 V194 7.985872711670751e-12
C49_194 V49 V194 -4.9957155990993075e-20

R49_195 V49 V195 3091.554230612716
L49_195 V49 V195 7.372575532626525e-12
C49_195 V49 V195 4.0906204846939973e-20

R49_196 V49 V196 1497.5053352552295
L49_196 V49 V196 5.603270097521945e-12
C49_196 V49 V196 9.675636980762718e-20

R49_197 V49 V197 -845.8136458674517
L49_197 V49 V197 1.1161927449273087e-11
C49_197 V49 V197 1.0212799726776008e-19

R49_198 V49 V198 1604.3606737144778
L49_198 V49 V198 7.170100433342107e-11
C49_198 V49 V198 2.1639824410944834e-21

R49_199 V49 V199 987.732918519326
L49_199 V49 V199 -2.308890513417125e-11
C49_199 V49 V199 -1.1027133912470879e-20

R49_200 V49 V200 68523.78882161452
L49_200 V49 V200 -5.297548023193461e-12
C49_200 V49 V200 3.807604788407266e-20

R50_50 V50 0 7065.4686080244755
L50_50 V50 0 -1.7256962933657381e-12
C50_50 V50 0 -1.468729673635517e-19

R50_51 V50 V51 -28569.241554514763
L50_51 V50 V51 -3.1800763678424246e-12
C50_51 V50 V51 -1.6655719102788927e-19

R50_52 V50 V52 -512567.986101318
L50_52 V50 V52 -2.6723394805127553e-12
C50_52 V50 V52 -2.12306424101106e-19

R50_53 V50 V53 -186840.73616324115
L50_53 V50 V53 1.745218187409007e-11
C50_53 V50 V53 1.7652385124009192e-19

R50_54 V50 V54 3347.393718550223
L50_54 V50 V54 6.188254247986665e-12
C50_54 V50 V54 2.386776293835008e-19

R50_55 V50 V55 372739.98872180766
L50_55 V50 V55 5.908660456502107e-12
C50_55 V50 V55 1.869977309981318e-19

R50_56 V50 V56 -916915.2164680351
L50_56 V50 V56 1.1731115567041903e-11
C50_56 V50 V56 1.7137304129356845e-19

R50_57 V50 V57 -37728.41185838746
L50_57 V50 V57 6.6016054023917535e-12
C50_57 V50 V57 3.08667117421491e-20

R50_58 V50 V58 -89094.99866128842
L50_58 V50 V58 2.227659152939458e-12
C50_58 V50 V58 3.0073315063273374e-19

R50_59 V50 V59 207740.99451600979
L50_59 V50 V59 4.719236118434143e-12
C50_59 V50 V59 8.63669478679138e-20

R50_60 V50 V60 -72643.66740064211
L50_60 V50 V60 2.8018907218353575e-12
C50_60 V50 V60 1.5145598215553603e-19

R50_61 V50 V61 86133.2761872349
L50_61 V50 V61 -1.0664846885678836e-11
C50_61 V50 V61 -9.067611187067839e-20

R50_62 V50 V62 3654.334534298134
L50_62 V50 V62 -1.1574997152985787e-11
C50_62 V50 V62 -1.8937502863273626e-19

R50_63 V50 V63 77905.44811635213
L50_63 V50 V63 -7.628499109820991e-12
C50_63 V50 V63 -8.494716219252976e-20

R50_64 V50 V64 -102233.41496299587
L50_64 V50 V64 -9.523552677382125e-12
C50_64 V50 V64 -1.1707474068119115e-19

R50_65 V50 V65 13640.976194423829
L50_65 V50 V65 1.5641079489359517e-11
C50_65 V50 V65 4.359865668946196e-20

R50_66 V50 V66 -2081.3281360503843
L50_66 V50 V66 -1.2654026973339395e-11
C50_66 V50 V66 6.516027879246701e-21

R50_67 V50 V67 -25079.207433116197
L50_67 V50 V67 -8.578168025366442e-12
C50_67 V50 V67 -5.609253600565041e-20

R50_68 V50 V68 -40254.37142575346
L50_68 V50 V68 -2.3175173645664e-11
C50_68 V50 V68 -5.832086632671663e-20

R50_69 V50 V69 75229.91269605802
L50_69 V50 V69 -5.036299663366777e-12
C50_69 V50 V69 -2.973360430286507e-20

R50_70 V50 V70 -5473.178563164628
L50_70 V50 V70 -1.1271093144020926e-11
C50_70 V50 V70 5.119412100504077e-22

R50_71 V50 V71 -490373.2217071827
L50_71 V50 V71 8.296499336716974e-12
C50_71 V50 V71 3.5041318371786975e-20

R50_72 V50 V72 30222.58570039178
L50_72 V50 V72 1.4605480960759357e-11
C50_72 V50 V72 3.510712467108968e-20

R50_73 V50 V73 -9715.991850973105
L50_73 V50 V73 -1.5218108986730643e-10
C50_73 V50 V73 1.5578786538550352e-20

R50_74 V50 V74 1637.3083620491961
L50_74 V50 V74 -6.286410874721093e-11
C50_74 V50 V74 -7.643248020214837e-20

R50_75 V50 V75 117237.7451348596
L50_75 V50 V75 8.283296701566802e-12
C50_75 V50 V75 8.156700047840088e-20

R50_76 V50 V76 -126888.15264678826
L50_76 V50 V76 -1.8935752977529893e-11
C50_76 V50 V76 5.332406627283163e-20

R50_77 V50 V77 9156.976967235787
L50_77 V50 V77 6.806961521722945e-12
C50_77 V50 V77 3.2391388785285345e-20

R50_78 V50 V78 -1741.7841093639731
L50_78 V50 V78 -5.799362691900348e-12
C50_78 V50 V78 4.269666606567805e-20

R50_79 V50 V79 -29138.17971740826
L50_79 V50 V79 -6.464287807885736e-12
C50_79 V50 V79 -2.6306762679573495e-20

R50_80 V50 V80 -13772.580299411387
L50_80 V50 V80 -1.7079327038389357e-10
C50_80 V50 V80 -1.0462139712999352e-20

R50_81 V50 V81 -11136.347474678054
L50_81 V50 V81 -1.1378313259927861e-11
C50_81 V50 V81 1.5452719791421566e-20

R50_82 V50 V82 5943.38235575511
L50_82 V50 V82 2.3392851804064265e-12
C50_82 V50 V82 1.443606087986536e-19

R50_83 V50 V83 -138289.91190303367
L50_83 V50 V83 -2.312471005282917e-11
C50_83 V50 V83 -7.97741926460481e-20

R50_84 V50 V84 -18452.92119597654
L50_84 V50 V84 6.531359294174185e-12
C50_84 V50 V84 -4.15190300966135e-20

R50_85 V50 V85 9795.833100420901
L50_85 V50 V85 1.7600942563761386e-11
C50_85 V50 V85 -7.70348143537297e-21

R50_86 V50 V86 -21721.19702075551
L50_86 V50 V86 3.957091979515549e-12
C50_86 V50 V86 -5.802823804754937e-20

R50_87 V50 V87 10778.115927391076
L50_87 V50 V87 7.762249972983007e-12
C50_87 V50 V87 1.6715116799127836e-20

R50_88 V50 V88 5739.033681137538
L50_88 V50 V88 2.723578621615361e-11
C50_88 V50 V88 1.8663752156833354e-20

R50_89 V50 V89 16030.916797533111
L50_89 V50 V89 -3.3000551951079376e-12
C50_89 V50 V89 -8.178742004732857e-20

R50_90 V50 V90 -6200.00119864632
L50_90 V50 V90 -1.0408604324822236e-12
C50_90 V50 V90 -2.4588251370189897e-19

R50_91 V50 V91 -34055.381715443866
L50_91 V50 V91 5.7647214478744897e-11
C50_91 V50 V91 7.689668567665347e-20

R50_92 V50 V92 1060219.3679426808
L50_92 V50 V92 -1.5765586157200285e-11
C50_92 V50 V92 -6.517737411340185e-21

R50_93 V50 V93 -20333.633434518324
L50_93 V50 V93 1.6647125720815555e-11
C50_93 V50 V93 4.834998730113475e-20

R50_94 V50 V94 2687.29003533937
L50_94 V50 V94 2.16458776426648e-12
C50_94 V50 V94 2.319879401880331e-19

R50_95 V50 V95 -8431.685537113688
L50_95 V50 V95 -1.8046419754856178e-11
C50_95 V50 V95 1.3611820354953594e-20

R50_96 V50 V96 -4237.999713968728
L50_96 V50 V96 -1.1333005774275633e-11
C50_96 V50 V96 2.5920058579154715e-20

R50_97 V50 V97 4268.542428208335
L50_97 V50 V97 3.3115481412175687e-12
C50_97 V50 V97 1.514101237468399e-19

R50_98 V50 V98 -5602.636808402872
L50_98 V50 V98 2.3155610864382746e-12
C50_98 V50 V98 1.0153473961664942e-19

R50_99 V50 V99 5724.1485304872685
L50_99 V50 V99 -7.580920632623982e-12
C50_99 V50 V99 -1.2931984861293028e-19

R50_100 V50 V100 4276.2647945679755
L50_100 V50 V100 4.73520007588848e-12
C50_100 V50 V100 -1.3396773370651788e-20

R50_101 V50 V101 -2689.5199178832563
L50_101 V50 V101 -2.1021945237523335e-12
C50_101 V50 V101 -1.3812265074670124e-19

R50_102 V50 V102 -12284.16523334811
L50_102 V50 V102 -1.253238907101022e-12
C50_102 V50 V102 -3.262970500437827e-19

R50_103 V50 V103 11647.130548283907
L50_103 V50 V103 1.5192170476094432e-11
C50_103 V50 V103 8.251436175898589e-21

R50_104 V50 V104 13155.99583046372
L50_104 V50 V104 7.115782489207716e-12
C50_104 V50 V104 -2.6616460513211744e-21

R50_105 V50 V105 2957.458178155387
L50_105 V50 V105 7.194620663006704e-11
C50_105 V50 V105 -6.594117569560298e-20

R50_106 V50 V106 -3069.4050144507096
L50_106 V50 V106 1.9595168047506997e-12
C50_106 V50 V106 1.4807860408145778e-19

R50_107 V50 V107 -3941.288015387455
L50_107 V50 V107 4.7649148553255046e-11
C50_107 V50 V107 8.365742808884839e-20

R50_108 V50 V108 -4954.664834054616
L50_108 V50 V108 -2.5968369921168023e-12
C50_108 V50 V108 -2.6718013641059944e-20

R50_109 V50 V109 3391.4330143200755
L50_109 V50 V109 5.099467122512913e-12
C50_109 V50 V109 9.602831987598698e-20

R50_110 V50 V110 4953.181554870854
L50_110 V50 V110 -1.2807823059849535e-10
C50_110 V50 V110 1.857615159976899e-19

R50_111 V50 V111 -11509.434636803107
L50_111 V50 V111 6.092021408122231e-12
C50_111 V50 V111 1.4411121550320735e-21

R50_112 V50 V112 -24563.88140697296
L50_112 V50 V112 5.7928793884593634e-12
C50_112 V50 V112 -2.3227763901451937e-20

R50_113 V50 V113 -1762.2803396534325
L50_113 V50 V113 -3.2269608294291385e-12
C50_113 V50 V113 7.893802489368318e-20

R50_114 V50 V114 17186.10746348591
L50_114 V50 V114 -2.9462961586849847e-12
C50_114 V50 V114 -1.385782873187613e-19

R50_115 V50 V115 3598.6073639994147
L50_115 V50 V115 -4.176677529558731e-12
C50_115 V50 V115 -7.957329402298347e-20

R50_116 V50 V116 6762.67890844919
L50_116 V50 V116 1.2503985364678207e-11
C50_116 V50 V116 4.7369856527699466e-20

R50_117 V50 V117 -123485.7235896572
L50_117 V50 V117 1.9118065970475516e-11
C50_117 V50 V117 -3.0348013905780125e-20

R50_118 V50 V118 2335.23420834911
L50_118 V50 V118 2.3379886277127645e-12
C50_118 V50 V118 -1.770180214171065e-19

R50_119 V50 V119 40099.458495507984
L50_119 V50 V119 -1.794143171120512e-11
C50_119 V50 V119 1.3202362079679347e-20

R50_120 V50 V120 5929.7851984792305
L50_120 V50 V120 -3.5487892719653177e-12
C50_120 V50 V120 -2.7043610103154938e-20

R50_121 V50 V121 2568.284465324391
L50_121 V50 V121 -1.3353263150888668e-11
C50_121 V50 V121 -1.1078134079234541e-19

R50_122 V50 V122 -2045.18056488763
L50_122 V50 V122 -2.780507717370316e-11
C50_122 V50 V122 2.3098660194032192e-19

R50_123 V50 V123 -3738.8948732545978
L50_123 V50 V123 3.177156988944225e-12
C50_123 V50 V123 3.626886224245926e-20

R50_124 V50 V124 -2495.079991183665
L50_124 V50 V124 3.084916801215896e-12
C50_124 V50 V124 -4.127577115372024e-20

R50_125 V50 V125 4340.630031687535
L50_125 V50 V125 -1.7024149954178357e-11
C50_125 V50 V125 -7.938252400823714e-21

R50_126 V50 V126 -1161.503304716623
L50_126 V50 V126 -3.174493930986917e-12
C50_126 V50 V126 6.378490000902494e-20

R50_127 V50 V127 -8536.18424253118
L50_127 V50 V127 -4.600046441742007e-12
C50_127 V50 V127 -1.0570117301558524e-20

R50_128 V50 V128 -6062.244083462108
L50_128 V50 V128 -7.379148641774087e-12
C50_128 V50 V128 4.401486014327933e-20

R50_129 V50 V129 -1800.1695677034124
L50_129 V50 V129 7.354337660883906e-12
C50_129 V50 V129 1.8458827703106596e-19

R50_130 V50 V130 1040.6707463226119
L50_130 V50 V130 1.506311941183896e-11
C50_130 V50 V130 -2.1801074863190234e-19

R50_131 V50 V131 2760.1770004581413
L50_131 V50 V131 6.486318700480888e-12
C50_131 V50 V131 -9.901962775451184e-22

R50_132 V50 V132 1669.182116828078
L50_132 V50 V132 2.0572000041880404e-11
C50_132 V50 V132 -2.3682481594144695e-20

R50_133 V50 V133 -27215.014991160617
L50_133 V50 V133 -4.347256420023166e-12
C50_133 V50 V133 -7.739463739834879e-20

R50_134 V50 V134 14356.33180223617
L50_134 V50 V134 3.463881419989598e-12
C50_134 V50 V134 2.0181242474430682e-19

R50_135 V50 V135 57571.215899035444
L50_135 V50 V135 5.171617086079387e-12
C50_135 V50 V135 1.8572586214808503e-20

R50_136 V50 V136 14934.189272194102
L50_136 V50 V136 3.031276400521825e-12
C50_136 V50 V136 -9.564133189174795e-21

R50_137 V50 V137 3437.007081359646
L50_137 V50 V137 -8.56102616024882e-12
C50_137 V50 V137 -1.2841992788165553e-19

R50_138 V50 V138 -1522.083834333268
L50_138 V50 V138 -6.640492032125617e-12
C50_138 V50 V138 -3.0186996886400373e-20

R50_139 V50 V139 -2726.8361891147447
L50_139 V50 V139 -1.405055404531792e-12
C50_139 V50 V139 -7.627570290927738e-20

R50_140 V50 V140 -1533.9668293546026
L50_140 V50 V140 -1.337635974610296e-12
C50_140 V50 V140 2.5487153365292106e-22

R50_141 V50 V141 2900.1491094693015
L50_141 V50 V141 1.5127220145578563e-12
C50_141 V50 V141 1.640553333429146e-19

R50_142 V50 V142 2753.3584844784973
L50_142 V50 V142 -4.94156896084638e-12
C50_142 V50 V142 -5.795223240687527e-20

R50_143 V50 V143 16640.676424335878
L50_143 V50 V143 2.324914094050349e-12
C50_143 V50 V143 9.271082287671644e-20

R50_144 V50 V144 6937.061077224238
L50_144 V50 V144 4.50404217263849e-12
C50_144 V50 V144 3.322690849047229e-20

R50_145 V50 V145 -2840.0504777664432
L50_145 V50 V145 2.8445374197983186e-11
C50_145 V50 V145 9.434196887419297e-20

R50_146 V50 V146 -1089.0293880567417
L50_146 V50 V146 1.926977303163384e-12
C50_146 V50 V146 -1.986498287159001e-20

R50_147 V50 V147 713781.287159961
L50_147 V50 V147 2.147543352399888e-12
C50_147 V50 V147 2.7084987815642504e-20

R50_148 V50 V148 -4965.08074322751
L50_148 V50 V148 1.7864813804022433e-12
C50_148 V50 V148 -2.477774985967721e-21

R50_149 V50 V149 -1721.9435382392155
L50_149 V50 V149 -7.383209044392981e-13
C50_149 V50 V149 -3.258535300798069e-19

R50_150 V50 V150 623.2800636821916
L50_150 V50 V150 -5.025821384140777e-12
C50_150 V50 V150 1.4039628846372184e-19

R50_151 V50 V151 6016.709865675799
L50_151 V50 V151 -4.707108229091634e-12
C50_151 V50 V151 -6.90565758928937e-20

R50_152 V50 V152 1882.4252955529048
L50_152 V50 V152 -6.8070512325399985e-12
C50_152 V50 V152 1.4743456984512604e-20

R50_153 V50 V153 2240.863335878079
L50_153 V50 V153 1.1724609598723379e-11
C50_153 V50 V153 2.5163397963177664e-20

R50_154 V50 V154 -3338.6603753019986
L50_154 V50 V154 -8.067385126620665e-12
C50_154 V50 V154 -8.399313276443306e-20

R50_155 V50 V155 -52846.40251119077
L50_155 V50 V155 -1.9142480418073717e-12
C50_155 V50 V155 -5.859439119939285e-20

R50_156 V50 V156 -1754.2544780097046
L50_156 V50 V156 -3.471015224900469e-12
C50_156 V50 V156 -2.4794530516946197e-20

R50_157 V50 V157 1193.007771004329
L50_157 V50 V157 7.725966940193233e-13
C50_157 V50 V157 2.885070399916189e-19

R50_158 V50 V158 -1798.897218749112
L50_158 V50 V158 3.841084258955597e-12
C50_158 V50 V158 8.241605226153081e-21

R50_159 V50 V159 -2550.269591500507
L50_159 V50 V159 3.9562690542436715e-12
C50_159 V50 V159 4.238276581862877e-21

R50_160 V50 V160 -5111.972149797967
L50_160 V50 V160 1.465697657759323e-11
C50_160 V50 V160 -4.6156475379954057e-20

R50_161 V50 V161 -2254.616329271538
L50_161 V50 V161 -2.7523920966006037e-12
C50_161 V50 V161 -4.1104627279622944e-20

R50_162 V50 V162 -2270.858188833408
L50_162 V50 V162 -3.1113162982022187e-12
C50_162 V50 V162 -4.734271297864312e-20

R50_163 V50 V163 -8490.013229958273
L50_163 V50 V163 5.249306374180184e-12
C50_163 V50 V163 6.585845732100196e-20

R50_164 V50 V164 -6765.732124195332
L50_164 V50 V164 7.118425505282888e-12
C50_164 V50 V164 1.473197447745792e-20

R50_165 V50 V165 -1911.249366507454
L50_165 V50 V165 -1.4394937147691413e-12
C50_165 V50 V165 -1.7273704115130166e-19

R50_166 V50 V166 1690.7261526975658
L50_166 V50 V166 -3.2046206119429323e-12
C50_166 V50 V166 1.4876141205123662e-20

R50_167 V50 V167 -43177.88839837428
L50_167 V50 V167 -1.6548118016806933e-11
C50_167 V50 V167 -5.59902633089308e-22

R50_168 V50 V168 -27347.20352985957
L50_168 V50 V168 -6.3545659899543125e-12
C50_168 V50 V168 4.5480878753941977e-20

R50_169 V50 V169 1278.3337340224055
L50_169 V50 V169 2.0584883820373436e-12
C50_169 V50 V169 4.4049067990755415e-20

R50_170 V50 V170 4235.476145525956
L50_170 V50 V170 2.189182293569649e-12
C50_170 V50 V170 -9.65904640576811e-20

R50_171 V50 V171 4576.55332719578
L50_171 V50 V171 -3.800640217839133e-12
C50_171 V50 V171 -1.4756182112975427e-19

R50_172 V50 V172 14230.771063325748
L50_172 V50 V172 5.7092427657227805e-11
C50_172 V50 V172 -7.921213961975759e-20

R50_173 V50 V173 -3056.234120918218
L50_173 V50 V173 5.159178246201175e-12
C50_173 V50 V173 8.744879923972782e-20

R50_174 V50 V174 273126.2335654915
L50_174 V50 V174 8.308772197106595e-12
C50_174 V50 V174 9.755062792810439e-20

R50_175 V50 V175 6644.663942798582
L50_175 V50 V175 8.835320839512013e-12
C50_175 V50 V175 9.824329022597298e-21

R50_176 V50 V176 21785.315208569806
L50_176 V50 V176 8.04736671825987e-12
C50_176 V50 V176 2.9087961426150756e-20

R50_177 V50 V177 -1065.2672726369858
L50_177 V50 V177 -3.119597673076247e-12
C50_177 V50 V177 -8.096943699463073e-20

R50_178 V50 V178 -1615.4730698388453
L50_178 V50 V178 -2.928115429338628e-12
C50_178 V50 V178 6.220898849593709e-20

R50_179 V50 V179 -3142.7939972248028
L50_179 V50 V179 4.512350845369019e-12
C50_179 V50 V179 1.414945022567347e-19

R50_180 V50 V180 -2153.0509923580594
L50_180 V50 V180 9.381427910347614e-12
C50_180 V50 V180 7.185202187502447e-20

R50_181 V50 V181 1382.1958492785684
L50_181 V50 V181 7.473782187953919e-12
C50_181 V50 V181 1.7632931292768793e-20

R50_182 V50 V182 1244.7402632591982
L50_182 V50 V182 -7.98851016524223e-12
C50_182 V50 V182 -8.412002953503035e-20

R50_183 V50 V183 -3390.7988803397625
L50_183 V50 V183 4.5100009446225115e-12
C50_183 V50 V183 1.774276398638e-20

R50_184 V50 V184 -13529.906822988576
L50_184 V50 V184 1.1730654148527073e-11
C50_184 V50 V184 -1.0041042197091712e-20

R50_185 V50 V185 1704.610462478788
L50_185 V50 V185 5.11079572010526e-12
C50_185 V50 V185 2.843768837894327e-20

R50_186 V50 V186 1250.930390000182
L50_186 V50 V186 7.456193213390097e-12
C50_186 V50 V186 -2.774320094455892e-20

R50_187 V50 V187 2477.969293728255
L50_187 V50 V187 -2.848641283111214e-12
C50_187 V50 V187 -1.2049230115733093e-19

R50_188 V50 V188 2174.6757803030823
L50_188 V50 V188 -2.441579386142882e-12
C50_188 V50 V188 -8.615477277660551e-20

R50_189 V50 V189 -939.9661903478162
L50_189 V50 V189 -3.1337942674431693e-12
C50_189 V50 V189 -9.062268846794529e-20

R50_190 V50 V190 -1060.7293431768655
L50_190 V50 V190 -4.116155770105263e-12
C50_190 V50 V190 8.362764593624501e-20

R50_191 V50 V191 9560.990351054172
L50_191 V50 V191 -2.307554505460507e-12
C50_191 V50 V191 -8.112985195581996e-20

R50_192 V50 V192 -3819.4077061366756
L50_192 V50 V192 -1.0865788068383088e-11
C50_192 V50 V192 -5.3343974480673615e-20

R50_193 V50 V193 -11882.193791036263
L50_193 V50 V193 -1.3345856150418553e-11
C50_193 V50 V193 7.098532367969676e-20

R50_194 V50 V194 1432.7577835063412
L50_194 V50 V194 1.6987803201249587e-12
C50_194 V50 V194 3.900686452835589e-20

R50_195 V50 V195 -6480.909892811855
L50_195 V50 V195 1.5119526738324434e-12
C50_195 V50 V195 1.4235659209259666e-19

R50_196 V50 V196 -19038.101430027633
L50_196 V50 V196 1.79233742077386e-12
C50_196 V50 V196 1.8134428412575278e-19

R50_197 V50 V197 2034.048298712402
L50_197 V50 V197 2.7116947011818307e-12
C50_197 V50 V197 3.9129058633208547e-20

R50_198 V50 V198 1010.2673785052299
L50_198 V50 V198 -1.7290210109315848e-11
C50_198 V50 V198 -6.305514401877913e-20

R50_199 V50 V199 49521.63634205735
L50_199 V50 V199 6.340819738013398e-12
C50_199 V50 V199 5.403961982465141e-20

R50_200 V50 V200 -3682.52275768636
L50_200 V50 V200 -3.725304598106283e-11
C50_200 V50 V200 1.3395981109271989e-21

R51_51 V51 0 -2568.9142293000673
L51_51 V51 0 8.802197046465316e-13
C51_51 V51 0 -4.778969684656087e-20

R51_52 V51 V52 -10299.28930900873
L51_52 V51 V52 -7.205696209631319e-12
C51_52 V51 V52 -1.534880497890745e-19

R51_53 V51 V53 -42002.81090198475
L51_53 V51 V53 9.008831833034194e-12
C51_53 V51 V53 1.5857215033863694e-19

R51_54 V51 V54 -34003.63571404952
L51_54 V51 V54 4.1523954399309644e-12
C51_54 V51 V54 1.7439828979293781e-19

R51_55 V51 V55 3009.8011464616557
L51_55 V51 V55 4.4029141373901456e-12
C51_55 V51 V55 2.1242470897326117e-19

R51_56 V51 V56 13478.061971361982
L51_56 V51 V56 3.4866333745085085e-12
C51_56 V51 V56 2.0943027647693302e-19

R51_57 V51 V57 71917.62313450569
L51_57 V51 V57 4.204524163867748e-12
C51_57 V51 V57 7.462273098774333e-20

R51_58 V51 V58 -14113.973189395796
L51_58 V51 V58 3.5898294093302895e-11
C51_58 V51 V58 -1.6004396302039527e-21

R51_59 V51 V59 1962.528945312674
L51_59 V51 V59 6.959728130682085e-13
C51_59 V51 V59 9.914641143142576e-19

R51_60 V51 V60 4618.5303448672385
L51_60 V51 V60 5.9992814509214225e-12
C51_60 V51 V60 1.0453414988030067e-19

R51_61 V51 V61 60668.83039170663
L51_61 V51 V61 -3.4326838115690915e-12
C51_61 V51 V61 -1.8488942350146672e-19

R51_62 V51 V62 8351.394786317458
L51_62 V51 V62 -2.93886246306924e-11
C51_62 V51 V62 -2.0233056855811624e-20

R51_63 V51 V63 -8293.706071766448
L51_63 V51 V63 -1.0357277558156421e-12
C51_63 V51 V63 -8.4750549114983925e-19

R51_64 V51 V64 -10168.878479389281
L51_64 V51 V64 -5.607805143172059e-12
C51_64 V51 V64 -1.4482096435738953e-19

R51_65 V51 V65 11894.027614149089
L51_65 V51 V65 1.6806826111968313e-11
C51_65 V51 V65 5.915321030105649e-20

R51_66 V51 V66 -16637.39665615943
L51_66 V51 V66 9.606811457972833e-12
C51_66 V51 V66 7.54171153312637e-20

R51_67 V51 V67 -1891.7996078298945
L51_67 V51 V67 -2.2055891667005435e-12
C51_67 V51 V67 -2.308770636227456e-19

R51_68 V51 V68 -5315.161299159857
L51_68 V51 V68 1.3864032565850433e-11
C51_68 V51 V68 -1.7514034684611093e-20

R51_69 V51 V69 -6273.820446216375
L51_69 V51 V69 5.043115560850674e-11
C51_69 V51 V69 7.909133587651233e-20

R51_70 V51 V70 -94689.2132786381
L51_70 V51 V70 -4.9950629109850486e-12
C51_70 V51 V70 -1.341646440289848e-19

R51_71 V51 V71 14525.469637073367
L51_71 V51 V71 1.1111944356666991e-12
C51_71 V51 V71 7.571354306653044e-19

R51_72 V51 V72 -121957.90252768098
L51_72 V51 V72 -4.998964023331951e-12
C51_72 V51 V72 -9.405266926109922e-20

R51_73 V51 V73 31504.213182962187
L51_73 V51 V73 -1.4681309011021368e-11
C51_73 V51 V73 -5.546874475144438e-20

R51_74 V51 V74 9575.246180891994
L51_74 V51 V74 1.7523275682514758e-11
C51_74 V51 V74 3.8828653956943395e-20

R51_75 V51 V75 1667.7102132078514
L51_75 V51 V75 -4.831693205824256e-12
C51_75 V51 V75 -3.310971409910096e-19

R51_76 V51 V76 4844.649020353467
L51_76 V51 V76 8.279772729412588e-12
C51_76 V51 V76 1.6335167679224987e-19

R51_77 V51 V77 3147.592949599459
L51_77 V51 V77 8.740940778723694e-12
C51_77 V51 V77 6.04496211254459e-20

R51_78 V51 V78 -9861.536293591613
L51_78 V51 V78 5.936835226263316e-11
C51_78 V51 V78 1.1138651260034643e-19

R51_79 V51 V79 -1845.543705893645
L51_79 V51 V79 -2.0847596183679513e-12
C51_79 V51 V79 -2.6072914936503677e-19

R51_80 V51 V80 -24236.428762981985
L51_80 V51 V80 1.1015732842229286e-11
C51_80 V51 V80 1.8436011420683756e-20

R51_81 V51 V81 -3287.796122244415
L51_81 V51 V81 -5.654828723917329e-12
C51_81 V51 V81 -1.6213147674128437e-20

R51_82 V51 V82 43319.76626584593
L51_82 V51 V82 3.0834773097601775e-11
C51_82 V51 V82 1.241645802089942e-21

R51_83 V51 V83 12670.207289325956
L51_83 V51 V83 2.3174954241624675e-12
C51_83 V51 V83 3.85423708625754e-19

R51_84 V51 V84 -8262.616103642493
L51_84 V51 V84 -3.838572476681555e-11
C51_84 V51 V84 -7.428460003306489e-20

R51_85 V51 V85 28253.689737215056
L51_85 V51 V85 5.0536799034445256e-11
C51_85 V51 V85 -8.660583331177545e-21

R51_86 V51 V86 10016.925770051444
L51_86 V51 V86 1.2954903247576785e-11
C51_86 V51 V86 -5.01311637942115e-20

R51_87 V51 V87 1512.5907965847982
L51_87 V51 V87 -5.938500760587731e-12
C51_87 V51 V87 -2.040058480362517e-19

R51_88 V51 V88 5752.522537708226
L51_88 V51 V88 -1.5623139638361967e-09
C51_88 V51 V88 4.24024407078472e-20

R51_89 V51 V89 7538.101370471845
L51_89 V51 V89 -9.230687738693442e-12
C51_89 V51 V89 -3.038321902118306e-20

R51_90 V51 V90 -12168.430233313897
L51_90 V51 V90 -4.604822249230509e-12
C51_90 V51 V90 -6.171479104424708e-20

R51_91 V51 V91 -580.9231831426894
L51_91 V51 V91 1.6521209563870633e-11
C51_91 V51 V91 1.1914201779200553e-19

R51_92 V51 V92 -4238.256017797616
L51_92 V51 V92 4.28562134792873e-11
C51_92 V51 V92 -2.4994868202557894e-20

R51_93 V51 V93 -12272.47334668772
L51_93 V51 V93 -5.568554405746076e-11
C51_93 V51 V93 2.6189754479901843e-20

R51_94 V51 V94 -365886.511562783
L51_94 V51 V94 5.379740939135505e-12
C51_94 V51 V94 1.2394766701150648e-19

R51_95 V51 V95 3254.569476432483
L51_95 V51 V95 2.6605744822827457e-12
C51_95 V51 V95 1.3032020604298407e-19

R51_96 V51 V96 -740335.5787312058
L51_96 V51 V96 -1.3912136424248167e-11
C51_96 V51 V96 1.518926627384082e-20

R51_97 V51 V97 6052.602402118395
L51_97 V51 V97 5.278348092652597e-12
C51_97 V51 V97 8.831705081483574e-20

R51_98 V51 V98 -18185.501461234868
L51_98 V51 V98 1.1126472665607343e-10
C51_98 V51 V98 -1.94456299593327e-20

R51_99 V51 V99 612.6440785187932
L51_99 V51 V99 -2.2563580909338755e-12
C51_99 V51 V99 -2.6009352745793503e-19

R51_100 V51 V100 4216.027082084239
L51_100 V51 V100 5.343415589183846e-12
C51_100 V51 V100 7.308431794153389e-20

R51_101 V51 V101 -2706.4369013459695
L51_101 V51 V101 -5.048513474612673e-12
C51_101 V51 V101 -1.16839009964644e-19

R51_102 V51 V102 6634.531719766782
L51_102 V51 V102 -4.4558679733486794e-12
C51_102 V51 V102 -1.5110711925643521e-19

R51_103 V51 V103 -974.4054278614668
L51_103 V51 V103 5.16458947178601e-10
C51_103 V51 V103 9.961477534115391e-20

R51_104 V51 V104 -19524.715523114646
L51_104 V51 V104 1.978578645949825e-11
C51_104 V51 V104 -8.794140415180813e-20

R51_105 V51 V105 4306.385713249117
L51_105 V51 V105 -4.975691168065891e-12
C51_105 V51 V105 -3.5281246515624984e-20

R51_106 V51 V106 12927.615262583977
L51_106 V51 V106 5.514186007252177e-12
C51_106 V51 V106 1.4228208570816385e-19

R51_107 V51 V107 -1024.688411607702
L51_107 V51 V107 2.417283093170801e-12
C51_107 V51 V107 6.366084077789153e-20

R51_108 V51 V108 -4848.001397383211
L51_108 V51 V108 -3.248154586570454e-12
C51_108 V51 V108 2.6306878699637464e-22

R51_109 V51 V109 2346.0330715162627
L51_109 V51 V109 1.1305146077929662e-11
C51_109 V51 V109 5.548460848381008e-20

R51_110 V51 V110 -8487.65298254385
L51_110 V51 V110 -1.1104865895211969e-10
C51_110 V51 V110 2.8728598696372815e-20

R51_111 V51 V111 1287.9041650448746
L51_111 V51 V111 -2.1040427101287393e-12
C51_111 V51 V111 -7.341640397461483e-20

R51_112 V51 V112 40271.56491863038
L51_112 V51 V112 4.63924853446869e-12
C51_112 V51 V112 1.5395627874922155e-20

R51_113 V51 V113 -1278.050208239447
L51_113 V51 V113 1.5377365886930844e-11
C51_113 V51 V113 4.81724212332466e-20

R51_114 V51 V114 -90657.70132494101
L51_114 V51 V114 -1.479480588808016e-11
C51_114 V51 V114 -7.396640133330949e-20

R51_115 V51 V115 957.8142216393746
L51_115 V51 V115 1.17161138179763e-11
C51_115 V51 V115 -7.370222880816063e-21

R51_116 V51 V116 2755.0997728395946
L51_116 V51 V116 1.4761062416444226e-11
C51_116 V51 V116 2.9169070736491623e-22

R51_117 V51 V117 -42917.15836006848
L51_117 V51 V117 7.979338827616194e-12
C51_117 V51 V117 1.77256939617866e-20

R51_118 V51 V118 15621.245428050459
L51_118 V51 V118 2.0855705546203584e-11
C51_118 V51 V118 -3.874215198410555e-20

R51_119 V51 V119 -615.2838640380727
L51_119 V51 V119 1.0756680641071524e-12
C51_119 V51 V119 4.4612550159891284e-20

R51_120 V51 V120 -2277.808459268967
L51_120 V51 V120 -4.117338683133475e-12
C51_120 V51 V120 3.605709891123393e-20

R51_121 V51 V121 1649.0539936604252
L51_121 V51 V121 -3.2395773343878035e-12
C51_121 V51 V121 -1.4883657037583308e-19

R51_122 V51 V122 13143.74455499154
L51_122 V51 V122 2.483816901535453e-11
C51_122 V51 V122 1.0699412587435322e-19

R51_123 V51 V123 1795.5669448632289
L51_123 V51 V123 -9.662055171971199e-13
C51_123 V51 V123 -4.1215532956991224e-20

R51_124 V51 V124 24243.409785387437
L51_124 V51 V124 3.654928831903527e-12
C51_124 V51 V124 -8.272285661629408e-20

R51_125 V51 V125 -6204.821793712114
L51_125 V51 V125 -5.820875252870022e-12
C51_125 V51 V125 6.725171243509333e-21

R51_126 V51 V126 -2619.2381163568407
L51_126 V51 V126 -4.61203609817276e-12
C51_126 V51 V126 -1.2664716420866582e-20

R51_127 V51 V127 2463.2631112205377
L51_127 V51 V127 -2.5329745937609083e-12
C51_127 V51 V127 5.39777483227846e-20

R51_128 V51 V128 2842.6526038862103
L51_128 V51 V128 -5.070671304591549e-12
C51_128 V51 V128 2.2317100526970952e-20

R51_129 V51 V129 -4700.792612691913
L51_129 V51 V129 4.633612344027993e-12
C51_129 V51 V129 1.7414062931916927e-19

R51_130 V51 V130 3785.545487187793
L51_130 V51 V130 1.2712887394940443e-11
C51_130 V51 V130 -7.698314500102373e-20

R51_131 V51 V131 -3004.79737532733
L51_131 V51 V131 1.0059314371195153e-12
C51_131 V51 V131 -6.083626234378463e-20

R51_132 V51 V132 -2072.5787416872868
L51_132 V51 V132 2.9598249666036893e-12
C51_132 V51 V132 1.1137789004755715e-20

R51_133 V51 V133 -5277.201631181844
L51_133 V51 V133 1.1769663289655982e-11
C51_133 V51 V133 -8.454899372983647e-20

R51_134 V51 V134 -15923.264037383846
L51_134 V51 V134 2.8428947128490845e-12
C51_134 V51 V134 1.7852736180982858e-19

R51_135 V51 V135 682.2124303781849
L51_135 V51 V135 -1.3208082399771471e-12
C51_135 V51 V135 -2.8326174205849386e-20

R51_136 V51 V136 7081.236137040725
L51_136 V51 V136 2.236663115142038e-12
C51_136 V51 V136 -4.1221733322479576e-20

R51_137 V51 V137 2273.061263864502
L51_137 V51 V137 -6.983980657722119e-12
C51_137 V51 V137 -9.994673738953438e-20

R51_138 V51 V138 14889.70560623628
L51_138 V51 V138 -2.331187761386483e-12
C51_138 V51 V138 -1.0541523461601383e-19

R51_139 V51 V139 -437.5947998424123
L51_139 V51 V139 1.9297137847287244e-12
C51_139 V51 V139 8.257360042986884e-20

R51_140 V51 V140 -4213.493179695389
L51_140 V51 V140 -1.130072135754733e-12
C51_140 V51 V140 5.3125664828762983e-20

R51_141 V51 V141 3692.3694301812293
L51_141 V51 V141 3.488704451424458e-11
C51_141 V51 V141 1.401987297214162e-19

R51_142 V51 V142 -19520.7148711883
L51_142 V51 V142 -2.934982596626177e-12
C51_142 V51 V142 -4.157055634608469e-20

R51_143 V51 V143 -1956.830656616062
L51_143 V51 V143 1.888501663087002e-12
C51_143 V51 V143 2.7968151874426384e-20

R51_144 V51 V144 -2378.543687082758
L51_144 V51 V144 6.526804805230591e-12
C51_144 V51 V144 2.4047436552308904e-20

R51_145 V51 V145 -1974.94552116203
L51_145 V51 V145 6.25299367171313e-11
C51_145 V51 V145 5.1065011075706793e-20

R51_146 V51 V146 -5577.681216238925
L51_146 V51 V146 1.2998085816578995e-12
C51_146 V51 V146 3.413148621306309e-20

R51_147 V51 V147 290.5096765051888
L51_147 V51 V147 -1.032378946412927e-12
C51_147 V51 V147 -5.443770220025241e-20

R51_148 V51 V148 1594.428144833233
L51_148 V51 V148 1.420573127720225e-12
C51_148 V51 V148 -3.51842257527381e-20

R51_149 V51 V149 -2919.2193410356253
L51_149 V51 V149 -2.8321339551344896e-12
C51_149 V51 V149 -2.6667622188257503e-19

R51_150 V51 V150 4567.9005023009895
L51_150 V51 V150 -9.761542649142233e-11
C51_150 V51 V150 1.1743628170514222e-19

R51_151 V51 V151 -575.026902697245
L51_151 V51 V151 -1.9561126903528253e-12
C51_151 V51 V151 -2.5105091696408984e-20

R51_152 V51 V152 -4023.986350677183
L51_152 V51 V152 -4.398047558174121e-12
C51_152 V51 V152 1.3758281745319276e-20

R51_153 V51 V153 2116.2207930215063
L51_153 V51 V153 6.57560556690286e-12
C51_153 V51 V153 2.5626163428733173e-20

R51_154 V51 V154 -58311.17037507377
L51_154 V51 V154 -3.334597301962708e-12
C51_154 V51 V154 -1.1057851927987366e-19

R51_155 V51 V155 588.9454553005222
L51_155 V51 V155 1.0254707754525984e-12
C51_155 V51 V155 -4.405252812987388e-20

R51_156 V51 V156 6583.0138479486595
L51_156 V51 V156 -2.7682792215511176e-12
C51_156 V51 V156 -3.612757713610411e-21

R51_157 V51 V157 2134.87639010553
L51_157 V51 V157 2.9129496896267462e-12
C51_157 V51 V157 2.653577490788488e-19

R51_158 V51 V158 -4252.174453459724
L51_158 V51 V158 -1.3051720385540682e-11
C51_158 V51 V158 -1.707709635780073e-21

R51_159 V51 V159 -1051.6982717854467
L51_159 V51 V159 2.8998257402955758e-12
C51_159 V51 V159 2.230373047282223e-21

R51_160 V51 V160 -10260.987472687038
L51_160 V51 V160 6.9470682334886114e-12
C51_160 V51 V160 -2.9242552534522146e-20

R51_161 V51 V161 -2811.197067268816
L51_161 V51 V161 -2.489400757326799e-12
C51_161 V51 V161 -6.194918875580276e-20

R51_162 V51 V162 -6730.646670210828
L51_162 V51 V162 1.0793281951347809e-11
C51_162 V51 V162 5.608359182352711e-21

R51_163 V51 V163 -17732.588181698597
L51_163 V51 V163 -1.1230317908397108e-12
C51_163 V51 V163 6.279336126718904e-20

R51_164 V51 V164 -2213.2517201041346
L51_164 V51 V164 4.7272928265815756e-11
C51_164 V51 V164 1.33571763288472e-20

R51_165 V51 V165 -3022.2785482415793
L51_165 V51 V165 -2.8594019836515204e-12
C51_165 V51 V165 -1.7290434591036638e-19

R51_166 V51 V166 1892.1927652980391
L51_166 V51 V166 -4.20073427295929e-12
C51_166 V51 V166 -1.146288428979328e-20

R51_167 V51 V167 -1230.967222131492
L51_167 V51 V167 1.8073904758705035e-12
C51_167 V51 V167 -1.3683284356444797e-21

R51_168 V51 V168 3529.5717039411957
L51_168 V51 V168 -3.5392712921447682e-12
C51_168 V51 V168 3.977959702532263e-20

R51_169 V51 V169 2759.4491682983917
L51_169 V51 V169 2.645647356252288e-12
C51_169 V51 V169 6.6520322084852466e-21

R51_170 V51 V170 -3529.6132546099393
L51_170 V51 V170 9.156401124517485e-12
C51_170 V51 V170 -9.260562482360196e-20

R51_171 V51 V171 661.1367735347026
L51_171 V51 V171 -3.461385053697815e-12
C51_171 V51 V171 -1.7446376880202577e-19

R51_172 V51 V172 3970.667655130067
L51_172 V51 V172 6.485896043170552e-12
C51_172 V51 V172 -8.410050272905612e-20

R51_173 V51 V173 2917.9904509987327
L51_173 V51 V173 1.651567943523345e-11
C51_173 V51 V173 1.3982210777864177e-19

R51_174 V51 V174 -10813.680951631677
L51_174 V51 V174 2.758870751070409e-12
C51_174 V51 V174 1.110047853370812e-19

R51_175 V51 V175 -2938.14152607704
L51_175 V51 V175 2.754909793873901e-10
C51_175 V51 V175 6.917720967352751e-20

R51_176 V51 V176 11718.613250623568
L51_176 V51 V176 6.56985776443114e-12
C51_176 V51 V176 5.593695264529491e-20

R51_177 V51 V177 -1083.4950188580474
L51_177 V51 V177 -4.4321078589226185e-12
C51_177 V51 V177 -8.22544007862699e-20

R51_178 V51 V178 17606.202216360056
L51_178 V51 V178 -2.9626576199821524e-12
C51_178 V51 V178 5.050593709029827e-20

R51_179 V51 V179 15937.211170828032
L51_179 V51 V179 2.0941526772884338e-12
C51_179 V51 V179 9.234722220773675e-20

R51_180 V51 V180 -2881.194279848817
L51_180 V51 V180 -6.7648363212098015e-12
C51_180 V51 V180 6.340149789828478e-20

R51_181 V51 V181 2286.8670044762653
L51_181 V51 V181 1.3177247024563655e-11
C51_181 V51 V181 -2.2788300310261164e-20

R51_182 V51 V182 1843.9595846295138
L51_182 V51 V182 -1.5165498237184913e-11
C51_182 V51 V182 -9.778578532300124e-20

R51_183 V51 V183 -1261.5766607212145
L51_183 V51 V183 -4.812362776896497e-12
C51_183 V51 V183 2.5803377227420907e-20

R51_184 V51 V184 -5011.478286685172
L51_184 V51 V184 2.0889334222238914e-11
C51_184 V51 V184 -1.4839983934365115e-20

R51_185 V51 V185 1504.4173936686816
L51_185 V51 V185 9.592050044756853e-12
C51_185 V51 V185 4.8753216499875083e-20

R51_186 V51 V186 -3642.0527183971058
L51_186 V51 V186 7.559956050653674e-12
C51_186 V51 V186 -4.271447387154283e-20

R51_187 V51 V187 1492.088879969799
L51_187 V51 V187 -4.254405008756593e-12
C51_187 V51 V187 -7.343849036854357e-20

R51_188 V51 V188 1796.6877392534134
L51_188 V51 V188 -4.65635370633997e-12
C51_188 V51 V188 -8.698412042130842e-20

R51_189 V51 V189 -1586.3071541723868
L51_189 V51 V189 -1.2683197380284563e-11
C51_189 V51 V189 -9.312552913940654e-20

R51_190 V51 V190 -5215.611799368931
L51_190 V51 V190 -8.936366257148553e-12
C51_190 V51 V190 8.86424097262915e-20

R51_191 V51 V191 1614.838672383573
L51_191 V51 V191 -2.0097861783372084e-11
C51_191 V51 V191 -1.0873652782791035e-19

R51_192 V51 V192 3435.077735777905
L51_192 V51 V192 9.559185490555546e-12
C51_192 V51 V192 -5.48620758903893e-20

R51_193 V51 V193 -4020.1855224108094
L51_193 V51 V193 -9.117744415297906e-12
C51_193 V51 V193 8.064006467005514e-20

R51_194 V51 V194 1820.4422068336758
L51_194 V51 V194 4.235961184053861e-12
C51_194 V51 V194 1.3808815800600514e-21

R51_195 V51 V195 -1284.1801771516975
L51_195 V51 V195 1.8379888051055668e-12
C51_195 V51 V195 1.6773671415794913e-19

R51_196 V51 V196 -1185.245130090165
L51_196 V51 V196 7.522949519458934e-12
C51_196 V51 V196 1.989578358385792e-19

R51_197 V51 V197 5037.206984782135
L51_197 V51 V197 8.095375824712377e-12
C51_197 V51 V197 2.5941684425520165e-20

R51_198 V51 V198 -12152.829732330592
L51_198 V51 V198 1.5791142043381783e-11
C51_198 V51 V198 -3.433767583108457e-20

R51_199 V51 V199 17903.43637292092
L51_199 V51 V199 -4.10627829355154e-12
C51_199 V51 V199 2.8868830157315955e-20

R51_200 V51 V200 -5987.75779251399
L51_200 V51 V200 -1.1243592444871933e-11
C51_200 V51 V200 5.9163404734526784e-21

R52_52 V52 0 -781.7946445149809
L52_52 V52 0 -5.546862559251846e-12
C52_52 V52 0 -1.5473841875216134e-18

R52_53 V52 V53 17133.559947683072
L52_53 V52 V53 4.264304866296931e-12
C52_53 V52 V53 1.640421681860393e-19

R52_54 V52 V54 -32035.511017885347
L52_54 V52 V54 3.29465036341427e-12
C52_54 V52 V54 1.5182589173748807e-19

R52_55 V52 V55 29776.820971737372
L52_55 V52 V55 2.9882283957217277e-12
C52_55 V52 V55 1.98011124517129e-19

R52_56 V52 V56 3191.8729495332345
L52_56 V52 V56 7.083931998675105e-12
C52_56 V52 V56 1.598142734864312e-20

R52_57 V52 V57 -129379.03362138505
L52_57 V52 V57 1.4224065175067336e-11
C52_57 V52 V57 7.07665857612131e-20

R52_58 V52 V58 55955.64564428518
L52_58 V52 V58 -1.602805321562665e-11
C52_58 V52 V58 7.571944281222844e-21

R52_59 V52 V59 9223.615470463585
L52_59 V52 V59 4.121911325784276e-12
C52_59 V52 V59 2.1903564157415163e-19

R52_60 V52 V60 2121.1666831787247
L52_60 V52 V60 6.93851005338228e-13
C52_60 V52 V60 1.0863880119255854e-18

R52_61 V52 V61 67932.13758513791
L52_61 V52 V61 -3.577670245199551e-12
C52_61 V52 V61 -1.603199764003056e-19

R52_62 V52 V62 24888.46936801825
L52_62 V52 V62 1.5918161826778057e-10
C52_62 V52 V62 7.25926167298783e-20

R52_63 V52 V63 -14931.565272682223
L52_63 V52 V63 -3.5946631295959424e-12
C52_63 V52 V63 -2.00180572341976e-19

R52_64 V52 V64 -3335.3657911255864
L52_64 V52 V64 -1.1823510097161324e-12
C52_64 V52 V64 -7.463267968422356e-19

R52_65 V52 V65 4729.78952482973
L52_65 V52 V65 6.3208358646269604e-12
C52_65 V52 V65 1.435035128398518e-19

R52_66 V52 V66 -140882.58601323905
L52_66 V52 V66 6.3799850512985e-12
C52_66 V52 V66 1.0212711826974762e-19

R52_67 V52 V67 -14569.69732250154
L52_67 V52 V67 1.7442171112814937e-11
C52_67 V52 V67 -4.950131560433739e-20

R52_68 V52 V68 -2219.6189306895244
L52_68 V52 V68 -1.9966898794357556e-12
C52_68 V52 V68 -2.820698439866453e-19

R52_69 V52 V69 -6307.10412735494
L52_69 V52 V69 1.3852808466256589e-11
C52_69 V52 V69 5.2698418534759746e-21

R52_70 V52 V70 31303.693933348273
L52_70 V52 V70 -3.3821765285403428e-12
C52_70 V52 V70 -2.6845205807769e-19

R52_71 V52 V71 10972.084288826807
L52_71 V52 V71 1.9670670964527408e-10
C52_71 V52 V71 6.280497537848538e-20

R52_72 V52 V72 2954.991555682145
L52_72 V52 V72 1.270415281194812e-12
C52_72 V52 V72 7.053766815778379e-19

R52_73 V52 V73 7429.956092832265
L52_73 V52 V73 -1.28698678062638e-11
C52_73 V52 V73 -6.4546823714227004e-21

R52_74 V52 V74 13138.728548971701
L52_74 V52 V74 1.5518549653914138e-11
C52_74 V52 V74 1.1367134734496832e-19

R52_75 V52 V75 7892.663273984637
L52_75 V52 V75 6.093020844722688e-12
C52_75 V52 V75 1.355257339268219e-19

R52_76 V52 V76 1743.9854524402892
L52_76 V52 V76 -1.2016972449572055e-11
C52_76 V52 V76 -3.8058808467489177e-19

R52_77 V52 V77 3025.1633536022696
L52_77 V52 V77 7.285522968473535e-11
C52_77 V52 V77 8.474223473697769e-20

R52_78 V52 V78 -9331.931076829656
L52_78 V52 V78 1.982134495529896e-11
C52_78 V52 V78 8.184258664058202e-20

R52_79 V52 V79 -5056.484666516842
L52_79 V52 V79 -5.223416961540851e-11
C52_79 V52 V79 -2.728778953366566e-20

R52_80 V52 V80 -848.9008975023689
L52_80 V52 V80 -1.855587616377308e-12
C52_80 V52 V80 -1.6892036184542542e-19

R52_81 V52 V81 -2973.2841202845248
L52_81 V52 V81 -1.055654717308554e-11
C52_81 V52 V81 1.0299391699762962e-21

R52_82 V52 V82 27249.308191515673
L52_82 V52 V82 2.0018842755150206e-11
C52_82 V52 V82 5.48649284618142e-20

R52_83 V52 V83 -24565.92212690307
L52_83 V52 V83 -5.461304933337999e-11
C52_83 V52 V83 -3.978383178083996e-20

R52_84 V52 V84 5125.610740733633
L52_84 V52 V84 2.032832546126503e-12
C52_84 V52 V84 4.1934166034916777e-19

R52_85 V52 V85 67220.74885596715
L52_85 V52 V85 1.312251005135736e-11
C52_85 V52 V85 4.4235138098069156e-20

R52_86 V52 V86 3773.2801578309673
L52_86 V52 V86 8.430938079706359e-12
C52_86 V52 V86 1.869131303018737e-20

R52_87 V52 V87 2120.5566076354476
L52_87 V52 V87 2.066540509337247e-11
C52_87 V52 V87 -4.6088727804045814e-20

R52_88 V52 V88 743.3133458905936
L52_88 V52 V88 -4.504483677713709e-12
C52_88 V52 V88 -3.507853185069348e-19

R52_89 V52 V89 2650.336921673883
L52_89 V52 V89 -1.3854879410495525e-11
C52_89 V52 V89 -1.1670611142554883e-19

R52_90 V52 V90 -14723.130762390158
L52_90 V52 V90 -3.5365727331548712e-12
C52_90 V52 V90 -2.426165789171067e-19

R52_91 V52 V91 -1753.8671984682674
L52_91 V52 V91 6.111265062337565e-12
C52_91 V52 V91 1.8200705716638038e-19

R52_92 V52 V92 -400.81622563741456
L52_92 V52 V92 2.190310866212961e-11
C52_92 V52 V92 1.8290487657288383e-19

R52_93 V52 V93 18937.73434639644
L52_93 V52 V93 -9.186031068061811e-12
C52_93 V52 V93 -7.23700731230869e-21

R52_94 V52 V94 15909.213391323667
L52_94 V52 V94 3.834116144611844e-12
C52_94 V52 V94 2.0613019786063802e-19

R52_95 V52 V95 -3424.9127822206265
L52_95 V52 V95 -2.7196787952754966e-11
C52_95 V52 V95 3.262189855402594e-20

R52_96 V52 V96 -11410.997229479222
L52_96 V52 V96 2.1769731558732356e-12
C52_96 V52 V96 1.9933669244052263e-19

R52_97 V52 V97 -76364.36773805489
L52_97 V52 V97 3.664831228618867e-12
C52_97 V52 V97 3.1157233936931626e-19

R52_98 V52 V98 -4188.210646618508
L52_98 V52 V98 1.6556659316527853e-11
C52_98 V52 V98 1.3654613459435566e-19

R52_99 V52 V99 1265.4279108390826
L52_99 V52 V99 -2.0186384778864153e-11
C52_99 V52 V99 -1.9330744860226977e-19

R52_100 V52 V100 389.9377061954125
L52_100 V52 V100 -1.865126049780361e-12
C52_100 V52 V100 -4.397723738204336e-19

R52_101 V52 V101 -2628.027955963943
L52_101 V52 V101 -6.018067174428028e-12
C52_101 V52 V101 -1.9077483882760904e-19

R52_102 V52 V102 10912.641389419503
L52_102 V52 V102 -2.6723437323605754e-12
C52_102 V52 V102 -2.9736883360305844e-19

R52_103 V52 V103 -10957.81754576465
L52_103 V52 V103 7.146103762518078e-11
C52_103 V52 V103 -1.3268057234136164e-20

R52_104 V52 V104 -1056.4532923972488
L52_104 V52 V104 7.0941575647667685e-12
C52_104 V52 V104 2.525803923991214e-19

R52_105 V52 V105 1380.2622257176802
L52_105 V52 V105 -4.369117953208082e-12
C52_105 V52 V105 -8.406190832842605e-20

R52_106 V52 V106 1500.660567429764
L52_106 V52 V106 5.726297070196658e-12
C52_106 V52 V106 6.915856915401727e-20

R52_107 V52 V107 -1907.9523018468847
L52_107 V52 V107 9.042054904724368e-12
C52_107 V52 V107 1.933171855975985e-19

R52_108 V52 V108 -545.7209143140543
L52_108 V52 V108 3.9330052105713045e-12
C52_108 V52 V108 -3.183496994495036e-20

R52_109 V52 V109 2263.8128544908127
L52_109 V52 V109 3.667596969703741e-12
C52_109 V52 V109 1.9762944104900893e-19

R52_110 V52 V110 -1470.1743956916584
L52_110 V52 V110 8.99912185882383e-12
C52_110 V52 V110 1.1866653428504294e-19

R52_111 V52 V111 2077.2937636158194
L52_111 V52 V111 1.9748927184393578e-11
C52_111 V52 V111 -3.084248746559258e-20

R52_112 V52 V112 631.9276560207863
L52_112 V52 V112 -2.9583170722652264e-12
C52_112 V52 V112 -9.601661413196486e-21

R52_113 V52 V113 -777.9726298145825
L52_113 V52 V113 -1.6336668945240613e-11
C52_113 V52 V113 3.326622254011542e-20

R52_114 V52 V114 -2616.1704804132523
L52_114 V52 V114 -5.673210194630827e-12
C52_114 V52 V114 -4.810173545260718e-21

R52_115 V52 V115 20223.41100098526
L52_115 V52 V115 -5.075939628110617e-12
C52_115 V52 V115 -1.5103072902092039e-19

R52_116 V52 V116 734.2543508070261
L52_116 V52 V116 -2.4100266824182173e-09
C52_116 V52 V116 3.5234032456529844e-20

R52_117 V52 V117 -45153.73987810026
L52_117 V52 V117 4.836862295382021e-11
C52_117 V52 V117 -1.3576244287131553e-20

R52_118 V52 V118 1048.8766762519788
L52_118 V52 V118 -1.092989746986999e-11
C52_118 V52 V118 -1.9486378258468022e-19

R52_119 V52 V119 -2500.287419611943
L52_119 V52 V119 -5.1173260214569446e-11
C52_119 V52 V119 1.6406717013360926e-20

R52_120 V52 V120 -347.6301264325539
L52_120 V52 V120 1.7239479543930799e-12
C52_120 V52 V120 -1.252721500949229e-19

R52_121 V52 V121 1143.6170908291315
L52_121 V52 V121 -6.691874195701523e-12
C52_121 V52 V121 -1.5296862212425926e-19

R52_122 V52 V122 -3521.8656267963906
L52_122 V52 V122 5.086688614010812e-12
C52_122 V52 V122 1.2423508414064468e-19

R52_123 V52 V123 3021.5555790855674
L52_123 V52 V123 6.072387145779783e-12
C52_123 V52 V123 4.627004737334927e-20

R52_124 V52 V124 591.8917465973874
L52_124 V52 V124 -1.5920705447759817e-12
C52_124 V52 V124 1.7716526199391554e-19

R52_125 V52 V125 13315.58444303267
L52_125 V52 V125 -7.339276876721548e-12
C52_125 V52 V125 9.695846391965868e-21

R52_126 V52 V126 -1005.9219961121827
L52_126 V52 V126 -7.505125199149037e-12
C52_126 V52 V126 9.459315122749948e-20

R52_127 V52 V127 -2205.6307015466714
L52_127 V52 V127 -1.0088490456655673e-11
C52_127 V52 V127 4.1730819517726966e-20

R52_128 V52 V128 1807.5850037002892
L52_128 V52 V128 -2.7754742366160627e-12
C52_128 V52 V128 -1.508311275142488e-21

R52_129 V52 V129 -1745.596177821112
L52_129 V52 V129 3.4658719468340894e-12
C52_129 V52 V129 3.1833194256564847e-19

R52_130 V52 V130 1983.3477114957013
L52_130 V52 V130 -6.872587331637549e-12
C52_130 V52 V130 -2.151516012000716e-19

R52_131 V52 V131 4414.925255622015
L52_131 V52 V131 1.071798221631178e-11
C52_131 V52 V131 -7.500105179753959e-20

R52_132 V52 V132 -1063.1088558764122
L52_132 V52 V132 9.214240815367625e-13
C52_132 V52 V132 -1.0805322775742085e-19

R52_133 V52 V133 -1326.2741550652563
L52_133 V52 V133 -1.9113615031503993e-11
C52_133 V52 V133 -2.4012958527213566e-19

R52_134 V52 V134 -5157.017594610781
L52_134 V52 V134 2.7859050792428115e-12
C52_134 V52 V134 1.6442575926289254e-19

R52_135 V52 V135 1785.8201931410213
L52_135 V52 V135 9.163243471597176e-12
C52_135 V52 V135 -1.6484300381531458e-20

R52_136 V52 V136 450.3130400192796
L52_136 V52 V136 -2.565987792315302e-12
C52_136 V52 V136 1.1335520634363068e-19

R52_137 V52 V137 710.3409485090892
L52_137 V52 V137 -2.4611895820468757e-12
C52_137 V52 V137 -1.5081823031090232e-19

R52_138 V52 V138 9311.602205053465
L52_138 V52 V138 -2.926903902647687e-12
C52_138 V52 V138 -5.24697325017268e-20

R52_139 V52 V139 -978.991454155152
L52_139 V52 V139 -1.7425714052492348e-12
C52_139 V52 V139 -6.927912014772935e-20

R52_140 V52 V140 -287.0424179363424
L52_140 V52 V140 -2.3413141379320224e-12
C52_140 V52 V140 -9.336167875469729e-20

R52_141 V52 V141 1676.2880685071411
L52_141 V52 V141 3.2150129515186714e-12
C52_141 V52 V141 3.2010125056952984e-19

R52_142 V52 V142 -1850.383555695281
L52_142 V52 V142 -2.6290078286640323e-12
C52_142 V52 V142 -5.617591475611315e-20

R52_143 V52 V143 -13329.469390025048
L52_143 V52 V143 3.4610894637391216e-12
C52_143 V52 V143 1.199484888959796e-19

R52_144 V52 V144 22039.065741665865
L52_144 V52 V144 1.3630555051360275e-12
C52_144 V52 V144 3.0030548945884253e-20

R52_145 V52 V145 -662.8422573253821
L52_145 V52 V145 2.93641113152762e-12
C52_145 V52 V145 8.566389035200676e-20

R52_146 V52 V146 3146.4823692195127
L52_146 V52 V146 1.022821821858071e-12
C52_146 V52 V146 4.572181005890986e-21

R52_147 V52 V147 1288.7072022016227
L52_147 V52 V147 2.8087391762712844e-12
C52_147 V52 V147 5.010474208330903e-20

R52_148 V52 V148 464.6203993293884
L52_148 V52 V148 -1.1797239412558416e-12
C52_148 V52 V148 7.739752892761601e-21

R52_149 V52 V149 -2900.6370841435187
L52_149 V52 V149 -1.06951143474666e-12
C52_149 V52 V149 -4.529926208346726e-19

R52_150 V52 V150 837.8100457821034
L52_150 V52 V150 -5.39993537159259e-12
C52_150 V52 V150 2.9215073111275863e-19

R52_151 V52 V151 1585.1384296552246
L52_151 V52 V151 -5.687122569741495e-12
C52_151 V52 V151 -8.901996526495381e-20

R52_152 V52 V152 1465.428346818961
L52_152 V52 V152 -1.9809705643064947e-12
C52_152 V52 V152 4.829936867944355e-20

R52_153 V52 V153 785.4643727429532
L52_153 V52 V153 1.0866546907257976e-11
C52_153 V52 V153 3.046317784192778e-20

R52_154 V52 V154 13376.70911242137
L52_154 V52 V154 -3.874308252811407e-12
C52_154 V52 V154 -1.8232620927329554e-19

R52_155 V52 V155 -1073.413870340209
L52_155 V52 V155 -3.742844508680179e-12
C52_155 V52 V155 -9.308934578930695e-20

R52_156 V52 V156 -391.9384194834439
L52_156 V52 V156 1.1251310436327175e-12
C52_156 V52 V156 -6.463367859595307e-20

R52_157 V52 V157 1947.8442299545657
L52_157 V52 V157 1.3978992957499328e-12
C52_157 V52 V157 5.056002514949188e-19

R52_158 V52 V158 -1583.6973831274058
L52_158 V52 V158 -6.32582390293734e-12
C52_158 V52 V158 -6.679778655446112e-21

R52_159 V52 V159 7623.304241136558
L52_159 V52 V159 4.049831715248029e-12
C52_159 V52 V159 3.952370861538948e-20

R52_160 V52 V160 -10167.575092717954
L52_160 V52 V160 1.5782384135197948e-12
C52_160 V52 V160 -9.601220863836829e-20

R52_161 V52 V161 -2277.8946091708503
L52_161 V52 V161 -3.705783532624759e-12
C52_161 V52 V161 -8.563818604608777e-20

R52_162 V52 V162 -5915.260662531878
L52_162 V52 V162 7.37308684590668e-12
C52_162 V52 V162 -1.0950534166045295e-20

R52_163 V52 V163 -2677.592760157576
L52_163 V52 V163 1.5130473208798936e-11
C52_163 V52 V163 1.011025158921173e-19

R52_164 V52 V164 1538.1705573854836
L52_164 V52 V164 -1.0269800886444583e-12
C52_164 V52 V164 3.4824156946302015e-20

R52_165 V52 V165 -2260.2353105502807
L52_165 V52 V165 -1.872415392865255e-12
C52_165 V52 V165 -2.1019275263183122e-19

R52_166 V52 V166 1079.9363532189143
L52_166 V52 V166 -4.229323806322985e-12
C52_166 V52 V166 6.31650204734806e-20

R52_167 V52 V167 3137.51109742818
L52_167 V52 V167 -8.306431299793909e-12
C52_167 V52 V167 1.2502024438290312e-20

R52_168 V52 V168 -1474.513006700452
L52_168 V52 V168 2.2580066137660375e-12
C52_168 V52 V168 3.3322651341359504e-20

R52_169 V52 V169 950.6602818126344
L52_169 V52 V169 2.1528732748845358e-12
C52_169 V52 V169 8.55927917922428e-20

R52_170 V52 V170 29966.544935331567
L52_170 V52 V170 3.904519900433677e-12
C52_170 V52 V170 -1.3453565332272538e-19

R52_171 V52 V171 2115.5507701678707
L52_171 V52 V171 -1.3021307398939075e-10
C52_171 V52 V171 -1.923744849351427e-19

R52_172 V52 V172 -7498.854559506333
L52_172 V52 V172 -4.38241062290442e-12
C52_172 V52 V172 -1.2802196205521582e-19

R52_173 V52 V173 6199.223702713925
L52_173 V52 V173 1.8888280522914313e-10
C52_173 V52 V173 9.766606074840704e-20

R52_174 V52 V174 -922.1160134023174
L52_174 V52 V174 5.044396613611616e-12
C52_174 V52 V174 1.5665394949166406e-19

R52_175 V52 V175 -2444.49955735396
L52_175 V52 V175 -2.188697628624087e-11
C52_175 V52 V175 -2.3180484668227035e-20

R52_176 V52 V176 1462.551579146667
L52_176 V52 V176 1.5752221007217383e-11
C52_176 V52 V176 1.0148268039745497e-20

R52_177 V52 V177 -1188.2824251448974
L52_177 V52 V177 -3.799424253205296e-12
C52_177 V52 V177 -5.593338741857747e-20

R52_178 V52 V178 1853.586726023379
L52_178 V52 V178 -2.6806629771777595e-12
C52_178 V52 V178 7.451745932165294e-20

R52_179 V52 V179 -4057.2376112242528
L52_179 V52 V179 2.0701940395864358e-11
C52_179 V52 V179 2.282052268931589e-19

R52_180 V52 V180 -1035.841640863535
L52_180 V52 V180 2.0855100627125463e-12
C52_180 V52 V180 1.2328959549015005e-19

R52_181 V52 V181 3340.2265089232937
L52_181 V52 V181 1.747998437535491e-11
C52_181 V52 V181 5.271723632426771e-21

R52_182 V52 V182 1551.5850872025455
L52_182 V52 V182 -4.3180576299783e-12
C52_182 V52 V182 -1.588196138522183e-19

R52_183 V52 V183 -13914.3998430152
L52_183 V52 V183 6.253198224985339e-12
C52_183 V52 V183 2.6567032877644177e-20

R52_184 V52 V184 -2925.901461919164
L52_184 V52 V184 -8.80362797341307e-12
C52_184 V52 V184 7.7098160774124555e-22

R52_185 V52 V185 1150.2269577627246
L52_185 V52 V185 4.07633588242314e-12
C52_185 V52 V185 1.588768450253095e-20

R52_186 V52 V186 -884.7861758817244
L52_186 V52 V186 3.6748159529881625e-12
C52_186 V52 V186 3.8663393534219755e-21

R52_187 V52 V187 -1813.9982441866455
L52_187 V52 V187 -6.786701145072885e-12
C52_187 V52 V187 -1.9187831126665397e-19

R52_188 V52 V188 511.2789303322336
L52_188 V52 V188 -1.7990050778901899e-12
C52_188 V52 V188 -1.9180974599804711e-19

R52_189 V52 V189 -1680.6094347427436
L52_189 V52 V189 -5.267117170725387e-12
C52_189 V52 V189 -1.1026068724065146e-19

R52_190 V52 V190 10754.927277610084
L52_190 V52 V190 -8.10724844898601e-12
C52_190 V52 V190 1.6474083053414642e-19

R52_191 V52 V191 932.712870700137
L52_191 V52 V191 -4.138776912094203e-12
C52_191 V52 V191 -9.642072343907464e-20

R52_192 V52 V192 -1692.0458892871425
L52_192 V52 V192 1.9732264526369485e-11
C52_192 V52 V192 6.102034182709804e-21

R52_193 V52 V193 -1870.416449179446
L52_193 V52 V193 -3.837815659956025e-12
C52_193 V52 V193 9.510021949915567e-20

R52_194 V52 V194 1523.539237802907
L52_194 V52 V194 8.247165564183203e-12
C52_194 V52 V194 9.192765185072098e-20

R52_195 V52 V195 -2796.9019192551664
L52_195 V52 V195 3.405171372543614e-12
C52_195 V52 V195 2.586349877716423e-19

R52_196 V52 V196 -11559.642888197608
L52_196 V52 V196 1.0346778101277071e-12
C52_196 V52 V196 1.6122923917316767e-19

R52_197 V52 V197 3070.103689508313
L52_197 V52 V197 2.9889897787215204e-12
C52_197 V52 V197 5.806724327343584e-20

R52_198 V52 V198 7299.88355694413
L52_198 V52 V198 9.672500971298439e-12
C52_198 V52 V198 7.282168179070272e-21

R52_199 V52 V199 -2463.800288931725
L52_199 V52 V199 4.582219739270965e-12
C52_199 V52 V199 1.515356020653105e-19

R52_200 V52 V200 -5002.115951932244
L52_200 V52 V200 -1.5243797508806813e-12
C52_200 V52 V200 -8.012861818993365e-20

R53_53 V53 0 202.0364684018012
L53_53 V53 0 1.2767278614107159e-11
C53_53 V53 0 -1.077497060274322e-18

R53_54 V53 V54 -3921.4932445975846
L53_54 V53 V54 -2.8831871845943196e-12
C53_54 V53 V54 -1.7433891431809796e-19

R53_55 V53 V55 -5011.6654876897555
L53_55 V53 V55 -2.9945244453093013e-12
C53_55 V53 V55 -1.593509036808467e-19

R53_56 V53 V56 -4615.268027071167
L53_56 V53 V56 -2.4473534659232272e-12
C53_56 V53 V56 -2.2644585436272787e-19

R53_57 V53 V57 29408.050628740515
L53_57 V53 V57 1.129030743683868e-12
C53_57 V53 V57 2.5076536630403505e-19

R53_58 V53 V58 6969.380704221215
L53_58 V53 V58 -1.1796736373380897e-11
C53_58 V53 V58 -1.0494662725548191e-19

R53_59 V53 V59 3882.180054054835
L53_59 V53 V59 6.916868307095247e-12
C53_59 V53 V59 1.2051003264548794e-20

R53_60 V53 V60 2946.440031413993
L53_60 V53 V60 5.262757153481629e-12
C53_60 V53 V60 -1.7837845366130562e-20

R53_61 V53 V61 4236.138126913599
L53_61 V53 V61 2.4120772549861296e-12
C53_61 V53 V61 3.490827356934935e-19

R53_62 V53 V62 8892.353245898768
L53_62 V53 V62 4.032715940636128e-12
C53_62 V53 V62 1.353665668729009e-19

R53_63 V53 V63 14584.47112688824
L53_63 V53 V63 1.5766031709354506e-11
C53_63 V53 V63 -1.9111809732039624e-20

R53_64 V53 V64 10572.77592274378
L53_64 V53 V64 6.788436503392073e-12
C53_64 V53 V64 2.013646138900341e-20

R53_65 V53 V65 82496.35206677201
L53_65 V53 V65 2.5891614322983845e-11
C53_65 V53 V65 1.052955491164562e-20

R53_66 V53 V66 14396.763369643491
L53_66 V53 V66 4.26822018322414e-12
C53_66 V53 V66 1.5193344521115436e-19

R53_67 V53 V67 -59611.05312016734
L53_67 V53 V67 2.0000264947544102e-11
C53_67 V53 V67 7.004345873136807e-20

R53_68 V53 V68 288172.3130836479
L53_68 V53 V68 6.104510771064242e-12
C53_68 V53 V68 1.479787741789497e-19

R53_69 V53 V69 -2536.6553776891706
L53_69 V53 V69 -1.1552106618241487e-12
C53_69 V53 V69 -2.6261405186335265e-19

R53_70 V53 V70 -10056.649746149276
L53_70 V53 V70 -3.0047977614596425e-12
C53_70 V53 V70 -1.418758642727699e-19

R53_71 V53 V71 -20385.46566687992
L53_71 V53 V71 1.022008095405593e-11
C53_71 V53 V71 6.54272257959714e-20

R53_72 V53 V72 -7915.510591264986
L53_72 V53 V72 -4.4783059989301965e-11
C53_72 V53 V72 1.4350664020784714e-20

R53_73 V53 V73 -1669.8802131359591
L53_73 V53 V73 -4.0490115974098855e-12
C53_73 V53 V73 -1.0044114986815609e-19

R53_74 V53 V74 -8692.01333363438
L53_74 V53 V74 -3.394560318312766e-12
C53_74 V53 V74 -1.614840606703412e-19

R53_75 V53 V75 16555.417659527204
L53_75 V53 V75 -3.4616002619412575e-12
C53_75 V53 V75 -1.6567035524202263e-19

R53_76 V53 V76 13501.10992804234
L53_76 V53 V76 -2.015033143109987e-12
C53_76 V53 V76 -3.070443300257655e-19

R53_77 V53 V77 72766.02579883294
L53_77 V53 V77 1.0907077743037527e-12
C53_77 V53 V77 2.81210814565674e-19

R53_78 V53 V78 8553.856531290283
L53_78 V53 V78 1.0357266601120769e-11
C53_78 V53 V78 3.601494741172828e-21

R53_79 V53 V79 6919.2274413409605
L53_79 V53 V79 7.0102217024432174e-12
C53_79 V53 V79 6.860556190735547e-20

R53_80 V53 V80 4193.778230295306
L53_80 V53 V80 2.230698832062704e-12
C53_80 V53 V80 1.9005215219183946e-19

R53_81 V53 V81 -18201.15074638853
L53_81 V53 V81 -2.5190412240905598e-12
C53_81 V53 V81 -1.9251146520620368e-20

R53_82 V53 V82 20199.247396954244
L53_82 V53 V82 2.1757345025694587e-12
C53_82 V53 V82 2.9608441440132917e-19

R53_83 V53 V83 -66471.96493380834
L53_83 V53 V83 3.76622041667795e-12
C53_83 V53 V83 1.0498712547317253e-19

R53_84 V53 V84 9634.076363487598
L53_84 V53 V84 1.9078124265122977e-12
C53_84 V53 V84 2.143574517299296e-19

R53_85 V53 V85 5608.327940425837
L53_85 V53 V85 -8.993111977787402e-11
C53_85 V53 V85 3.2058020258290524e-20

R53_86 V53 V86 -18748.334189900623
L53_86 V53 V86 1.1785048352513983e-11
C53_86 V53 V86 4.8962437433243856e-20

R53_87 V53 V87 -6847.906896262718
L53_87 V53 V87 -2.7767765753992357e-12
C53_87 V53 V87 -1.8246502472625286e-19

R53_88 V53 V88 -4600.07199600399
L53_88 V53 V88 -1.6536948120012472e-12
C53_88 V53 V88 -2.5984173227300046e-19

R53_89 V53 V89 -1230.693730725869
L53_89 V53 V89 -1.6911479494146796e-12
C53_89 V53 V89 -2.1248559724677366e-19

R53_90 V53 V90 87637.53764891096
L53_90 V53 V90 -1.0586827906537696e-12
C53_90 V53 V90 -5.210642255924577e-19

R53_91 V53 V91 2733.952784406816
L53_91 V53 V91 3.489629027535099e-12
C53_91 V53 V91 1.836964123476517e-19

R53_92 V53 V92 2813.7732304021374
L53_92 V53 V92 3.318464108389365e-12
C53_92 V53 V92 9.418363459963261e-20

R53_93 V53 V93 11332.073458922368
L53_93 V53 V93 3.0327867848902385e-12
C53_93 V53 V93 1.222775549618906e-19

R53_94 V53 V94 -14747.005503758899
L53_94 V53 V94 4.3597541974187145e-12
C53_94 V53 V94 1.9410282310615872e-19

R53_95 V53 V95 8175.949213453275
L53_95 V53 V95 4.808579825719178e-12
C53_95 V53 V95 1.146796135753506e-19

R53_96 V53 V96 6702.86153742271
L53_96 V53 V96 4.471088857893618e-12
C53_96 V53 V96 1.5667322285003703e-19

R53_97 V53 V97 -2150.5351408580436
L53_97 V53 V97 1.6626900273803232e-12
C53_97 V53 V97 2.0816766709678612e-19

R53_98 V53 V98 5061.253143149383
L53_98 V53 V98 1.6551895164929798e-12
C53_98 V53 V98 2.9127204956796057e-19

R53_99 V53 V99 -2833.618467917742
L53_99 V53 V99 -1.844638877648556e-12
C53_99 V53 V99 -3.2362245966025654e-19

R53_100 V53 V100 -4648.383817840259
L53_100 V53 V100 -6.025786393503593e-12
C53_100 V53 V100 -1.9620225141194611e-19

R53_101 V53 V101 78277.42366937202
L53_101 V53 V101 -1.3873181710467695e-12
C53_101 V53 V101 -2.358493933690877e-19

R53_102 V53 V102 29160.47040122747
L53_102 V53 V102 -5.598610531662788e-12
C53_102 V53 V102 -1.9153389244765187e-19

R53_103 V53 V103 5407.349282669466
L53_103 V53 V103 4.0871576740055516e-12
C53_103 V53 V103 6.835824307373307e-20

R53_104 V53 V104 4004.6692584412954
L53_104 V53 V104 3.3314051979577136e-12
C53_104 V53 V104 6.424210344174837e-20

R53_105 V53 V105 -5254.096958709249
L53_105 V53 V105 -2.6134040411401574e-12
C53_105 V53 V105 -4.846220770119531e-20

R53_106 V53 V106 -5044.283601570923
L53_106 V53 V106 -1.4430218907100128e-12
C53_106 V53 V106 -2.3511488976903115e-19

R53_107 V53 V107 3337.8099964099883
L53_107 V53 V107 4.791124864048017e-12
C53_107 V53 V107 1.6264493613615307e-19

R53_108 V53 V108 7622.923303307139
L53_108 V53 V108 -2.7774364907537613e-12
C53_108 V53 V108 -3.8579623653870035e-20

R53_109 V53 V109 -3263.1336932722743
L53_109 V53 V109 6.5879534353935385e-12
C53_109 V53 V109 2.2970180518775562e-19

R53_110 V53 V110 4419.648647093691
L53_110 V53 V110 2.9572916025350104e-12
C53_110 V53 V110 1.7688416993766889e-19

R53_111 V53 V111 -2545.6015220283252
L53_111 V53 V111 -3.4465384046135028e-12
C53_111 V53 V111 -2.1584844316952702e-20

R53_112 V53 V112 -3148.5347826224947
L53_112 V53 V112 2.3120076073963912e-10
C53_112 V53 V112 7.224203973395652e-20

R53_113 V53 V113 -7580.886555145303
L53_113 V53 V113 1.5340786930551403e-12
C53_113 V53 V113 1.0751608636240685e-19

R53_114 V53 V114 6173.649206147812
L53_114 V53 V114 1.5890537612487414e-12
C53_114 V53 V114 2.1365194690284064e-19

R53_115 V53 V115 23399.822925114357
L53_115 V53 V115 -5.603056083802062e-12
C53_115 V53 V115 -1.29389614112063e-19

R53_116 V53 V116 82590.32614122209
L53_116 V53 V116 1.0615750402226394e-11
C53_116 V53 V116 -1.3466289925745429e-21

R53_117 V53 V117 -13690.647642100803
L53_117 V53 V117 -2.2048406530120333e-12
C53_117 V53 V117 -2.6023633214606755e-19

R53_118 V53 V118 -4124.310558726466
L53_118 V53 V118 -1.3799631684387207e-12
C53_118 V53 V118 -2.709421777171268e-19

R53_119 V53 V119 4730.539466095807
L53_119 V53 V119 -3.8156468311712826e-11
C53_119 V53 V119 -8.296002851948414e-20

R53_120 V53 V120 3513.9195725139007
L53_120 V53 V120 -4.776774467915919e-12
C53_120 V53 V120 -2.145966503332819e-19

R53_121 V53 V121 -5312.195972635586
L53_121 V53 V121 -3.6228843900983057e-12
C53_121 V53 V121 1.1665464421565852e-19

R53_122 V53 V122 88370.92516014658
L53_122 V53 V122 1.516626501959811e-11
C53_122 V53 V122 3.8217171927973605e-20

R53_123 V53 V123 -5183.815703369293
L53_123 V53 V123 3.0376997335235095e-12
C53_123 V53 V123 1.9334017989335955e-19

R53_124 V53 V124 -6493.791582339743
L53_124 V53 V124 2.4960956280899983e-12
C53_124 V53 V124 2.9400843790359466e-19

R53_125 V53 V125 -24190.815795950115
L53_125 V53 V125 8.301290387715589e-11
C53_125 V53 V125 -3.7334591637306374e-20

R53_126 V53 V126 3120.793731885037
L53_126 V53 V126 1.8884894889387105e-12
C53_126 V53 V126 1.3247868583370248e-19

R53_127 V53 V127 4926.068052927737
L53_127 V53 V127 1.779215491255203e-11
C53_127 V53 V127 1.4555314277586547e-20

R53_128 V53 V128 -75267.00420228219
L53_128 V53 V128 -6.366978096484716e-12
C53_128 V53 V128 1.548132754283273e-20

R53_129 V53 V129 -16594.40429192693
L53_129 V53 V129 -3.942631140448785e-11
C53_129 V53 V129 1.562553653185294e-19

R53_130 V53 V130 -9983.347164780896
L53_130 V53 V130 -2.506464712799426e-12
C53_130 V53 V130 -1.0995847436681707e-19

R53_131 V53 V131 -6558.58953841295
L53_131 V53 V131 -3.408574513075005e-12
C53_131 V53 V131 -1.0458036427642288e-19

R53_132 V53 V132 -19276.604985873473
L53_132 V53 V132 -3.0583513160669718e-12
C53_132 V53 V132 -2.1505146077838404e-19

R53_133 V53 V133 -4713.701261766345
L53_133 V53 V133 3.0412374794609796e-11
C53_133 V53 V133 -9.730984930842148e-20

R53_134 V53 V134 12803.541592475642
L53_134 V53 V134 3.0951581802801633e-12
C53_134 V53 V134 6.873777263621682e-20

R53_135 V53 V135 -8017.013612848655
L53_135 V53 V135 7.80012137582811e-12
C53_135 V53 V135 8.676833470474598e-20

R53_136 V53 V136 -6531.850042966772
L53_136 V53 V136 3.444520136560464e-12
C53_136 V53 V136 1.8228433408925077e-19

R53_137 V53 V137 4990.785274174328
L53_137 V53 V137 2.608948450631593e-12
C53_137 V53 V137 -1.2922941320410872e-19

R53_138 V53 V138 21944.46051589954
L53_138 V53 V138 5.437959505754345e-12
C53_138 V53 V138 1.16622808643021e-20

R53_139 V53 V139 4378.185401145118
L53_139 V53 V139 -4.868653229455931e-12
C53_139 V53 V139 -2.001004564527016e-19

R53_140 V53 V140 3525.879829344557
L53_140 V53 V140 1.9998175080763568e-11
C53_140 V53 V140 -2.193289004460656e-19

R53_141 V53 V141 -51858.309220067844
L53_141 V53 V141 -1.017720420666279e-11
C53_141 V53 V141 2.069327735156455e-19

R53_142 V53 V142 -8210.524570217654
L53_142 V53 V142 -1.9351431982518883e-12
C53_142 V53 V142 -4.176502111644107e-20

R53_143 V53 V143 -20927.76849587871
L53_143 V53 V143 4.274065548963905e-12
C53_143 V53 V143 1.4933579747731068e-19

R53_144 V53 V144 10736.43671253083
L53_144 V53 V144 -3.794410751369159e-12
C53_144 V53 V144 8.9199998202384e-20

R53_145 V53 V145 -2081.659705639274
L53_145 V53 V145 -1.7396873600895546e-12
C53_145 V53 V145 1.9799875808607256e-19

R53_146 V53 V146 -11113.64573529134
L53_146 V53 V146 -5.067725846610005e-12
C53_146 V53 V146 3.3432220918398788e-21

R53_147 V53 V147 5691.260903976618
L53_147 V53 V147 1.727758935341184e-10
C53_147 V53 V147 2.035586765389336e-19

R53_148 V53 V148 -3913.54671408806
L53_148 V53 V148 4.135995395520457e-12
C53_148 V53 V148 1.4379496878080352e-19

R53_149 V53 V149 7030.130003215133
L53_149 V53 V149 -1.936040568328303e-12
C53_149 V53 V149 -5.238653853986268e-19

R53_150 V53 V150 4053.6773716872876
L53_150 V53 V150 1.669129024504895e-12
C53_150 V53 V150 2.4506504404770176e-19

R53_151 V53 V151 -1639.2654707713104
L53_151 V53 V151 -4.138170550146258e-12
C53_151 V53 V151 -1.7517652308435022e-19

R53_152 V53 V152 -20655.613305168936
L53_152 V53 V152 2.59717884650353e-10
C53_152 V53 V152 -3.456751444637938e-20

R53_153 V53 V153 3747.976628215959
L53_153 V53 V153 1.7642744740873347e-12
C53_153 V53 V153 -6.322695029401875e-20

R53_154 V53 V154 -42772.66838804209
L53_154 V53 V154 3.805909060659338e-12
C53_154 V53 V154 -2.010725724691461e-19

R53_155 V53 V155 1150.1528937652238
L53_155 V53 V155 -2.7745063604795677e-12
C53_155 V53 V155 -1.4500408661093917e-19

R53_156 V53 V156 -204446.96140295657
L53_156 V53 V156 6.098137813202779e-12
C53_156 V53 V156 -1.8804605474664172e-19

R53_157 V53 V157 -1684.5513358462285
L53_157 V53 V157 9.74311154893384e-13
C53_157 V53 V157 5.132802918839061e-19

R53_158 V53 V158 -6899.799688491259
L53_158 V53 V158 -1.5638495876388617e-12
C53_158 V53 V158 -5.779997001300064e-20

R53_159 V53 V159 -9007.53508827256
L53_159 V53 V159 3.1022357543525924e-12
C53_159 V53 V159 3.790673010585707e-20

R53_160 V53 V160 2763.7066579344582
L53_160 V53 V160 -6.457841170637877e-12
C53_160 V53 V160 3.2734536891646564e-20

R53_161 V53 V161 2469.7436815291176
L53_161 V53 V161 -2.880961279251197e-12
C53_161 V53 V161 2.5706795383701458e-20

R53_162 V53 V162 -11515.964980863893
L53_162 V53 V162 -2.570696363710568e-12
C53_162 V53 V162 -3.287996980533793e-20

R53_163 V53 V163 67902.1686756516
L53_163 V53 V163 2.4178728946983653e-12
C53_163 V53 V163 9.4933819733356e-20

R53_164 V53 V164 -3477.3790786148656
L53_164 V53 V164 6.540587539445072e-12
C53_164 V53 V164 -3.6494010210332165e-21

R53_165 V53 V165 -858.533231084012
L53_165 V53 V165 -6.779424950066608e-13
C53_165 V53 V165 -3.897350684022107e-19

R53_166 V53 V166 -30963.160533092087
L53_166 V53 V166 2.052814582697035e-12
C53_166 V53 V166 1.1260342513886433e-19

R53_167 V53 V167 -6597.632090526196
L53_167 V53 V167 -3.161266555348879e-12
C53_167 V53 V167 -2.8422808232543124e-20

R53_168 V53 V168 2404.740184146325
L53_168 V53 V168 -4.14536852683748e-12
C53_168 V53 V168 6.513263502181319e-20

R53_169 V53 V169 6802.71631701299
L53_169 V53 V169 1.914138297086039e-12
C53_169 V53 V169 1.719319315299312e-19

R53_170 V53 V170 -5450.185106181988
L53_170 V53 V170 -2.8746257713616467e-12
C53_170 V53 V170 -1.620668902701167e-19

R53_171 V53 V171 -12236.219516296884
L53_171 V53 V171 -1.4628228136531443e-12
C53_171 V53 V171 -1.2988223399063606e-19

R53_172 V53 V172 -3569.284657277886
L53_172 V53 V172 -1.3196486129547224e-11
C53_172 V53 V172 -8.004950455604547e-20

R53_173 V53 V173 2058.0214805749183
L53_173 V53 V173 1.5269026043999996e-12
C53_173 V53 V173 5.684855677842576e-20

R53_174 V53 V174 2835.7114268997548
L53_174 V53 V174 2.0115255079382363e-11
C53_174 V53 V174 7.74788114210799e-20

R53_175 V53 V175 12195.719207840675
L53_175 V53 V175 3.497927317401116e-12
C53_175 V53 V175 -9.497513495120811e-20

R53_176 V53 V176 8608.697955181273
L53_176 V53 V176 3.974474798827803e-12
C53_176 V53 V176 -1.1898797972076218e-19

R53_177 V53 V177 -1444.247699321235
L53_177 V53 V177 -4.154405948694891e-11
C53_177 V53 V177 2.034506422668766e-20

R53_178 V53 V178 8941.45165230833
L53_178 V53 V178 2.20062824826065e-12
C53_178 V53 V178 1.291213207632133e-19

R53_179 V53 V179 2747.5798718999845
L53_179 V53 V179 1.6771567112199342e-12
C53_179 V53 V179 2.7071931943633765e-19

R53_180 V53 V180 3434.349899064358
L53_180 V53 V180 2.8640258236979865e-12
C53_180 V53 V180 2.496449155647961e-19

R53_181 V53 V181 1313.1651801807568
L53_181 V53 V181 -6.341656459594061e-12
C53_181 V53 V181 -5.944523688208072e-20

R53_182 V53 V182 -3402.949877933066
L53_182 V53 V182 -1.7084677973038489e-12
C53_182 V53 V182 -1.610033000044081e-19

R53_183 V53 V183 -2931.2761833009513
L53_183 V53 V183 3.4253020032577825e-12
C53_183 V53 V183 1.662202995256802e-20

R53_184 V53 V184 -2188.0387740409637
L53_184 V53 V184 1.9093983676217586e-11
C53_184 V53 V184 -2.4282851353845367e-20

R53_185 V53 V185 -4650.6229417048335
L53_185 V53 V185 -1.9755219399264882e-12
C53_185 V53 V185 -3.799248427205651e-20

R53_186 V53 V186 -2299.138033165159
L53_186 V53 V186 -2.282023628733889e-12
C53_186 V53 V186 3.3243187558827253e-21

R53_187 V53 V187 -3220.385288598612
L53_187 V53 V187 -1.2035659630995012e-12
C53_187 V53 V187 -2.1129522533090836e-19

R53_188 V53 V188 -8454.326982590188
L53_188 V53 V188 -9.580552689847934e-13
C53_188 V53 V188 -1.8309125813586244e-19

R53_189 V53 V189 -19596.30908082576
L53_189 V53 V189 5.373855559808509e-12
C53_189 V53 V189 2.4309022593542188e-21

R53_190 V53 V190 2687.417609347059
L53_190 V53 V190 2.7874596965214694e-12
C53_190 V53 V190 1.322341333235454e-19

R53_191 V53 V191 2806.822746205154
L53_191 V53 V191 -1.9133364141537234e-12
C53_191 V53 V191 -6.000012517949978e-21

R53_192 V53 V192 2545.731340072239
L53_192 V53 V192 3.5229543039005222e-12
C53_192 V53 V192 9.248391098964075e-20

R53_193 V53 V193 -4150.30009101871
L53_193 V53 V193 1.4542434363496905e-12
C53_193 V53 V193 9.063645546561275e-20

R53_194 V53 V194 1451.9048059601607
L53_194 V53 V194 2.231993069343326e-12
C53_194 V53 V194 6.612313182129085e-20

R53_195 V53 V195 13918.04441616556
L53_195 V53 V195 1.2339582308529643e-12
C53_195 V53 V195 1.2784153655928308e-19

R53_196 V53 V196 14815.82340356505
L53_196 V53 V196 1.6725181884665617e-12
C53_196 V53 V196 -2.6185161501792152e-21

R53_197 V53 V197 2680.334829631128
L53_197 V53 V197 6.509947887949078e-12
C53_197 V53 V197 7.054000389612392e-20

R53_198 V53 V198 -1472.9852736460812
L53_198 V53 V198 -6.5559969021331015e-12
C53_198 V53 V198 -1.0800518489063827e-20

R53_199 V53 V199 -1327.6229563871495
L53_199 V53 V199 2.5646727569072204e-12
C53_199 V53 V199 4.193692857784603e-20

R53_200 V53 V200 -1966.9634889781385
L53_200 V53 V200 3.392914245682384e-11
C53_200 V53 V200 2.8343113173490025e-20

R54_54 V54 0 -1353.8312175105182
L54_54 V54 0 -3.477352294902722e-13
C54_54 V54 0 -2.4843253414856848e-18

R54_55 V54 V55 -6663.033153874002
L54_55 V54 V55 -3.4795269923439177e-12
C54_55 V54 V55 -1.8108852056428998e-19

R54_56 V54 V56 -3147.48064060447
L54_56 V54 V56 -1.7606282054258568e-12
C54_56 V54 V56 -3.487599915541197e-19

R54_57 V54 V57 122187.61378461898
L54_57 V54 V57 5.6740106429072096e-11
C54_57 V54 V57 -3.93110881166964e-20

R54_58 V54 V58 2832.8722949161406
L54_58 V54 V58 6.385817175710831e-13
C54_58 V54 V58 7.6978155743069815e-19

R54_59 V54 V59 5878.4823855472005
L54_59 V54 V59 3.8842732435591125e-11
C54_59 V54 V59 3.8533213890132277e-20

R54_60 V54 V60 6048.617664657577
L54_60 V54 V60 1.5002186578921643e-11
C54_60 V54 V60 3.7413108736762916e-20

R54_61 V54 V61 5298.894217283183
L54_61 V54 V61 3.3718726053679407e-12
C54_61 V54 V61 2.0577683752498907e-19

R54_62 V54 V62 -5057.002560206478
L54_62 V54 V62 5.621326526669749e-13
C54_62 V54 V62 1.1921338057512934e-18

R54_63 V54 V63 22480.59769366133
L54_63 V54 V63 1.281613981944674e-10
C54_63 V54 V63 -3.0295774500375164e-21

R54_64 V54 V64 6338.172429992964
L54_64 V54 V64 3.715906089013921e-12
C54_64 V54 V64 1.1461837975308584e-19

R54_65 V54 V65 42263.427433437035
L54_65 V54 V65 8.40511939982293e-12
C54_65 V54 V65 1.155606531244672e-19

R54_66 V54 V66 2684.3979182129196
L54_66 V54 V66 -1.1311247542380797e-12
C54_66 V54 V66 -5.974791837407368e-19

R54_67 V54 V67 -8972.553235341975
L54_67 V54 V67 -5.2021967134768065e-12
C54_67 V54 V67 -1.3384900645517035e-19

R54_68 V54 V68 -34961.09496293537
L54_68 V54 V68 3.183548198806971e-11
C54_68 V54 V68 -3.4540452480107684e-20

R54_69 V54 V69 -3053.5161914799633
L54_69 V54 V69 -1.7495358748310765e-12
C54_69 V54 V69 -2.9717627649363744e-19

R54_70 V54 V70 3226.7853170924577
L54_70 V54 V70 -1.2115576723289714e-12
C54_70 V54 V70 -4.267474121329662e-19

R54_71 V54 V71 15767.93189604918
L54_71 V54 V71 3.2109784314585753e-12
C54_71 V54 V71 1.6691592284732312e-19

R54_72 V54 V72 30729.0494131899
L54_72 V54 V72 2.706677404851472e-11
C54_72 V54 V72 4.5559882786508634e-21

R54_73 V54 V73 20514.213515123727
L54_73 V54 V73 5.301775280457511e-12
C54_73 V54 V73 1.2290620328521197e-19

R54_74 V54 V74 -1619.560163964763
L54_74 V54 V74 3.280788154246493e-12
C54_74 V54 V74 3.1460124257108684e-19

R54_75 V54 V75 6242.541400967828
L54_75 V54 V75 -1.8230302694432814e-11
C54_75 V54 V75 1.0821656002081688e-20

R54_76 V54 V76 -12741.959011721743
L54_76 V54 V76 -2.041083394966559e-12
C54_76 V54 V76 -2.0239986754505172e-19

R54_77 V54 V77 38754.15088976683
L54_77 V54 V77 9.361682694893325e-12
C54_77 V54 V77 4.5573845078893294e-20

R54_78 V54 V78 -348453.8513815195
L54_78 V54 V78 1.7055462744100025e-12
C54_78 V54 V78 1.0281847550208062e-19

R54_79 V54 V79 -6936.084429112274
L54_79 V54 V79 -9.000940578196327e-12
C54_79 V54 V79 -8.754810421276215e-20

R54_80 V54 V80 -315577.5137670457
L54_80 V54 V80 2.484443615823932e-12
C54_80 V54 V80 1.228967122247083e-19

R54_81 V54 V81 174563.6806351766
L54_81 V54 V81 1.7102560940804903e-11
C54_81 V54 V81 9.069158742952951e-20

R54_82 V54 V82 3760.151886345975
L54_82 V54 V82 2.810139787802023e-11
C54_82 V54 V82 1.1235276685473867e-19

R54_83 V54 V83 82028.48076113482
L54_83 V54 V83 2.3485098664721802e-11
C54_83 V54 V83 1.0209917783471849e-20

R54_84 V54 V84 6136.594496021944
L54_84 V54 V84 2.420116782107466e-12
C54_84 V54 V84 1.758520404379517e-19

R54_85 V54 V85 -28838.07490248764
L54_85 V54 V85 3.445383982444634e-12
C54_85 V54 V85 1.9374726411816377e-19

R54_86 V54 V86 1152.0710356126156
L54_86 V54 V86 -4.5389413359435995e-12
C54_86 V54 V86 -5.509482557351226e-20

R54_87 V54 V87 -15612.324817718221
L54_87 V54 V87 -3.4584568819068975e-12
C54_87 V54 V87 -1.355315317957255e-19

R54_88 V54 V88 -10251.681922000309
L54_88 V54 V88 -1.6766728190894883e-12
C54_88 V54 V88 -2.6477685102429645e-19

R54_89 V54 V89 -3413.7978262976744
L54_89 V54 V89 -1.2701281048028712e-12
C54_89 V54 V89 -3.7946656902960464e-19

R54_90 V54 V90 -1006.7391143148333
L54_90 V54 V90 -1.5340655361983384e-12
C54_90 V54 V90 -4.877215686411843e-19

R54_91 V54 V91 5330.5220441296515
L54_91 V54 V91 1.3837219979348566e-12
C54_91 V54 V91 3.1614595272089697e-19

R54_92 V54 V92 7285.560883799427
L54_92 V54 V92 1.9746706834321827e-12
C54_92 V54 V92 1.2275733414921747e-19

R54_93 V54 V93 11641.283551338773
L54_93 V54 V93 1.3296783874552942e-11
C54_93 V54 V93 2.0392791306849813e-20

R54_94 V54 V94 -3174.7967631783135
L54_94 V54 V94 2.2233505285939436e-12
C54_94 V54 V94 3.371157345303879e-19

R54_95 V54 V95 7576.57508962583
L54_95 V54 V95 1.3335430690878046e-11
C54_95 V54 V95 1.196108650166689e-19

R54_96 V54 V96 -51155.64263243368
L54_96 V54 V96 1.2658549124480091e-11
C54_96 V54 V96 1.9019496090617003e-19

R54_97 V54 V97 -4660.465497042347
L54_97 V54 V97 1.19152416839936e-12
C54_97 V54 V97 4.861523643424208e-19

R54_98 V54 V98 1311.9433914122583
L54_98 V54 V98 2.5778506240588695e-12
C54_98 V54 V98 2.629489160227643e-19

R54_99 V54 V99 -1647.0516537983617
L54_99 V54 V99 -9.930966072859994e-13
C54_99 V54 V99 -5.281481645080692e-19

R54_100 V54 V100 -3140.3829381712126
L54_100 V54 V100 -3.093632529573986e-12
C54_100 V54 V100 -2.70898983104042e-19

R54_101 V54 V101 -47138.91237105376
L54_101 V54 V101 -1.987146332311519e-12
C54_101 V54 V101 -2.574212246427221e-19

R54_102 V54 V102 -3046.8002751360395
L54_102 V54 V102 -2.1551118946974883e-12
C54_102 V54 V102 -3.0691331535022613e-19

R54_103 V54 V103 2250.3304800302567
L54_103 V54 V103 5.584504567985501e-12
C54_103 V54 V103 -1.1430195880773698e-20

R54_104 V54 V104 1844.4841503848736
L54_104 V54 V104 5.662861109691344e-12
C54_104 V54 V104 -2.351466253142449e-20

R54_105 V54 V105 119121.06509916116
L54_105 V54 V105 -1.3962582358026166e-12
C54_105 V54 V105 -2.33996375534025e-19

R54_106 V54 V106 1230.2420608703594
L54_106 V54 V106 -2.9663845994372683e-12
C54_106 V54 V106 -1.6475918101087786e-19

R54_107 V54 V107 4712.392239285561
L54_107 V54 V107 1.4308590316158524e-12
C54_107 V54 V107 4.487129685341839e-19

R54_108 V54 V108 -17006.31123103466
L54_108 V54 V108 -6.928927597865425e-12
C54_108 V54 V108 7.325216760299582e-20

R54_109 V54 V109 -6944.032413954209
L54_109 V54 V109 1.977319149082962e-12
C54_109 V54 V109 3.7201284895267394e-19

R54_110 V54 V110 -1203.0814988689876
L54_110 V54 V110 2.1493867456663266e-12
C54_110 V54 V110 1.8327762797102156e-19

R54_111 V54 V111 -2640.4332126804243
L54_111 V54 V111 8.392141741336331e-11
C54_111 V54 V111 2.885357115635321e-20

R54_112 V54 V112 -3080.0483438590827
L54_112 V54 V112 3.495502524339076e-12
C54_112 V54 V112 1.4138529974859943e-19

R54_113 V54 V113 -8483.561017716731
L54_113 V54 V113 1.2971116139187489e-12
C54_113 V54 V113 1.979669438282963e-19

R54_114 V54 V114 -2344.419715142529
L54_114 V54 V114 1.8184317697417465e-12
C54_114 V54 V114 2.7164497896590594e-19

R54_115 V54 V115 -11642.866195339195
L54_115 V54 V115 -1.1977947902754372e-12
C54_115 V54 V115 -3.9432808378133576e-19

R54_116 V54 V116 -76896.41060431358
L54_116 V54 V116 -2.979893982359686e-12
C54_116 V54 V116 -1.2798821127900284e-19

R54_117 V54 V117 -3709.8824309295273
L54_117 V54 V117 -1.4501604074218483e-12
C54_117 V54 V117 -2.981396926909997e-19

R54_118 V54 V118 709.6651077450601
L54_118 V54 V118 -8.018068198093775e-13
C54_118 V54 V118 -3.992448035419449e-19

R54_119 V54 V119 2492.5894803048536
L54_119 V54 V119 -4.038107430152174e-11
C54_119 V54 V119 -5.2909116090216775e-20

R54_120 V54 V120 2424.1511137731795
L54_120 V54 V120 -3.244439134138683e-12
C54_120 V54 V120 -2.545895433662616e-19

R54_121 V54 V121 3141.5362093761755
L54_121 V54 V121 -2.0598926810213934e-12
C54_121 V54 V121 -6.68767786484795e-20

R54_122 V54 V122 -4444.923270848213
L54_122 V54 V122 1.7763195850661844e-12
C54_122 V54 V122 1.8999961504018357e-19

R54_123 V54 V123 -38361.504476932074
L54_123 V54 V123 1.5130618290174436e-12
C54_123 V54 V123 2.987943623177808e-19

R54_124 V54 V124 -41113.92814496876
L54_124 V54 V124 1.1940487305330517e-12
C54_124 V54 V124 4.283612013883737e-19

R54_125 V54 V125 2502.2589621264724
L54_125 V54 V125 3.4233378300554583e-12
C54_125 V54 V125 7.237887703702895e-20

R54_126 V54 V126 -1056.5426036760186
L54_126 V54 V126 9.836366951750286e-13
C54_126 V54 V126 1.793626717180195e-19

R54_127 V54 V127 -1986.6286466289512
L54_127 V54 V127 6.089421739317196e-12
C54_127 V54 V127 7.790057069588074e-20

R54_128 V54 V128 -1570.3177080166236
L54_128 V54 V128 2.6844537369741725e-10
C54_128 V54 V128 8.122798188505812e-20

R54_129 V54 V129 -1216.336970404136
L54_129 V54 V129 1.260176710748367e-12
C54_129 V54 V129 5.058188352990831e-19

R54_130 V54 V130 3245.7769309955647
L54_130 V54 V130 -8.95606480165224e-13
C54_130 V54 V130 -3.6639577640751673e-19

R54_131 V54 V131 1731.3014376633564
L54_131 V54 V131 -1.7489262868067731e-12
C54_131 V54 V131 -2.2986288188101426e-19

R54_132 V54 V132 1258.0416627732775
L54_132 V54 V132 -1.0869473277837538e-12
C54_132 V54 V132 -4.609332723634267e-19

R54_133 V54 V133 -4532.660687801007
L54_133 V54 V133 -1.1746367794720582e-12
C54_133 V54 V133 -5.07521218738486e-19

R54_134 V54 V134 864.7507134060603
L54_134 V54 V134 1.9702523983500212e-12
C54_134 V54 V134 4.337769864456116e-19

R54_135 V54 V135 3557.3259841326844
L54_135 V54 V135 2.9032162984454705e-11
C54_135 V54 V135 4.667661837343925e-20

R54_136 V54 V136 1717.9317641753635
L54_136 V54 V136 3.83440276295416e-12
C54_136 V54 V136 2.571920180163581e-19

R54_137 V54 V137 927.8957126978906
L54_137 V54 V137 -2.780776214432593e-12
C54_137 V54 V137 -3.338226206110317e-19

R54_138 V54 V138 -1200.1871511283707
L54_138 V54 V138 4.654496251865558e-12
C54_138 V54 V138 -1.483047293875599e-19

R54_139 V54 V139 -1319.221954341383
L54_139 V54 V139 -8.475365587873178e-11
C54_139 V54 V139 -1.607529279122682e-19

R54_140 V54 V140 -1048.6495971912295
L54_140 V54 V140 2.548168865022572e-12
C54_140 V54 V140 -1.9208706875172747e-19

R54_141 V54 V141 3845.896605296861
L54_141 V54 V141 9.602341073128293e-13
C54_141 V54 V141 8.171333915623956e-19

R54_142 V54 V142 -625.2182164922045
L54_142 V54 V142 -3.3176106138411635e-12
C54_142 V54 V142 -1.7566096709773834e-19

R54_143 V54 V143 4126.620267550707
L54_143 V54 V143 4.45943571732499e-12
C54_143 V54 V143 2.5553044719419585e-19

R54_144 V54 V144 -4130.033736697399
L54_144 V54 V144 -2.5063073067645963e-12
C54_144 V54 V144 1.2092851299441778e-19

R54_145 V54 V145 -748.5650361730686
L54_145 V54 V145 3.827875225824538e-12
C54_145 V54 V145 2.8187978805144805e-19

R54_146 V54 V146 542.3208560748214
L54_146 V54 V146 3.3623729856115277e-12
C54_146 V54 V146 6.080996316795518e-20

R54_147 V54 V147 9164.49588663268
L54_147 V54 V147 4.6672376208750515e-12
C54_147 V54 V147 1.8014878628128581e-19

R54_148 V54 V148 1002.7200162436783
L54_148 V54 V148 1.3250344978300753e-12
C54_148 V54 V148 1.826276922838263e-19

R54_149 V54 V149 -9389.153778559394
L54_149 V54 V149 -5.17194305215014e-13
C54_149 V54 V149 -1.190458827468806e-18

R54_150 V54 V150 711.3881153707246
L54_150 V54 V150 -1.6538364739639174e-12
C54_150 V54 V150 6.652695470718694e-19

R54_151 V54 V151 -2294.1608943091005
L54_151 V54 V151 6.7505098475204215e-12
C54_151 V54 V151 -2.4504872865567294e-19

R54_152 V54 V152 -820.3983637028734
L54_152 V54 V152 4.837153207455977e-12
C54_152 V54 V152 -3.716464166676559e-20

R54_153 V54 V153 890.201037885445
L54_153 V54 V153 -1.0797701387252942e-10
C54_153 V54 V153 -1.145499761539309e-19

R54_154 V54 V154 -1180.3009575339988
L54_154 V54 V154 -1.185533186933229e-11
C54_154 V54 V154 -5.166636145320977e-19

R54_155 V54 V155 -69216.78365655841
L54_155 V54 V155 -1.3143403240725827e-12
C54_155 V54 V155 -2.222558809006325e-19

R54_156 V54 V156 709.792518393644
L54_156 V54 V156 -7.340223577754062e-12
C54_156 V54 V156 -2.5129805045723276e-19

R54_157 V54 V157 3471.339884635115
L54_157 V54 V157 5.55053020418395e-13
C54_157 V54 V157 1.0955295334113361e-18

R54_158 V54 V158 -1411.5713403683671
L54_158 V54 V158 1.1920287874496987e-12
C54_158 V54 V158 -3.108203225474903e-20

R54_159 V54 V159 844.8611157910849
L54_159 V54 V159 -3.530222767590756e-12
C54_159 V54 V159 1.0373657202654712e-21

R54_160 V54 V160 3052.5541854939543
L54_160 V54 V160 -9.969215120107261e-13
C54_160 V54 V160 -3.132446179193845e-20

R54_161 V54 V161 -955.7897142673968
L54_161 V54 V161 4.696203524051679e-12
C54_161 V54 V161 7.602453938810534e-20

R54_162 V54 V162 -9758.270404986331
L54_162 V54 V162 2.3489095334862886e-11
C54_162 V54 V162 -1.0620725600306576e-19

R54_163 V54 V163 -1194.9592324346822
L54_163 V54 V163 1.2194856032061383e-12
C54_163 V54 V163 1.8932034034188897e-19

R54_164 V54 V164 -1168.1163544546002
L54_164 V54 V164 1.1576062459491176e-12
C54_164 V54 V164 -1.554242498716923e-20

R54_165 V54 V165 -30322.229322097155
L54_165 V54 V165 -8.731047716563632e-13
C54_165 V54 V165 -5.92474858630915e-19

R54_166 V54 V166 628.147900271081
L54_166 V54 V166 -7.448864456077742e-13
C54_166 V54 V166 1.8448618833614803e-19

R54_167 V54 V167 -10020.852048638151
L54_167 V54 V167 1.3222997588572638e-12
C54_167 V54 V167 3.565721110455073e-20

R54_168 V54 V168 -2304.721470740715
L54_168 V54 V168 1.191404671691375e-12
C54_168 V54 V168 2.2877633948530704e-19

R54_169 V54 V169 840.1892068385961
L54_169 V54 V169 -2.3840620390901863e-12
C54_169 V54 V169 9.553726233954738e-20

R54_170 V54 V170 -1519.5072534378478
L54_170 V54 V170 -3.4272677121992945e-12
C54_170 V54 V170 -3.0694802459012696e-19

R54_171 V54 V171 2809.991760972001
L54_171 V54 V171 -6.119943312775561e-13
C54_171 V54 V171 -3.805979126575435e-19

R54_172 V54 V172 1834.0765788655635
L54_172 V54 V172 -1.0227959758653637e-12
C54_172 V54 V172 -2.584361127948493e-19

R54_173 V54 V173 -1902.884426673246
L54_173 V54 V173 9.82746170210307e-13
C54_173 V54 V173 1.4987899917829557e-19

R54_174 V54 V174 -711.0593005977437
L54_174 V54 V174 6.025327269835388e-13
C54_174 V54 V174 2.5386712081305653e-19

R54_175 V54 V175 71149.34164788807
L54_175 V54 V175 -2.7573884269477197e-12
C54_175 V54 V175 -1.7494945488343488e-19

R54_176 V54 V176 12058.573007097906
L54_176 V54 V176 -1.6991308918376208e-12
C54_176 V54 V176 -2.2488373683375495e-19

R54_177 V54 V177 -5328.277300357014
L54_177 V54 V177 2.9792180697858133e-12
C54_177 V54 V177 -3.982118282505298e-20

R54_178 V54 V178 963.36053936529
L54_178 V54 V178 4.914366581816611e-12
C54_178 V54 V178 1.613608550657514e-19

R54_179 V54 V179 9020.738508442877
L54_179 V54 V179 6.968107691668532e-13
C54_179 V54 V179 5.611363156256379e-19

R54_180 V54 V180 4333.354728314198
L54_180 V54 V180 6.716623078091135e-13
C54_180 V54 V180 4.850482809639733e-19

R54_181 V54 V181 2278.007109014691
L54_181 V54 V181 -1.4811194985734192e-12
C54_181 V54 V181 1.1215978272146935e-19

R54_182 V54 V182 2357.5153085531347
L54_182 V54 V182 -4.915309834479429e-13
C54_182 V54 V182 -3.1326998599146285e-19

R54_183 V54 V183 6786.370000491528
L54_183 V54 V183 2.2832368941452105e-12
C54_183 V54 V183 7.247321100256946e-20

R54_184 V54 V184 -9708.27098838111
L54_184 V54 V184 5.41762874111866e-12
C54_184 V54 V184 -2.796692406951915e-20

R54_185 V54 V185 -15471.830641105844
L54_185 V54 V185 -2.2529010081142653e-11
C54_185 V54 V185 -8.088173156133198e-20

R54_186 V54 V186 -1168.7555766892353
L54_186 V54 V186 -2.8948540432967876e-11
C54_186 V54 V186 1.2011113316964648e-19

R54_187 V54 V187 -1761.3179927742801
L54_187 V54 V187 -9.737078991442107e-13
C54_187 V54 V187 -4.1985872800749256e-19

R54_188 V54 V188 -1100.133575783023
L54_188 V54 V188 -6.855255944900496e-13
C54_188 V54 V188 -3.305073164523913e-19

R54_189 V54 V189 3196.155791318131
L54_189 V54 V189 4.592169306910299e-12
C54_189 V54 V189 -2.336148900412798e-19

R54_190 V54 V190 2301.865597616165
L54_190 V54 V190 7.904779205064973e-13
C54_190 V54 V190 2.824193840008707e-19

R54_191 V54 V191 9875.454820089524
L54_191 V54 V191 -1.5345734524368187e-12
C54_191 V54 V191 -2.0739025015847196e-19

R54_192 V54 V192 2020.3999937730596
L54_192 V54 V192 6.149733080774427e-12
C54_192 V54 V192 -9.429250478700281e-20

R54_193 V54 V193 -1893.6856309267014
L54_193 V54 V193 8.984171345287895e-12
C54_193 V54 V193 1.710972036669106e-19

R54_194 V54 V194 2457.242180699061
L54_194 V54 V194 -6.179441403686999e-11
C54_194 V54 V194 5.720207250702506e-20

R54_195 V54 V195 2022.0483540298137
L54_195 V54 V195 8.025903941267649e-13
C54_195 V54 V195 4.931110762597426e-19

R54_196 V54 V196 1982.5097747260868
L54_196 V54 V196 9.962093427012542e-13
C54_196 V54 V196 3.115577860433598e-19

R54_197 V54 V197 -45038.39802951536
L54_197 V54 V197 6.401652262509239e-12
C54_197 V54 V197 2.3868250653459104e-19

R54_198 V54 V198 -2412.3515751654486
L54_198 V54 V198 -8.785781637602503e-13
C54_198 V54 V198 -5.006990670810013e-20

R54_199 V54 V199 -4566.143778581429
L54_199 V54 V199 5.426112322570051e-12
C54_199 V54 V199 1.59638841798334e-19

R54_200 V54 V200 -1177.0318031322015
L54_200 V54 V200 2.090294381457398e-11
C54_200 V54 V200 8.635166676668852e-20

R55_55 V55 0 761.7683448076725
L55_55 V55 0 -2.012023828720865e-12
C55_55 V55 0 -1.166372386500966e-18

R55_56 V55 V56 -4327.113563280169
L55_56 V55 V56 -3.7596769718444815e-12
C55_56 V55 V56 -1.4045291155569399e-19

R55_57 V55 V57 -110246.50396451127
L55_57 V55 V57 1.2829321581828392e-11
C55_57 V55 V57 -2.3152361189241736e-20

R55_58 V55 V58 5962.139588823207
L55_58 V55 V58 -6.12737434882893e-12
C55_58 V55 V58 -1.1559004765220701e-19

R55_59 V55 V59 -29466.40191200487
L55_59 V55 V59 8.656277981580593e-13
C55_59 V55 V59 5.875863084815007e-19

R55_60 V55 V60 11519.101055045521
L55_60 V55 V60 -1.110536965600316e-11
C55_60 V55 V60 -6.986683681506814e-20

R55_61 V55 V61 6894.05168768809
L55_61 V55 V61 4.947738726118777e-12
C55_61 V55 V61 1.3466301693041423e-19

R55_62 V55 V62 -30176.029475839103
L55_62 V55 V62 3.855014622667484e-12
C55_62 V55 V62 1.5774821132971942e-19

R55_63 V55 V63 200810.28331935065
L55_63 V55 V63 9.020105383405044e-13
C55_63 V55 V63 7.250392713920972e-19

R55_64 V55 V64 6916.487020815847
L55_64 V55 V64 1.0119495752083798e-11
C55_64 V55 V64 2.2291842804458438e-20

R55_65 V55 V65 -12950.360545342228
L55_65 V55 V65 -1.8080427053246745e-11
C55_65 V55 V65 1.5735073827918945e-20

R55_66 V55 V66 25709.11992600198
L55_66 V55 V66 9.3711962750473e-12
C55_66 V55 V66 9.312641290849505e-20

R55_67 V55 V67 2912.7295226238584
L55_67 V55 V67 -1.089731251908012e-12
C55_67 V55 V67 -6.369000723142844e-19

R55_68 V55 V68 17766.73508873277
L55_68 V55 V68 1.546477620964058e-11
C55_68 V55 V68 7.200281692688292e-22

R55_69 V55 V69 -5674.868652285264
L55_69 V55 V69 -2.8774823256337687e-12
C55_69 V55 V69 -1.6063723082649912e-19

R55_70 V55 V70 61491.337135124704
L55_70 V55 V70 -5.701142010256825e-12
C55_70 V55 V70 -8.54560362073131e-20

R55_71 V55 V71 4491.94667872794
L55_71 V55 V71 -7.334927107665499e-12
C55_71 V55 V71 -7.131409590016303e-20

R55_72 V55 V72 -46567.48839802815
L55_72 V55 V72 7.758153124301235e-12
C55_72 V55 V72 8.537792269643559e-20

R55_73 V55 V73 -76440.14951262774
L55_73 V55 V73 5.050151189983575e-12
C55_73 V55 V73 1.4707577321247352e-19

R55_74 V55 V74 -13649.643146663644
L55_74 V55 V74 -3.916650042818075e-11
C55_74 V55 V74 -4.027775887696827e-21

R55_75 V55 V75 -2007.5625884002063
L55_75 V55 V75 2.7634059644091594e-12
C55_75 V55 V75 3.791078567318644e-19

R55_76 V55 V76 -11837.146536369859
L55_76 V55 V76 -2.3532874799543467e-12
C55_76 V55 V76 -1.6688882126340796e-19

R55_77 V55 V77 -11394.807194791281
L55_77 V55 V77 1.3856896645018015e-11
C55_77 V55 V77 -5.074127507870278e-22

R55_78 V55 V78 21749.635146631284
L55_78 V55 V78 -7.19836530500124e-12
C55_78 V55 V78 -1.5090697160063593e-19

R55_79 V55 V79 -9279.83345292571
L55_79 V55 V79 2.5414755830012042e-12
C55_79 V55 V79 1.1541200990171082e-19

R55_80 V55 V80 37521.750120975834
L55_80 V55 V80 4.314945566047216e-12
C55_80 V55 V80 3.015944200711869e-20

R55_81 V55 V81 -14315.912327784805
L55_81 V55 V81 -7.811457278768611e-12
C55_81 V55 V81 -3.4052088224562733e-20

R55_82 V55 V82 40057.68460982105
L55_82 V55 V82 3.1494915969568444e-12
C55_82 V55 V82 2.2696372968628386e-19

R55_83 V55 V83 6195.418425789797
L55_83 V55 V83 -2.2347719832789887e-12
C55_83 V55 V83 -3.856953686638393e-19

R55_84 V55 V84 6822.2793024045795
L55_84 V55 V84 3.3308107579606885e-12
C55_84 V55 V84 9.633759878585835e-20

R55_85 V55 V85 72275.88261116999
L55_85 V55 V85 4.091795387789782e-12
C55_85 V55 V85 1.474214535880833e-19

R55_86 V55 V86 5269.814702939607
L55_86 V55 V86 7.242041238998997e-12
C55_86 V55 V86 1.2384371328448577e-19

R55_87 V55 V87 2725.9190165680134
L55_87 V55 V87 -1.6660581763712488e-12
C55_87 V55 V87 -1.3848790431929135e-19

R55_88 V55 V88 -5936.610777560748
L55_88 V55 V88 -2.2291436159710126e-12
C55_88 V55 V88 -1.5518271641550545e-19

R55_89 V55 V89 -5561.108937225706
L55_89 V55 V89 -1.9724201492512827e-12
C55_89 V55 V89 -2.0104999138309727e-19

R55_90 V55 V90 -10195.628680134136
L55_90 V55 V90 -1.2426675805679896e-12
C55_90 V55 V90 -4.78139796957182e-19

R55_91 V55 V91 13044.672374301754
L55_91 V55 V91 7.172880874501404e-13
C55_91 V55 V91 5.435790823783897e-19

R55_92 V55 V92 2759.3198282861063
L55_92 V55 V92 2.2638855162641054e-12
C55_92 V55 V92 9.579695036067963e-20

R55_93 V55 V93 -269240.96232421405
L55_93 V55 V93 -9.228342158474675e-12
C55_93 V55 V93 -4.7594373046504803e-20

R55_94 V55 V94 -4206.011987543991
L55_94 V55 V94 5.143746881564948e-12
C55_94 V55 V94 1.5008723209690897e-19

R55_95 V55 V95 -1346.9468632905573
L55_95 V55 V95 7.346016812010073e-12
C55_95 V55 V95 3.2911498746844466e-20

R55_96 V55 V96 -11566.21837771947
L55_96 V55 V96 2.2960992613318085e-11
C55_96 V55 V96 1.0584770919941378e-19

R55_97 V55 V97 -3497.3609740821407
L55_97 V55 V97 1.4289110835069852e-12
C55_97 V55 V97 3.4610183057627975e-19

R55_98 V55 V98 2669.5737490060874
L55_98 V55 V98 1.7478568800612144e-12
C55_98 V55 V98 2.839934267634696e-19

R55_99 V55 V99 3206.143404073494
L55_99 V55 V99 -6.57229182193432e-13
C55_99 V55 V99 -6.3489912674856685e-19

R55_100 V55 V100 -2616.9852915818083
L55_100 V55 V100 -3.125246965358153e-12
C55_100 V55 V100 -1.9325675003795463e-19

R55_101 V55 V101 15524.41508425714
L55_101 V55 V101 -3.6782864039899235e-12
C55_101 V55 V101 -1.6580782518234393e-19

R55_102 V55 V102 2940191.6541162534
L55_102 V55 V102 -3.4871742432573103e-12
C55_102 V55 V102 -1.717606675915104e-19

R55_103 V55 V103 2314.9959450801916
L55_103 V55 V103 2.4049265267907624e-12
C55_103 V55 V103 2.4055209515364416e-19

R55_104 V55 V104 2168.7347606674543
L55_104 V55 V104 4.26082844696572e-12
C55_104 V55 V104 4.187102848459338e-20

R55_105 V55 V105 -11089.079945085621
L55_105 V55 V105 -1.6974052943461624e-12
C55_105 V55 V105 -1.5375454790091093e-19

R55_106 V55 V106 -22722.27416686696
L55_106 V55 V106 -1.661818521648155e-12
C55_106 V55 V106 -2.6363462857004644e-19

R55_107 V55 V107 -5766.061655104444
L55_107 V55 V107 1.0581022796921e-12
C55_107 V55 V107 3.116961349796455e-19

R55_108 V55 V108 5773.908296288918
L55_108 V55 V108 -1.0928298217416809e-11
C55_108 V55 V108 2.800123451447147e-20

R55_109 V55 V109 26900.597201319026
L55_109 V55 V109 5.090687143192228e-12
C55_109 V55 V109 2.4198019921562607e-19

R55_110 V55 V110 -38283.73624265845
L55_110 V55 V110 2.170196964431181e-12
C55_110 V55 V110 2.0541261465877047e-19

R55_111 V55 V111 3171.964617187176
L55_111 V55 V111 -1.1463098488369946e-10
C55_111 V55 V111 -7.642497876105226e-20

R55_112 V55 V112 -3734.1145746033594
L55_112 V55 V112 1.3004633711318404e-11
C55_112 V55 V112 2.4098084058418047e-20

R55_113 V55 V113 -6100.532879485258
L55_113 V55 V113 1.4703366210135596e-12
C55_113 V55 V113 9.063328644438432e-20

R55_114 V55 V114 -22038.364281094284
L55_114 V55 V114 1.7598483032963402e-12
C55_114 V55 V114 2.5512749411369273e-19

R55_115 V55 V115 -1762.7814427078877
L55_115 V55 V115 -9.592062109635378e-13
C55_115 V55 V115 -2.2922262742068794e-19

R55_116 V55 V116 -3794.537488802842
L55_116 V55 V116 -4.775799490724037e-12
C55_116 V55 V116 -1.6735473398197477e-20

R55_117 V55 V117 -2358.2842011239354
L55_117 V55 V117 -3.678226512458835e-12
C55_117 V55 V117 -1.7625741014455787e-19

R55_118 V55 V118 6431.960593527276
L55_118 V55 V118 -1.174444484897318e-12
C55_118 V55 V118 -3.713301755795354e-19

R55_119 V55 V119 1681.3055682262743
L55_119 V55 V119 7.913255359292042e-12
C55_119 V55 V119 -4.346181654866673e-20

R55_120 V55 V120 1992.6868422426066
L55_120 V55 V120 -6.943140132062939e-12
C55_120 V55 V120 -1.915215813152007e-19

R55_121 V55 V121 3188.5717116619057
L55_121 V55 V121 -1.7385340952667187e-12
C55_121 V55 V121 4.4874927587895785e-20

R55_122 V55 V122 16038.629470282545
L55_122 V55 V122 5.999460764794743e-12
C55_122 V55 V122 9.049642731883784e-20

R55_123 V55 V123 5771.372632392921
L55_123 V55 V123 1.083639155053174e-12
C55_123 V55 V123 3.852474127601218e-19

R55_124 V55 V124 -136111.9062841625
L55_124 V55 V124 1.840808592354038e-12
C55_124 V55 V124 2.659584015543681e-19

R55_125 V55 V125 2111.2770375119167
L55_125 V55 V125 3.33326981312509e-10
C55_125 V55 V125 -2.7352526219663894e-20

R55_126 V55 V126 6103.535203808722
L55_126 V55 V126 1.1510585715667157e-12
C55_126 V55 V126 2.1904930824514876e-19

R55_127 V55 V127 -1692.27991688592
L55_127 V55 V127 -8.336268681743316e-12
C55_127 V55 V127 -1.7941777979408208e-19

R55_128 V55 V128 -2656.138996456343
L55_128 V55 V128 2.6827234332919668e-11
C55_128 V55 V128 7.724571247308822e-20

R55_129 V55 V129 -1228.8336374152718
L55_129 V55 V129 1.3320526163684104e-12
C55_129 V55 V129 2.34678641462465e-19

R55_130 V55 V130 -2698.750605662579
L55_130 V55 V130 -1.5489907075682818e-12
C55_130 V55 V130 -2.0515726478525382e-19

R55_131 V55 V131 2390.1160041671724
L55_131 V55 V131 -2.0537922632187367e-12
C55_131 V55 V131 -8.134923898099172e-20

R55_132 V55 V132 2669.082250400944
L55_132 V55 V132 -1.2684102772909605e-12
C55_132 V55 V132 -3.4996190637665972e-19

R55_133 V55 V133 -4410.025552291494
L55_133 V55 V133 -3.2231478659747257e-12
C55_133 V55 V133 -1.957791765912535e-19

R55_134 V55 V134 2489.797237414431
L55_134 V55 V134 2.3061645565180064e-11
C55_134 V55 V134 7.078802809925595e-20

R55_135 V55 V135 30398.293031448677
L55_135 V55 V135 1.5259125893794346e-11
C55_135 V55 V135 3.7582625822918756e-19

R55_136 V55 V136 22583.838867411167
L55_136 V55 V136 9.889901760744571e-12
C55_136 V55 V136 1.4744144924790406e-19

R55_137 V55 V137 1269.7140781357411
L55_137 V55 V137 -1.824675175138394e-12
C55_137 V55 V137 -1.3177440896347912e-19

R55_138 V55 V138 -4775.792318706859
L55_138 V55 V138 2.5037625099018932e-12
C55_138 V55 V138 8.430138824765039e-20

R55_139 V55 V139 24855.387324792337
L55_139 V55 V139 -3.797460391381884e-12
C55_139 V55 V139 -5.638996729037882e-19

R55_140 V55 V140 -7531.028072350232
L55_140 V55 V140 2.0020794342940075e-12
C55_140 V55 V140 -8.988312259757804e-20

R55_141 V55 V141 3292.7726727243958
L55_141 V55 V141 2.171132828666779e-12
C55_141 V55 V141 3.6093014559476427e-19

R55_142 V55 V142 -2754.98909678331
L55_142 V55 V142 1.7628353716288257e-11
C55_142 V55 V142 -4.184344655024802e-20

R55_143 V55 V143 9120.696477036496
L55_143 V55 V143 9.437902521096663e-13
C55_143 V55 V143 2.1159128326153032e-19

R55_144 V55 V144 3247.2353433417265
L55_144 V55 V144 -3.798508508597133e-12
C55_144 V55 V144 4.4210175372211215e-20

R55_145 V55 V145 -862.8535382876352
L55_145 V55 V145 1.6640523541124513e-12
C55_145 V55 V145 1.3593345516234863e-19

R55_146 V55 V146 10158.311208553037
L55_146 V55 V146 -2.803356708407666e-12
C55_146 V55 V146 -6.003794045809395e-20

R55_147 V55 V147 -699.3604368185415
L55_147 V55 V147 -2.592903290158828e-12
C55_147 V55 V147 3.487875331681763e-19

R55_148 V55 V148 -1315.8826025308917
L55_148 V55 V148 1.957688110813657e-12
C55_148 V55 V148 9.883804993100352e-20

R55_149 V55 V149 13815.617886674881
L55_149 V55 V149 -8.126312272938117e-13
C55_149 V55 V149 -5.847297757594401e-19

R55_150 V55 V150 1024.656998358355
L55_150 V55 V150 2.4902091942613368e-11
C55_150 V55 V150 2.5027246725573214e-19

R55_151 V55 V151 426.0495346347457
L55_151 V55 V151 -8.302665310532385e-13
C55_151 V55 V151 -1.9536436397711565e-19

R55_152 V55 V152 4384.911661787568
L55_152 V55 V152 4.58654112284082e-12
C55_152 V55 V152 -2.946201322782438e-21

R55_153 V55 V153 1518.3142660143958
L55_153 V55 V153 -6.096052302114567e-12
C55_153 V55 V153 -1.1054609995580592e-20

R55_154 V55 V154 13255.89279584222
L55_154 V55 V154 -2.7702452361146014e-11
C55_154 V55 V154 -1.4812855468184387e-19

R55_155 V55 V155 -309.29190256154203
L55_155 V55 V155 -1.6338755704674785e-12
C55_155 V55 V155 -3.4607769917929163e-19

R55_156 V55 V156 2570.8572582129796
L55_156 V55 V156 -6.156501180448977e-12
C55_156 V55 V156 -1.1998538347019765e-19

R55_157 V55 V157 6700.175065265152
L55_157 V55 V157 1.3109694855490242e-12
C55_157 V55 V157 4.961563920381996e-19

R55_158 V55 V158 -3319.8808466730025
L55_158 V55 V158 -5.008285562219214e-12
C55_158 V55 V158 -5.3589847211039607e-20

R55_159 V55 V159 1921.84421541923
L55_159 V55 V159 4.761722006861694e-13
C55_159 V55 V159 2.0782304287323714e-19

R55_160 V55 V160 3924.4963052833546
L55_160 V55 V160 -1.2533601051214293e-12
C55_160 V55 V160 -1.0232134084566117e-20

R55_161 V55 V161 -2689.539577580135
L55_161 V55 V161 2.3493455831743462e-11
C55_161 V55 V161 -2.4521224290064945e-20

R55_162 V55 V162 -5086.7817858086
L55_162 V55 V162 -2.762717341043946e-12
C55_162 V55 V162 -8.486517496583922e-20

R55_163 V55 V163 2266.176443684071
L55_163 V55 V163 3.548304419874689e-12
C55_163 V55 V163 -3.2251929225221463e-21

R55_164 V55 V164 -3451.7900163113004
L55_164 V55 V164 1.5120886565951828e-12
C55_164 V55 V164 -2.6507352873287998e-20

R55_165 V55 V165 -1971.3680939051512
L55_165 V55 V165 -2.556105067580575e-12
C55_165 V55 V165 -2.241534077800138e-19

R55_166 V55 V166 2336.387764181886
L55_166 V55 V166 1.994967950952759e-12
C55_166 V55 V166 1.0672428340259734e-19

R55_167 V55 V167 1052.2751127514196
L55_167 V55 V167 -5.303414987126149e-13
C55_167 V55 V167 -4.031415840824618e-20

R55_168 V55 V168 -5758.779243063663
L55_168 V55 V168 3.474435130791823e-12
C55_168 V55 V168 4.7870300634825604e-20

R55_169 V55 V169 2071.2559148227665
L55_169 V55 V169 8.285223836247055e-12
C55_169 V55 V169 1.60506461922753e-19

R55_170 V55 V170 -3353.5774028629985
L55_170 V55 V170 -4.231672467484539e-12
C55_170 V55 V170 -1.3029642293742202e-19

R55_171 V55 V171 -633.3641611284373
L55_171 V55 V171 8.434118737577157e-12
C55_171 V55 V171 -5.301170318525554e-20

R55_172 V55 V172 -6834.708915978025
L55_172 V55 V172 -3.1391462635062182e-12
C55_172 V55 V172 -4.065123637955236e-20

R55_173 V55 V173 -4307.774483947608
L55_173 V55 V173 8.078859827808929e-12
C55_173 V55 V173 -2.9482680809577105e-20

R55_174 V55 V174 -6784.466118915579
L55_174 V55 V174 -2.5738345111628003e-12
C55_174 V55 V174 1.0655333961431151e-19

R55_175 V55 V175 2701.4615470196695
L55_175 V55 V175 1.2571576453826168e-12
C55_175 V55 V175 -2.1059271179840286e-19

R55_176 V55 V176 -11234.216908365463
L55_176 V55 V176 -1.0549116314676283e-11
C55_176 V55 V176 -1.104986918062203e-19

R55_177 V55 V177 4890.105202593778
L55_177 V55 V177 8.968549114374525e-12
C55_177 V55 V177 2.6533650456547898e-21

R55_178 V55 V178 2034.4560680543843
L55_178 V55 V178 1.6970537808990994e-12
C55_178 V55 V178 9.384709436556692e-20

R55_179 V55 V179 -2010.8620617335941
L55_179 V55 V179 -4.770499425627265e-11
C55_179 V55 V179 2.7559580310370127e-19

R55_180 V55 V180 1737.3823962701401
L55_180 V55 V180 2.2424768436737507e-12
C55_180 V55 V180 2.2096399544753193e-19

R55_181 V55 V181 13322.91528802345
L55_181 V55 V181 -3.921941711466419e-12
C55_181 V55 V181 3.723630880180104e-20

R55_182 V55 V182 -2298.733830235663
L55_182 V55 V182 -2.1313012908249574e-12
C55_182 V55 V182 -1.5865144284226003e-19

R55_183 V55 V183 936.2109204398752
L55_183 V55 V183 1.4162983716962364e-11
C55_183 V55 V183 5.029232758057031e-20

R55_184 V55 V184 -5246.497406877061
L55_184 V55 V184 6.638279871765497e-12
C55_184 V55 V184 8.667085521309242e-21

R55_185 V55 V185 -2469.91841354068
L55_185 V55 V185 -8.792501157612799e-12
C55_185 V55 V185 -5.376024727208244e-20

R55_186 V55 V186 -4411.2566977052875
L55_186 V55 V186 -3.4341915390889736e-12
C55_186 V55 V186 6.515290776025832e-20

R55_187 V55 V187 -2310.746895218522
L55_187 V55 V187 -1.8658811498197913e-12
C55_187 V55 V187 -2.6855085171776567e-19

R55_188 V55 V188 -1351.3067536400079
L55_188 V55 V188 -1.2297102741796537e-12
C55_188 V55 V188 -1.924103621637885e-19

R55_189 V55 V189 1997.9113572680133
L55_189 V55 V189 3.1443315836610583e-12
C55_189 V55 V189 -1.3735220036342987e-20

R55_190 V55 V190 2239.353353579766
L55_190 V55 V190 4.491435613437449e-12
C55_190 V55 V190 1.107781807657974e-19

R55_191 V55 V191 -1447.2735452846687
L55_191 V55 V191 3.5938466010228806e-11
C55_191 V55 V191 5.9842420661839e-20

R55_192 V55 V192 5560.334897161376
L55_192 V55 V192 7.768222552647247e-12
C55_192 V55 V192 3.433449247810502e-20

R55_193 V55 V193 -9175.778475108626
L55_193 V55 V193 4.1848703133169775e-11
C55_193 V55 V193 6.545393892141809e-20

R55_194 V55 V194 34804.621736220375
L55_194 V55 V194 2.750442688377398e-12
C55_194 V55 V194 1.155861572466867e-19

R55_195 V55 V195 1221.1346338695635
L55_195 V55 V195 4.101194689605983e-12
C55_195 V55 V195 -3.985525409872423e-20

R55_196 V55 V196 1146.9683961007004
L55_196 V55 V196 1.6709502469668753e-12
C55_196 V55 V196 1.3659766192984276e-19

R55_197 V55 V197 -433475.0135255141
L55_197 V55 V197 -1.2638845098620151e-11
C55_197 V55 V197 6.23394541852392e-20

R55_198 V55 V198 -7338.221649355404
L55_198 V55 V198 -4.914013627514999e-12
C55_198 V55 V198 -3.8726055907140084e-20

R55_199 V55 V199 -4332.860121116681
L55_199 V55 V199 -5.226662973478723e-12
C55_199 V55 V199 5.547782264898718e-20

R55_200 V55 V200 -3544.819232822922
L55_200 V55 V200 -5.216613955098915e-12
C55_200 V55 V200 -1.7125266619628987e-20

R56_56 V56 0 -217.5856770726981
L56_56 V56 0 -4.442355745557017e-13
C56_56 V56 0 -3.0821755083506386e-18

R56_57 V56 V57 -15354.377187029346
L56_57 V56 V57 -3.1571402350844025e-11
C56_57 V56 V57 2.063247241284927e-21

R56_58 V56 V58 2541.3701841236407
L56_58 V56 V58 -6.060911043754497e-11
C56_58 V56 V58 -4.1228667033973e-21

R56_59 V56 V59 332657.04309645627
L56_59 V56 V59 4.254107957706671e-11
C56_59 V56 V59 9.726359248160255e-20

R56_60 V56 V60 -4005.457492353126
L56_60 V56 V60 6.341066533007243e-13
C56_60 V56 V60 7.975989400617811e-19

R56_61 V56 V61 3963.390172085228
L56_61 V56 V61 2.7160203166831337e-12
C56_61 V56 V61 2.0143801531050702e-19

R56_62 V56 V62 -7539.561817593501
L56_62 V56 V62 2.1190868144386817e-12
C56_62 V56 V62 3.154756067750773e-19

R56_63 V56 V63 7390.976879207141
L56_63 V56 V63 -7.179891366624287e-12
C56_63 V56 V63 -1.1549642258329682e-19

R56_64 V56 V64 2474.915833655399
L56_64 V56 V64 7.860240075178974e-13
C56_64 V56 V64 7.412825530662667e-19

R56_65 V56 V65 25105.70913778317
L56_65 V56 V65 7.250557176174464e-12
C56_65 V56 V65 1.5476623793997585e-19

R56_66 V56 V66 12721.957098639172
L56_66 V56 V66 9.733817908107637e-12
C56_66 V56 V66 1.2157285034630631e-19

R56_67 V56 V67 -12583.270453722145
L56_67 V56 V67 -1.5887064497367793e-11
C56_67 V56 V67 -3.172655806615285e-20

R56_68 V56 V68 1638.3460387155278
L56_68 V56 V68 -1.4561750398407207e-12
C56_68 V56 V68 -5.26768814154699e-19

R56_69 V56 V69 -3257.769937474644
L56_69 V56 V69 -1.6067282465344862e-12
C56_69 V56 V69 -3.662363990994128e-19

R56_70 V56 V70 15329.500641942379
L56_70 V56 V70 -2.7159553944390786e-12
C56_70 V56 V70 -2.5435700770546045e-19

R56_71 V56 V71 6534.3902709279455
L56_71 V56 V71 2.306710886394623e-12
C56_71 V56 V71 2.0622773983760068e-19

R56_72 V56 V72 2245.462136203711
L56_72 V56 V72 -7.538875490868793e-12
C56_72 V56 V72 -1.5609078474990626e-19

R56_73 V56 V73 9666.416078227288
L56_73 V56 V73 3.433089634307784e-12
C56_73 V56 V73 2.1055879233208363e-19

R56_74 V56 V74 -5197.207025764876
L56_74 V56 V74 -2.565159460810585e-11
C56_74 V56 V74 2.653868381009475e-20

R56_75 V56 V75 7637.604993446042
L56_75 V56 V75 -1.46349443707266e-11
C56_75 V56 V75 5.2648329431992406e-20

R56_76 V56 V76 -684.2236542649846
L56_76 V56 V76 -1.4400623615264789e-12
C56_76 V56 V76 -7.763636656982523e-20

R56_77 V56 V77 -5558.099411491403
L56_77 V56 V77 5.580791581157907e-11
C56_77 V56 V77 4.076398581779068e-20

R56_78 V56 V78 4251.553462359562
L56_78 V56 V78 -7.689673922359483e-12
C56_78 V56 V78 -2.0071069595687577e-19

R56_79 V56 V79 -2900.437110694614
L56_79 V56 V79 -3.698419326388976e-12
C56_79 V56 V79 -1.652501542013963e-19

R56_80 V56 V80 2691.3666598093446
L56_80 V56 V80 7.94595567362063e-13
C56_80 V56 V80 4.208323166716109e-19

R56_81 V56 V81 4173.528850584604
L56_81 V56 V81 6.601174640460443e-12
C56_81 V56 V81 1.1841957383237603e-19

R56_82 V56 V82 -51342.55478800886
L56_82 V56 V82 1.9620511256676615e-12
C56_82 V56 V82 4.0069958235158524e-19

R56_83 V56 V83 6468.8126890795365
L56_83 V56 V83 5.390237961710499e-12
C56_83 V56 V83 7.845885330960096e-20

R56_84 V56 V84 2483.631857249745
L56_84 V56 V84 2.581409047444156e-08
C56_84 V56 V84 -1.6600344548046756e-19

R56_85 V56 V85 -34588.181258922545
L56_85 V56 V85 2.494842755548677e-12
C56_85 V56 V85 2.205272984395397e-19

R56_86 V56 V86 3253.44307912144
L56_86 V56 V86 3.921527331057958e-12
C56_86 V56 V86 2.209387140951582e-19

R56_87 V56 V87 84934.16001640544
L56_87 V56 V87 -2.5479472713654818e-12
C56_87 V56 V87 -1.4763013374211246e-19

R56_88 V56 V88 2598.942407170507
L56_88 V56 V88 -8.158330981208966e-13
C56_88 V56 V88 -4.819598909723995e-19

R56_89 V56 V89 -2891.6391721536334
L56_89 V56 V89 -1.100721734698933e-12
C56_89 V56 V89 -4.151639768946583e-19

R56_90 V56 V90 -4287.893172212191
L56_90 V56 V90 -7.14550299821408e-13
C56_90 V56 V90 -8.252844790042697e-19

R56_91 V56 V91 1613.6907687534047
L56_91 V56 V91 1.0751046464116463e-12
C56_91 V56 V91 3.713674701034091e-19

R56_92 V56 V92 11359.488480634998
L56_92 V56 V92 5.62748127644199e-13
C56_92 V56 V92 6.491828247527081e-19

R56_93 V56 V93 3315.303247684144
L56_93 V56 V93 -7.472094791852937e-12
C56_93 V56 V93 -3.583877268782493e-20

R56_94 V56 V94 -3003.3983581735606
L56_94 V56 V94 2.6510559676131337e-12
C56_94 V56 V94 3.1728357540867726e-19

R56_95 V56 V95 -2942.1689639619467
L56_95 V56 V95 1.3835748395590684e-11
C56_95 V56 V95 1.2057352619491641e-19

R56_96 V56 V96 -575.3962892726573
L56_96 V56 V96 -2.0617915474325846e-11
C56_96 V56 V96 1.4660300446014872e-19

R56_97 V56 V97 -1983.612841851092
L56_97 V56 V97 8.849714153576355e-13
C56_97 V56 V97 6.937913797567318e-19

R56_98 V56 V98 1524.7652097627335
L56_98 V56 V98 9.60598704860479e-13
C56_98 V56 V98 5.29545029903293e-19

R56_99 V56 V99 -1992.2726277074537
L56_99 V56 V99 -8.323890210997016e-13
C56_99 V56 V99 -5.288388707707163e-19

R56_100 V56 V100 753.5186342804516
L56_100 V56 V100 -7.674397595974097e-13
C56_100 V56 V100 -8.53225896222236e-19

R56_101 V56 V101 11168.927605665356
L56_101 V56 V101 -2.4680570311579212e-12
C56_101 V56 V101 -2.6050912868279324e-19

R56_102 V56 V102 -13357.026940052607
L56_102 V56 V102 -1.723834899336234e-12
C56_102 V56 V102 -3.6015404918649774e-19

R56_103 V56 V103 1491.8429147254171
L56_103 V56 V103 2.367036979700363e-12
C56_103 V56 V103 1.131887081441109e-19

R56_104 V56 V104 1312.3227578317249
L56_104 V56 V104 1.886189235375926e-12
C56_104 V56 V104 3.53258336549101e-19

R56_105 V56 V105 3034.740188299693
L56_105 V56 V105 -1.246648721652014e-12
C56_105 V56 V105 -2.8570276677983605e-19

R56_106 V56 V106 3737.9937747472386
L56_106 V56 V106 -1.1804471711683878e-12
C56_106 V56 V106 -3.907610572648187e-19

R56_107 V56 V107 3537.949281128646
L56_107 V56 V107 1.4245132385402113e-12
C56_107 V56 V107 3.8710591303751696e-19

R56_108 V56 V108 -1025.044015776815
L56_108 V56 V108 2.24899756765715e-12
C56_108 V56 V108 1.6733262994192895e-19

R56_109 V56 V109 -2939.352207798815
L56_109 V56 V109 2.463533471901056e-12
C56_109 V56 V109 4.840537158433218e-19

R56_110 V56 V110 -1810.8057527993515
L56_110 V56 V110 1.7698003143091528e-12
C56_110 V56 V110 2.6034633433994484e-19

R56_111 V56 V111 -6468.902617131498
L56_111 V56 V111 -1.0909138298431016e-11
C56_111 V56 V111 -7.280293887045633e-20

R56_112 V56 V112 1438.1750288682722
L56_112 V56 V112 2.114891174313327e-12
C56_112 V56 V112 2.0219708713350814e-19

R56_113 V56 V113 -10108.097601554391
L56_113 V56 V113 1.1445938207961727e-12
C56_113 V56 V113 1.2452630378968302e-19

R56_114 V56 V114 -4597.505969806851
L56_114 V56 V114 1.1808007135620046e-12
C56_114 V56 V114 4.2778426191926114e-19

R56_115 V56 V115 -1136.6823995845402
L56_115 V56 V115 -1.2218956702660738e-12
C56_115 V56 V115 -2.733879962584968e-19

R56_116 V56 V116 -1120.8073300295184
L56_116 V56 V116 -8.203002749776393e-13
C56_116 V56 V116 -2.5011030155179777e-19

R56_117 V56 V117 -1452.76001173525
L56_117 V56 V117 -1.6887376254713158e-12
C56_117 V56 V117 -3.2566053679877364e-19

R56_118 V56 V118 1142.6988480266916
L56_118 V56 V118 -8.103114669856679e-13
C56_118 V56 V118 -5.973470932832324e-19

R56_119 V56 V119 1241.1659500705775
L56_119 V56 V119 -6.434834487953754e-12
C56_119 V56 V119 -2.2764708072627375e-19

R56_120 V56 V120 654.9780366102477
L56_120 V56 V120 6.371116425505333e-11
C56_120 V56 V120 -4.901619290378223e-19

R56_121 V56 V121 2415.0316456065443
L56_121 V56 V121 -1.680829681777832e-12
C56_121 V56 V121 1.1226730285502329e-19

R56_122 V56 V122 -7956.90722252583
L56_122 V56 V122 3.913255592810502e-12
C56_122 V56 V122 8.738551655503784e-20

R56_123 V56 V123 4764.683482463519
L56_123 V56 V123 1.247875538152079e-12
C56_123 V56 V123 3.3380172119415695e-19

R56_124 V56 V124 -4607.361713171612
L56_124 V56 V124 6.624491115279247e-13
C56_124 V56 V124 1.045723536449711e-18

R56_125 V56 V125 760.8313052919277
L56_125 V56 V125 4.4451459652853615e-12
C56_125 V56 V125 -1.1003892255919992e-20

R56_126 V56 V126 41039.359104453266
L56_126 V56 V126 7.946329903060951e-13
C56_126 V56 V126 3.3951156230239164e-19

R56_127 V56 V127 -1335.2154782545172
L56_127 V56 V127 2.852072350499882e-12
C56_127 V56 V127 2.2773853494161074e-19

R56_128 V56 V128 -666.1810966564567
L56_128 V56 V128 -3.3538902626177324e-12
C56_128 V56 V128 -1.2499631538218662e-19

R56_129 V56 V129 -536.810397962181
L56_129 V56 V129 1.1263253176136956e-12
C56_129 V56 V129 4.1676844858781127e-19

R56_130 V56 V130 -1638.8003151981109
L56_130 V56 V130 -9.311705199541555e-13
C56_130 V56 V130 -3.8618354517701165e-19

R56_131 V56 V131 1249.7846116949709
L56_131 V56 V131 -1.209331868122972e-12
C56_131 V56 V131 -3.9737183497735754e-19

R56_132 V56 V132 612.7660681553009
L56_132 V56 V132 -8.385199851098572e-13
C56_132 V56 V132 -6.892319730639321e-19

R56_133 V56 V133 -2422.451945877165
L56_133 V56 V133 -1.6725798597179206e-12
C56_133 V56 V133 -4.621701314635656e-19

R56_134 V56 V134 957.8211774543379
L56_134 V56 V134 1.5037202777694285e-11
C56_134 V56 V134 -3.6714002934887056e-21

R56_135 V56 V135 -24268.07699662014
L56_135 V56 V135 -2.0636868818914882e-11
C56_135 V56 V135 -5.638182486973222e-20

R56_136 V56 V136 3682.301726140074
L56_136 V56 V136 2.440050443184303e-12
C56_136 V56 V136 9.009243240096404e-19

R56_137 V56 V137 593.3027202819192
L56_137 V56 V137 -1.2202315605974873e-12
C56_137 V56 V137 -1.8527219716885688e-19

R56_138 V56 V138 -1508.3271726350056
L56_138 V56 V138 1.6955817467161945e-12
C56_138 V56 V138 2.025670708328338e-19

R56_139 V56 V139 -1230.6905155116658
L56_139 V56 V139 6.332932256535921e-12
C56_139 V56 V139 8.607253795636417e-21

R56_140 V56 V140 4878.642975219191
L56_140 V56 V140 2.0221416421894326e-11
C56_140 V56 V140 -9.386212719400568e-19

R56_141 V56 V141 1871.3516889800733
L56_141 V56 V141 9.502606564052105e-13
C56_141 V56 V141 6.901318838494803e-19

R56_142 V56 V142 -908.151820549828
L56_142 V56 V142 1.692350225047654e-11
C56_142 V56 V142 -4.3909127646203164e-20

R56_143 V56 V143 1452.9670811374433
L56_143 V56 V143 3.0820860495268208e-12
C56_143 V56 V143 1.8183664054969071e-19

R56_144 V56 V144 -449.0827492019265
L56_144 V56 V144 1.9134852615533983e-12
C56_144 V56 V144 1.5234098036998525e-19

R56_145 V56 V145 -447.2847275505715
L56_145 V56 V145 1.199899630250633e-12
C56_145 V56 V145 1.8091659668952997e-19

R56_146 V56 V146 4732.147017888763
L56_146 V56 V146 -2.4340004424671055e-12
C56_146 V56 V146 -1.432417195459711e-19

R56_147 V56 V147 -886.9281633952313
L56_147 V56 V147 3.7282086601872e-12
C56_147 V56 V147 2.1166195906376475e-19

R56_148 V56 V148 319.25784133507165
L56_148 V56 V148 2.0317505349016577e-12
C56_148 V56 V148 7.439738044126121e-19

R56_149 V56 V149 -13460.251899774486
L56_149 V56 V149 -5.107016730090326e-13
C56_149 V56 V149 -8.935380715124939e-19

R56_150 V56 V150 419.3109256833572
L56_150 V56 V150 1.3097035985218276e-11
C56_150 V56 V150 5.378698692167625e-19

R56_151 V56 V151 1733.407261963847
L56_151 V56 V151 1.339799834145017e-10
C56_151 V56 V151 -1.3506920240602517e-19

R56_152 V56 V152 -1379.9923437915484
L56_152 V56 V152 -7.777977058030987e-13
C56_152 V56 V152 -2.353764694166425e-19

R56_153 V56 V153 919.1882440379723
L56_153 V56 V153 -1.539620588330763e-12
C56_153 V56 V153 -1.265425784150689e-19

R56_154 V56 V154 -1137.9963813760257
L56_154 V56 V154 -5.077280081416554e-12
C56_154 V56 V154 -2.7277926999756085e-19

R56_155 V56 V155 -621.9704269662387
L56_155 V56 V155 -9.809897541917078e-13
C56_155 V56 V155 -2.4121433052557054e-19

R56_156 V56 V156 468.82317013588363
L56_156 V56 V156 -2.9303394198889995e-12
C56_156 V56 V156 -5.403043787491594e-19

R56_157 V56 V157 770.6210304768974
L56_157 V56 V157 5.849543026497728e-13
C56_157 V56 V157 9.735771485260518e-19

R56_158 V56 V158 6087.2572759957575
L56_158 V56 V158 -5.919218483754882e-12
C56_158 V56 V158 -6.474752241016645e-20

R56_159 V56 V159 468.7575308903347
L56_159 V56 V159 -2.306268400120435e-12
C56_159 V56 V159 1.7089381256829386e-20

R56_160 V56 V160 -321.89650339942386
L56_160 V56 V160 5.432678994295313e-13
C56_160 V56 V160 2.174196495855644e-19

R56_161 V56 V161 -854.4200829896332
L56_161 V56 V161 -7.489146502302376e-12
C56_161 V56 V161 -4.0065733742693346e-20

R56_162 V56 V162 -2442.201806955719
L56_162 V56 V162 -1.6801506943688913e-12
C56_162 V56 V162 -1.1387305690009412e-19

R56_163 V56 V163 -8149.556342733722
L56_163 V56 V163 1.2486524028851932e-12
C56_163 V56 V163 1.5744726752763273e-19

R56_164 V56 V164 360.9884807381771
L56_164 V56 V164 7.251175918566499e-12
C56_164 V56 V164 -1.6148329007732832e-19

R56_165 V56 V165 4638.039741160199
L56_165 V56 V165 -1.7201067009687577e-12
C56_165 V56 V165 -3.044046760036749e-19

R56_166 V56 V166 703.9123030750674
L56_166 V56 V166 1.3195745417976013e-12
C56_166 V56 V166 2.8632252688139645e-19

R56_167 V56 V167 1315.2856895460186
L56_167 V56 V167 2.0560067775396383e-12
C56_167 V56 V167 2.457822182152521e-21

R56_168 V56 V168 -583.6911986551494
L56_168 V56 V168 -4.549123325599491e-13
C56_168 V56 V168 1.172434632793298e-19

R56_169 V56 V169 1251.0136564447705
L56_169 V56 V169 2.6379700396984712e-11
C56_169 V56 V169 2.7712469518369395e-19

R56_170 V56 V170 -1414.665213599578
L56_170 V56 V170 -1.567403005960321e-12
C56_170 V56 V170 -2.396156325108412e-19

R56_171 V56 V171 -764.5809201686307
L56_171 V56 V171 -7.419069363515146e-13
C56_171 V56 V171 -1.9945681052367473e-19

R56_172 V56 V172 -4292.681660424914
L56_172 V56 V172 1.1016654119959312e-12
C56_172 V56 V172 -9.920386112435986e-20

R56_173 V56 V173 -2210.9588693033393
L56_173 V56 V173 5.726742167091156e-12
C56_173 V56 V173 -7.834921428596183e-20

R56_174 V56 V174 -1024.4667509758365
L56_174 V56 V174 -3.038298805378959e-12
C56_174 V56 V174 1.6013358434533191e-19

R56_175 V56 V175 1545.824756134837
L56_175 V56 V175 -2.3182260512446258e-11
C56_175 V56 V175 -1.4930187150956725e-19

R56_176 V56 V176 2993.0802310268205
L56_176 V56 V176 -5.886771466165153e-10
C56_176 V56 V176 -5.05562372173503e-19

R56_177 V56 V177 1959.5813289541813
L56_177 V56 V177 4.030017290002061e-12
C56_177 V56 V177 4.8700490117163363e-20

R56_178 V56 V178 801.9932898839902
L56_178 V56 V178 1.0318340550808153e-12
C56_178 V56 V178 1.277683565993123e-19

R56_179 V56 V179 5884.913885554326
L56_179 V56 V179 8.869651549388779e-13
C56_179 V56 V179 4.0861429963277146e-19

R56_180 V56 V180 21175.245848286195
L56_180 V56 V180 1.6462161031475729e-12
C56_180 V56 V180 5.796547865095404e-19

R56_181 V56 V181 -13019.55241680291
L56_181 V56 V181 -3.3706645215823493e-12
C56_181 V56 V181 1.1128618998580945e-19

R56_182 V56 V182 -1279.0520075002323
L56_182 V56 V182 -1.1878857078197996e-12
C56_182 V56 V182 -1.931482906019176e-19

R56_183 V56 V183 3275.1473276883
L56_183 V56 V183 1.7738489627282917e-12
C56_183 V56 V183 1.1638886362917436e-19

R56_184 V56 V184 1225.9926536342045
L56_184 V56 V184 5.494375777736453e-12
C56_184 V56 V184 -1.0851649856691767e-19

R56_185 V56 V185 -6005.280259812766
L56_185 V56 V185 -2.208612159409991e-11
C56_185 V56 V185 -1.2439862877061524e-19

R56_186 V56 V186 -10501.9811781588
L56_186 V56 V186 -6.221704950778083e-12
C56_186 V56 V186 4.096058844769185e-20

R56_187 V56 V187 -2827.744734672116
L56_187 V56 V187 -1.1312139037942337e-12
C56_187 V56 V187 -4.2732974053491603e-19

R56_188 V56 V188 -363.6488488608644
L56_188 V56 V188 -5.658924314941161e-13
C56_188 V56 V188 -2.664255815739963e-19

R56_189 V56 V189 1981.1637470885692
L56_189 V56 V189 5.960702800731043e-12
C56_189 V56 V189 -8.197939038378446e-20

R56_190 V56 V190 1044.7694905611118
L56_190 V56 V190 3.491571848761823e-12
C56_190 V56 V190 2.2937197834773106e-19

R56_191 V56 V191 -1981.277981536754
L56_191 V56 V191 -9.776381354225922e-13
C56_191 V56 V191 -1.0460764333931331e-19

R56_192 V56 V192 2404.726973600048
L56_192 V56 V192 9.784118136395834e-13
C56_192 V56 V192 1.6777901657866807e-19

R56_193 V56 V193 -1265.3247500116613
L56_193 V56 V193 1.1835145101573046e-11
C56_193 V56 V193 1.3412666788686389e-19

R56_194 V56 V194 2893.8829319078463
L56_194 V56 V194 1.7603265171562177e-12
C56_194 V56 V194 2.685168815668234e-19

R56_195 V56 V195 903.0160803488449
L56_195 V56 V195 6.191224936896657e-13
C56_195 V56 V195 5.370338895677593e-19

R56_196 V56 V196 544.6753300953895
L56_196 V56 V196 -6.043966862272014e-12
C56_196 V56 V196 -3.1047097486996824e-19

R56_197 V56 V197 -18649.758204825306
L56_197 V56 V197 6.596029130938455e-12
C56_197 V56 V197 6.319521237435729e-20

R56_198 V56 V198 10221.518282589686
L56_198 V56 V198 -3.203466265841636e-12
C56_198 V56 V198 4.4162057833537353e-20

R56_199 V56 V199 847.5374914502135
L56_199 V56 V199 2.6717825378312824e-11
C56_199 V56 V199 9.514862519722932e-20

R56_200 V56 V200 -499.03104105775526
L56_200 V56 V200 -5.228455372789151e-12
C56_200 V56 V200 9.276812057428678e-20

R57_57 V57 0 10343.926131642578
L57_57 V57 0 -2.5105853148297534e-13
C57_57 V57 0 -8.2719125200764e-20

R57_58 V57 V58 -50096.867390723215
L57_58 V57 V58 -3.2639391712042494e-12
C57_58 V57 V58 -1.2943300985614142e-19

R57_59 V57 V59 -11563.677734033765
L57_59 V57 V59 -2.180559610345761e-12
C57_59 V57 V59 -2.286266725903139e-19

R57_60 V57 V60 -7533.858304392019
L57_60 V57 V60 -1.5134375360278106e-12
C57_60 V57 V60 -2.516705758244653e-19

R57_61 V57 V61 2072.2453595372594
L57_61 V57 V61 1.285588726668539e-12
C57_61 V57 V61 4.627155153729581e-19

R57_62 V57 V62 -13696.232680166417
L57_62 V57 V62 -1.4074101958067902e-11
C57_62 V57 V62 -4.5355797585936226e-20

R57_63 V57 V63 -35150.454027947024
L57_63 V57 V63 -1.4131900455140251e-11
C57_63 V57 V63 5.388659114881583e-20

R57_64 V57 V64 41036.565589439924
L57_64 V57 V64 1.78835114074116e-11
C57_64 V57 V64 1.0540691312871378e-19

R57_65 V57 V65 4692.4513089117545
L57_65 V57 V65 1.6231651779436546e-12
C57_65 V57 V65 3.095034474793398e-19

R57_66 V57 V66 -22112.210552716497
L57_66 V57 V66 1.8372735197754653e-11
C57_66 V57 V66 7.568324308045214e-21

R57_67 V57 V67 28335.27585098054
L57_67 V57 V67 4.054700399666495e-12
C57_67 V57 V67 1.3365521213433722e-19

R57_68 V57 V68 8603.909642405539
L57_68 V57 V68 2.312117838298223e-12
C57_68 V57 V68 2.1290274695080966e-19

R57_69 V57 V69 -2151.818510382596
L57_69 V57 V69 1.809787129892172e-12
C57_69 V57 V69 -1.9067238652649748e-20

R57_70 V57 V70 6014.608064671653
L57_70 V57 V70 3.895249109205802e-12
C57_70 V57 V70 1.5918905706256336e-19

R57_71 V57 V71 4649.873756040847
L57_71 V57 V71 9.774437223039904e-12
C57_71 V57 V71 -1.3143843176848576e-20

R57_72 V57 V72 4526.45433438018
L57_72 V57 V72 9.543750911106076e-12
C57_72 V57 V72 -2.9843021764424655e-20

R57_73 V57 V73 1813.788004368278
L57_73 V57 V73 -5.230618262426704e-10
C57_73 V57 V73 -1.4681371324287512e-19

R57_74 V57 V74 11898.925453263044
L57_74 V57 V74 -1.3707649721844753e-11
C57_74 V57 V74 -1.4771977777824662e-19

R57_75 V57 V75 -13729.259433749852
L57_75 V57 V75 -9.21188411453977e-12
C57_75 V57 V75 -7.151807241478395e-20

R57_76 V57 V76 -5304.983390655579
L57_76 V57 V76 -3.7761059792358e-12
C57_76 V57 V76 -5.2479715421200384e-20

R57_77 V57 V77 13396.502629919069
L57_77 V57 V77 -7.45052125952817e-13
C57_77 V57 V77 -4.686563836817352e-19

R57_78 V57 V78 -2990.9046620683584
L57_78 V57 V78 -9.383018781452738e-12
C57_78 V57 V78 4.5911451544595924e-20

R57_79 V57 V79 -2196.479667086099
L57_79 V57 V79 -4.740180032869537e-12
C57_79 V57 V79 -3.866601395052803e-20

R57_80 V57 V80 -2139.96882105839
L57_80 V57 V80 -3.606284372664022e-12
C57_80 V57 V80 -7.197264850896195e-20

R57_81 V57 V81 -1072.2583468855817
L57_81 V57 V81 1.0321189985895703e-12
C57_81 V57 V81 4.2139328541561543e-19

R57_82 V57 V82 9322.713495341275
L57_82 V57 V82 -1.570086052073109e-11
C57_82 V57 V82 -9.18395466898164e-20

R57_83 V57 V83 2530.791087677871
L57_83 V57 V83 -1.3896558962213932e-11
C57_83 V57 V83 -6.394314135553584e-20

R57_84 V57 V84 2598.886007755901
L57_84 V57 V84 -6.409070627157953e-11
C57_84 V57 V84 1.169081442909935e-20

R57_85 V57 V85 2967.227185107471
L57_85 V57 V85 9.018153501759289e-12
C57_85 V57 V85 1.4325864076081683e-19

R57_86 V57 V86 1299.6329462812566
L57_86 V57 V86 1.0353701994041283e-11
C57_86 V57 V86 5.8295440972391454e-21

R57_87 V57 V87 3597.0652599313553
L57_87 V57 V87 6.415289010575516e-12
C57_87 V57 V87 1.3266349093198444e-19

R57_88 V57 V88 2895.96637064016
L57_88 V57 V88 3.6050737307137556e-12
C57_88 V57 V88 1.9774587761372829e-19

R57_89 V57 V89 994.1852806721445
L57_89 V57 V89 1.0294041040850686e-12
C57_89 V57 V89 2.4054856479487064e-19

R57_90 V57 V90 -1727.296658170628
L57_90 V57 V90 3.858487768511241e-12
C57_90 V57 V90 2.078628302015557e-19

R57_91 V57 V91 -1955.9956979418364
L57_91 V57 V91 3.222510676227409e-12
C57_91 V57 V91 5.581123015322953e-20

R57_92 V57 V92 -2143.994349522142
L57_92 V57 V92 1.8224427342284858e-11
C57_92 V57 V92 -4.986283059853629e-20

R57_93 V57 V93 -751.8442010687834
L57_93 V57 V93 -1.831772127522183e-12
C57_93 V57 V93 -3.6758469763407426e-19

R57_94 V57 V94 -2896.041178833691
L57_94 V57 V94 -6.4511059148404026e-12
C57_94 V57 V94 -1.938725297753609e-19

R57_95 V57 V95 -8425.109133677488
L57_95 V57 V95 -2.830668776802104e-12
C57_95 V57 V95 -2.1636008678027118e-19

R57_96 V57 V96 -3475.635067662016
L57_96 V57 V96 -2.5022440722987464e-12
C57_96 V57 V96 -2.474859651368181e-19

R57_97 V57 V97 14361.859498559646
L57_97 V57 V97 -1.3175669940031499e-12
C57_97 V57 V97 -4.729355377541165e-19

R57_98 V57 V98 1247.3634177341658
L57_98 V57 V98 -1.633188004758563e-10
C57_98 V57 V98 -4.137823547850281e-20

R57_99 V57 V99 1960.2756113521502
L57_99 V57 V99 -1.504392530218926e-11
C57_99 V57 V99 7.75406057218276e-20

R57_100 V57 V100 1908.6742598614294
L57_100 V57 V100 -9.324011740187278e-12
C57_100 V57 V100 1.7913662101119003e-19

R57_101 V57 V101 954.735799845703
L57_101 V57 V101 1.4744410538245115e-12
C57_101 V57 V101 4.757199295814947e-19

R57_102 V57 V102 -11703.750967203157
L57_102 V57 V102 -4.7040903878710634e-12
C57_102 V57 V102 5.3906080201675516e-21

R57_103 V57 V103 -16129.976325107418
L57_103 V57 V103 -1.6093142077903635e-11
C57_103 V57 V103 -2.8204873076985066e-20

R57_104 V57 V104 15333.979221540247
L57_104 V57 V104 -1.300196434480809e-11
C57_104 V57 V104 -2.313772223284361e-20

R57_105 V57 V105 -852.3543181547668
L57_105 V57 V105 1.4412757072678246e-12
C57_105 V57 V105 2.6238258487602237e-19

R57_106 V57 V106 -3225.2800321962277
L57_106 V57 V106 3.285388631779938e-12
C57_106 V57 V106 1.659171283504507e-19

R57_107 V57 V107 -14193.673190682804
L57_107 V57 V107 7.050452731228041e-12
C57_107 V57 V107 4.6041172629050745e-20

R57_108 V57 V108 -8599.629304284665
L57_108 V57 V108 2.342342806878483e-12
C57_108 V57 V108 1.2283034463299653e-19

R57_109 V57 V109 -3348.5009843274343
L57_109 V57 V109 -3.287155832066424e-11
C57_109 V57 V109 -1.4725969629890568e-19

R57_110 V57 V110 3491.5366974691956
L57_110 V57 V110 2.7259333983499247e-11
C57_110 V57 V110 -2.7355197075767366e-20

R57_111 V57 V111 7460.047880389316
L57_111 V57 V111 2.531408121192284e-12
C57_111 V57 V111 8.53508050262786e-20

R57_112 V57 V112 14687.30408847157
L57_112 V57 V112 1.180331351542583e-11
C57_112 V57 V112 -9.406023771445725e-20

R57_113 V57 V113 1029.2747504370366
L57_113 V57 V113 -1.9942894339530443e-12
C57_113 V57 V113 -3.9743715594891346e-19

R57_114 V57 V114 -28822.429395921135
L57_114 V57 V114 -2.6028070464325427e-12
C57_114 V57 V114 -2.0218216788847248e-19

R57_115 V57 V115 -5338.278787456464
L57_115 V57 V115 -2.8075087594065724e-12
C57_115 V57 V115 -1.3686713716214354e-19

R57_116 V57 V116 -7458.840767469702
L57_116 V57 V116 -2.0117159938487545e-12
C57_116 V57 V116 -1.8738627772413304e-19

R57_117 V57 V117 -1870.1508958573545
L57_117 V57 V117 -4.324896053415336e-12
C57_117 V57 V117 -8.407547516597718e-20

R57_118 V57 V118 -189679.0169374077
L57_118 V57 V118 3.205307191652967e-12
C57_118 V57 V118 1.9400290738990994e-19

R57_119 V57 V119 7289.410028144378
L57_119 V57 V119 -3.505776173904831e-11
C57_119 V57 V119 1.4238185235415957e-19

R57_120 V57 V120 3653.446418508181
L57_120 V57 V120 7.0715783643343965e-12
C57_120 V57 V120 2.584581474048049e-19

R57_121 V57 V121 -1836.0229264331479
L57_121 V57 V121 1.4377704937046488e-12
C57_121 V57 V121 4.596219851844894e-19

R57_122 V57 V122 -21556.009128089994
L57_122 V57 V122 -1.1963205612436067e-11
C57_122 V57 V122 -2.937896823024458e-20

R57_123 V57 V123 -53626.90560602027
L57_123 V57 V123 -4.746163817628852e-11
C57_123 V57 V123 -1.4753300417451313e-19

R57_124 V57 V124 -5433.802772050309
L57_124 V57 V124 -2.92587127787959e-10
C57_124 V57 V124 -1.8684887843072696e-19

R57_125 V57 V125 1920.5376716945386
L57_125 V57 V125 2.280547095675333e-12
C57_125 V57 V125 2.045868144569478e-19

R57_126 V57 V126 5687.301868291683
L57_126 V57 V126 9.436198952038354e-11
C57_126 V57 V126 6.624449058856274e-20

R57_127 V57 V127 81966.83342511831
L57_127 V57 V127 1.2134429440293002e-11
C57_127 V57 V127 5.2746379875214086e-20

R57_128 V57 V128 124184.50534772853
L57_128 V57 V128 3.211973254867652e-12
C57_128 V57 V128 8.349127926624773e-20

R57_129 V57 V129 -4361.064119044305
L57_129 V57 V129 -4.409807805730072e-12
C57_129 V57 V129 -3.5264365652996755e-19

R57_130 V57 V130 -22413.613877724878
L57_130 V57 V130 -4.6744430688809946e-11
C57_130 V57 V130 -3.00019022823999e-20

R57_131 V57 V131 11575.483911457006
L57_131 V57 V131 1.1408359335052651e-11
C57_131 V57 V131 4.27687314285244e-20

R57_132 V57 V132 6728.390658649992
L57_132 V57 V132 -5.941500436957134e-12
C57_132 V57 V132 2.398224031407232e-21

R57_133 V57 V133 -7947.533336039982
L57_133 V57 V133 -7.942873187543668e-12
C57_133 V57 V133 -8.996907310187058e-20

R57_134 V57 V134 -4535.868516108731
L57_134 V57 V134 -3.4404137515332096e-12
C57_134 V57 V134 -3.9462474759350085e-20

R57_135 V57 V135 -4504.879227731997
L57_135 V57 V135 -7.02784020392074e-12
C57_135 V57 V135 -8.976326623769782e-20

R57_136 V57 V136 -3087.6639642783452
L57_136 V57 V136 -3.5450536355462574e-12
C57_136 V57 V136 -2.4016185242428156e-19

R57_137 V57 V137 55376.471584595354
L57_137 V57 V137 -1.3786563053799276e-12
C57_137 V57 V137 -1.0430379456068986e-19

R57_138 V57 V138 4934.605125744976
L57_138 V57 V138 7.743717737494588e-12
C57_138 V57 V138 2.055629721727602e-20

R57_139 V57 V139 6896.724691589207
L57_139 V57 V139 1.0856829750571229e-11
C57_139 V57 V139 1.4289530521783658e-19

R57_140 V57 V140 2911.287891056128
L57_140 V57 V140 -1.659707826313874e-11
C57_140 V57 V140 1.6050798753419953e-19

R57_141 V57 V141 -11061.226352827638
L57_141 V57 V141 2.4000525016931716e-12
C57_141 V57 V141 2.6863229539819563e-19

R57_142 V57 V142 4002.389070845576
L57_142 V57 V142 2.9307026985718807e-12
C57_142 V57 V142 5.80052174257833e-20

R57_143 V57 V143 5192.8513676004095
L57_143 V57 V143 -7.564614214403629e-12
C57_143 V57 V143 -1.395390302313343e-19

R57_144 V57 V144 20480.6853550699
L57_144 V57 V144 3.0805036915505316e-12
C57_144 V57 V144 1.102194238911776e-19

R57_145 V57 V145 -46499.48846387008
L57_145 V57 V145 7.874877666716803e-13
C57_145 V57 V145 1.417761567308273e-19

R57_146 V57 V146 -3946.0199147434096
L57_146 V57 V146 -2.2296115152356348e-11
C57_146 V57 V146 -5.341203705233418e-20

R57_147 V57 V147 -3549.494350131371
L57_147 V57 V147 3.6544109087943525e-12
C57_147 V57 V147 7.406277390589038e-20

R57_148 V57 V148 -23081.456766854586
L57_148 V57 V148 5.227674692724603e-12
C57_148 V57 V148 -2.647675923886437e-20

R57_149 V57 V149 2443.2401724855895
L57_149 V57 V149 -5.0813224973982934e-12
C57_149 V57 V149 6.431841209305732e-20

R57_150 V57 V150 -4932.675874023562
L57_150 V57 V150 -6.160692410606053e-11
C57_150 V57 V150 -2.3916591138225962e-20

R57_151 V57 V151 -373191.44451522134
L57_151 V57 V151 3.0031405788454544e-12
C57_151 V57 V151 1.1073671238838646e-19

R57_152 V57 V152 -10774.572013933517
L57_152 V57 V152 -7.848132155400575e-12
C57_152 V57 V152 -5.064857747388105e-20

R57_153 V57 V153 -1782.3393605549163
L57_153 V57 V153 -8.900717514643419e-13
C57_153 V57 V153 -3.3589618492327335e-19

R57_154 V57 V154 -120070.05830965615
L57_154 V57 V154 -1.869768285226834e-12
C57_154 V57 V154 -2.5157645614225208e-20

R57_155 V57 V155 -4051.81842152078
L57_155 V57 V155 -4.2837636362230985e-12
C57_155 V57 V155 1.184952102687179e-19

R57_156 V57 V156 6798.510126137068
L57_156 V57 V156 -3.136110510714043e-12
C57_156 V57 V156 -1.84549579288454e-20

R57_157 V57 V157 -1701.2918514767605
L57_157 V57 V157 -1.9647787164618e-12
C57_157 V57 V157 -3.549046577787454e-19

R57_158 V57 V158 3064.3206642645023
L57_158 V57 V158 3.1193597984880884e-12
C57_158 V57 V158 -8.221858871667078e-21

R57_159 V57 V159 3069.3410565267723
L57_159 V57 V159 -2.441425624778763e-12
C57_159 V57 V159 -2.717424456812836e-19

R57_160 V57 V160 -76309.05082278787
L57_160 V57 V160 -4.694769497432096e-12
C57_160 V57 V160 -7.217785651202241e-20

R57_161 V57 V161 1713.8796405661346
L57_161 V57 V161 1.190273439681088e-12
C57_161 V57 V161 4.118952942350553e-19

R57_162 V57 V162 9130.569580078047
L57_162 V57 V162 3.0148300020312636e-12
C57_162 V57 V162 -1.1923803965413166e-19

R57_163 V57 V163 3898.1630283248705
L57_163 V57 V163 -6.431787929678939e-12
C57_163 V57 V163 -1.3469169326454452e-19

R57_164 V57 V164 2316.7132088480043
L57_164 V57 V164 3.5489115269272494e-12
C57_164 V57 V164 4.0224288927062206e-20

R57_165 V57 V165 -6133.120885945671
L57_165 V57 V165 7.216793505563539e-13
C57_165 V57 V165 3.249060644276121e-19

R57_166 V57 V166 -3261.0384082374308
L57_166 V57 V166 8.362337579682057e-12
C57_166 V57 V166 1.471508951521407e-19

R57_167 V57 V167 35185.13158518942
L57_167 V57 V167 2.1116797926449047e-12
C57_167 V57 V167 2.1201332766490278e-19

R57_168 V57 V168 -9325.268003993451
L57_168 V57 V168 2.059687424898738e-12
C57_168 V57 V168 2.968174923377459e-19

R57_169 V57 V169 -1631.5817425309478
L57_169 V57 V169 -7.436379567232161e-13
C57_169 V57 V169 -5.035006004593708e-19

R57_170 V57 V170 3781.6171068527196
L57_170 V57 V170 1.1813953920721073e-11
C57_170 V57 V170 1.1658912859838154e-19

R57_171 V57 V171 -3118.598444014491
L57_171 V57 V171 2.2211696431533543e-12
C57_171 V57 V171 1.8691290409450412e-19

R57_172 V57 V172 -7974.457545227779
L57_172 V57 V172 -1.495552900761822e-11
C57_172 V57 V172 -3.7028520182510016e-20

R57_173 V57 V173 3587.7826787350045
L57_173 V57 V173 -1.898862401323703e-12
C57_173 V57 V173 -1.7602726541304953e-19

R57_174 V57 V174 -8859.809747197234
L57_174 V57 V174 -1.2338256621050077e-12
C57_174 V57 V174 -4.2294038909518235e-19

R57_175 V57 V175 466692.24599697505
L57_175 V57 V175 -1.2555176534857839e-12
C57_175 V57 V175 -2.5771559244758412e-19

R57_176 V57 V176 -31438.41243582454
L57_176 V57 V176 -1.0982913770465922e-12
C57_176 V57 V176 -2.9281650875560983e-19

R57_177 V57 V177 -28953.13821121996
L57_177 V57 V177 1.3140883670956503e-12
C57_177 V57 V177 2.4556174644637206e-19

R57_178 V57 V178 -12098.973058098192
L57_178 V57 V178 1.4367841759533926e-11
C57_178 V57 V178 5.807374860709285e-21

R57_179 V57 V179 6951.741913253364
L57_179 V57 V179 -1.694760154231802e-11
C57_179 V57 V179 -1.0176470495058062e-19

R57_180 V57 V180 7737.6515294105775
L57_180 V57 V180 4.514862655678978e-12
C57_180 V57 V180 -1.1122620563620963e-20

R57_181 V57 V181 2023.7477196414509
L57_181 V57 V181 4.221847846419737e-12
C57_181 V57 V181 4.2196050335025565e-19

R57_182 V57 V182 -40384.78457315545
L57_182 V57 V182 1.966673295008237e-12
C57_182 V57 V182 1.4218076862184257e-19

R57_183 V57 V183 6978.94374618119
L57_183 V57 V183 3.365563651193809e-11
C57_183 V57 V183 -6.120992461094252e-21

R57_184 V57 V184 11508.421240550188
L57_184 V57 V184 3.055710216725555e-12
C57_184 V57 V184 1.216852830859309e-19

R57_185 V57 V185 -3934.823055312652
L57_185 V57 V185 2.2364695497149957e-10
C57_185 V57 V185 -4.1346315578644015e-19

R57_186 V57 V186 68862.25339628675
L57_186 V57 V186 1.6721511560007876e-12
C57_186 V57 V186 2.3597869815323054e-19

R57_187 V57 V187 -4480.237483141868
L57_187 V57 V187 2.355172665511669e-12
C57_187 V57 V187 1.9188506844951132e-19

R57_188 V57 V188 -2418.123304533633
L57_188 V57 V188 2.020475006605091e-12
C57_188 V57 V188 2.0785262852560113e-19

R57_189 V57 V189 -2251.154122423003
L57_189 V57 V189 -1.1542506136931784e-12
C57_189 V57 V189 -5.955973270208031e-20

R57_190 V57 V190 -266896.29882736236
L57_190 V57 V190 -2.6610973420473387e-12
C57_190 V57 V190 -1.4226379873966571e-19

R57_191 V57 V191 -4046.9503855689472
L57_191 V57 V191 6.60662702085277e-12
C57_191 V57 V191 1.215709021255627e-20

R57_192 V57 V192 -13974.591314864261
L57_192 V57 V192 -2.0685776690581407e-12
C57_192 V57 V192 -2.627453218644256e-19

R57_193 V57 V193 2435.4977932265406
L57_193 V57 V193 -9.43722264913772e-11
C57_193 V57 V193 -1.3165551285961569e-19

R57_194 V57 V194 -5252.461317122723
L57_194 V57 V194 -9.011678626903572e-13
C57_194 V57 V194 -3.906590263085928e-19

R57_195 V57 V195 6055.858593398743
L57_195 V57 V195 -2.1146301890915306e-12
C57_195 V57 V195 -1.2620168604678195e-19

R57_196 V57 V196 6482.113082025446
L57_196 V57 V196 -1.556306826018318e-12
C57_196 V57 V196 -7.894941304241161e-20

R57_197 V57 V197 6623.018327231788
L57_197 V57 V197 2.128967684785873e-12
C57_197 V57 V197 2.9346209203653574e-19

R57_198 V57 V198 9290.289182496037
L57_198 V57 V198 1.8978465193390167e-12
C57_198 V57 V198 5.381959128000521e-20

R57_199 V57 V199 3105.2917389253
L57_199 V57 V199 1.1721221661814797e-11
C57_199 V57 V199 -1.8520269694231146e-19

R57_200 V57 V200 4931.819786199399
L57_200 V57 V200 1.523640437568635e-12
C57_200 V57 V200 2.1149014809792e-19

R58_58 V58 0 418.468253457903
L58_58 V58 0 7.611479077351212e-12
C58_58 V58 0 1.1492304592016499e-18

R58_59 V58 V59 -22212.045124501466
L58_59 V58 V59 -1.0795747889754154e-11
C58_59 V58 V59 -8.202100091888818e-20

R58_60 V58 V60 -19621.942646006817
L58_60 V58 V60 -5.726758330826634e-12
C58_60 V58 V60 -7.935863599762928e-20

R58_61 V58 V61 -6463.455655328409
L58_61 V58 V61 5.1872036723115685e-12
C58_61 V58 V61 1.3224023509491433e-19

R58_62 V58 V62 3647.0876995253416
L58_62 V58 V62 -5.181715283817967e-12
C58_62 V58 V62 -1.3969320084748693e-19

R58_63 V58 V63 -17194.05552124639
L58_63 V58 V63 1.0851110811663253e-11
C58_63 V58 V63 1.0378707368737589e-19

R58_64 V58 V64 -6469.892120182633
L58_64 V58 V64 -4.7755253183333776e-11
C58_64 V58 V64 4.981376607402021e-20

R58_65 V58 V65 9237.450446527544
L58_65 V58 V65 4.267066134296363e-12
C58_65 V58 V65 1.7066328928441944e-20

R58_66 V58 V66 15394.36728546425
L58_66 V58 V66 1.3450609400093472e-12
C58_66 V58 V66 4.647111591751418e-19

R58_67 V58 V67 27916.750700817192
L58_67 V58 V67 4.627801561488798e-12
C58_67 V58 V67 8.450349559754836e-20

R58_68 V58 V68 -18793.132300188423
L58_68 V58 V68 5.883252672472161e-12
C58_68 V58 V68 6.533397404903597e-20

R58_69 V58 V69 2907.7008938018025
L58_69 V58 V69 1.207823510262173e-11
C58_69 V58 V69 2.883402066943001e-20

R58_70 V58 V70 -1904.63267484101
L58_70 V58 V70 -5.6865099104884435e-12
C58_70 V58 V70 -1.5944358075064377e-19

R58_71 V58 V71 -4741.998813484232
L58_71 V58 V71 -5.111307918447871e-12
C58_71 V58 V71 -8.381823738791594e-20

R58_72 V58 V72 -3571.4318831758073
L58_72 V58 V72 -1.0259227974154379e-11
C58_72 V58 V72 -7.5816647535096e-21

R58_73 V58 V73 -5671.906159566072
L58_73 V58 V73 -4.316340801114283e-12
C58_73 V58 V73 -1.7495783624851794e-19

R58_74 V58 V74 7777.21164991306
L58_74 V58 V74 -5.369312425734548e-12
C58_74 V58 V74 -1.0219708934217007e-19

R58_75 V58 V75 -20127.86906437627
L58_75 V58 V75 -7.408717643981724e-12
C58_75 V58 V75 -7.63248543378184e-20

R58_76 V58 V76 3312.1818463717755
L58_76 V58 V76 -5.364283908702772e-11
C58_76 V58 V76 2.937225290142931e-21

R58_77 V58 V77 -6556.907865819856
L58_77 V58 V77 -1.4622151461005047e-11
C58_77 V58 V77 1.6792733831346696e-21

R58_78 V58 V78 1335.4604444522552
L58_78 V58 V78 -3.6852988668246543e-11
C58_78 V58 V78 -4.1340788310718436e-20

R58_79 V58 V79 2132.1361607658087
L58_79 V58 V79 6.89895019368125e-12
C58_79 V58 V79 5.3919110491809865e-20

R58_80 V58 V80 2548.2033729343443
L58_80 V58 V80 -1.8501589518546346e-11
C58_80 V58 V80 -4.051512918076845e-20

R58_81 V58 V81 1823.1059041381432
L58_81 V58 V81 3.1223995396639528e-12
C58_81 V58 V81 1.0498897457425292e-19

R58_82 V58 V82 -1849.1952644287812
L58_82 V58 V82 -3.293168817715104e-11
C58_82 V58 V82 -2.76334973387867e-20

R58_83 V58 V83 -3581.560485745654
L58_83 V58 V83 2.6987915217613758e-11
C58_83 V58 V83 3.595991621659933e-20

R58_84 V58 V84 -2915.406753679255
L58_84 V58 V84 -2.209697251161647e-09
C58_84 V58 V84 4.9169538573000013e-20

R58_85 V58 V85 -20011.70426028025
L58_85 V58 V85 -3.927663713163485e-12
C58_85 V58 V85 -1.6413615269197421e-19

R58_86 V58 V86 -704.1090753696362
L58_86 V58 V86 -1.479475030257702e-11
C58_86 V58 V86 1.9470660898361486e-19

R58_87 V58 V87 -2518.6145733810204
L58_87 V58 V87 -2.105775765887698e-11
C58_87 V58 V87 7.948901727756413e-21

R58_88 V58 V88 -2039.3987138574046
L58_88 V58 V88 2.449006930771644e-11
C58_88 V58 V88 6.510686836207112e-20

R58_89 V58 V89 52361.53009298976
L58_89 V58 V89 1.991058057489873e-12
C58_89 V58 V89 2.0045805669527798e-19

R58_90 V58 V90 663.1060557145748
L58_90 V58 V90 6.298093361556616e-12
C58_90 V58 V90 -6.558547212696317e-20

R58_91 V58 V91 3286.6501045477808
L58_91 V58 V91 -1.0954061613606863e-11
C58_91 V58 V91 -1.1424572862740035e-19

R58_92 V58 V92 2607.2063993942606
L58_92 V58 V92 -5.5254841120246276e-12
C58_92 V58 V92 -9.607537643701078e-20

R58_93 V58 V93 10286.212297013273
L58_93 V58 V93 -2.174363289874931e-11
C58_93 V58 V93 -2.065804571172718e-20

R58_94 V58 V94 4024.136138303215
L58_94 V58 V94 7.073439937208338e-11
C58_94 V58 V94 -1.2887393043746954e-19

R58_95 V58 V95 2634.375115314073
L58_95 V58 V95 1.7717471049120097e-11
C58_95 V58 V95 -8.638531750908437e-21

R58_96 V58 V96 1477.6246534096508
L58_96 V58 V96 6.667659481221485e-12
C58_96 V58 V96 -2.7335668870087877e-20

R58_97 V58 V97 2359.1795551983378
L58_97 V58 V97 -3.352875751147943e-12
C58_97 V58 V97 -3.0847515782240507e-19

R58_98 V58 V98 -957.3854991792889
L58_98 V58 V98 -7.268189243708223e-12
C58_98 V58 V98 -3.697570405800379e-20

R58_99 V58 V99 -2520.798888228153
L58_99 V58 V99 8.169452198907066e-12
C58_99 V58 V99 1.3224105367365955e-19

R58_100 V58 V100 -1400.8825775863493
L58_100 V58 V100 -9.873259636960225e-12
C58_100 V58 V100 1.3443066952205227e-19

R58_101 V58 V101 5637.902773628793
L58_101 V58 V101 4.448641784618071e-12
C58_101 V58 V101 1.371099158843162e-19

R58_102 V58 V102 1929.3289301216755
L58_102 V58 V102 6.247513961139207e-12
C58_102 V58 V102 1.2364108401268413e-19

R58_103 V58 V103 -1973.9432616625495
L58_103 V58 V103 -4.909899071437378e-12
C58_103 V58 V103 -3.1122027429337314e-20

R58_104 V58 V104 -1562.8860100466215
L58_104 V58 V104 -3.936012507483501e-12
C58_104 V58 V104 -5.272053561177105e-20

R58_105 V58 V105 -2542.7647269429635
L58_105 V58 V105 3.39845351083475e-12
C58_105 V58 V105 1.6596119260381532e-19

R58_106 V58 V106 -772.9273212195284
L58_106 V58 V106 -1.3913317438538148e-11
C58_106 V58 V106 1.3164619258114948e-19

R58_107 V58 V107 2261.2530602758334
L58_107 V58 V107 1.54156361452486e-11
C58_107 V58 V107 -9.834814968712086e-20

R58_108 V58 V108 1452.7855394502749
L58_108 V58 V108 2.6792067499986e-12
C58_108 V58 V108 1.1012379834898959e-20

R58_109 V58 V109 14569.29801630849
L58_109 V58 V109 6.746189123012364e-11
C58_109 V58 V109 -1.3907286025289456e-19

R58_110 V58 V110 730.3291816507423
L58_110 V58 V110 -3.0159644682806283e-12
C58_110 V58 V110 -3.2568882991854433e-19

R58_111 V58 V111 -6776.070040724115
L58_111 V58 V111 2.4452688479258867e-11
C58_111 V58 V111 2.5074310897117245e-20

R58_112 V58 V112 -6353.5665932553375
L58_112 V58 V112 -8.632203750111412e-12
C58_112 V58 V112 -5.562495200802465e-20

R58_113 V58 V113 888.1462347768055
L58_113 V58 V113 -9.574549123746744e-12
C58_113 V58 V113 -1.6470783838761299e-19

R58_114 V58 V114 1036.5718390176096
L58_114 V58 V114 4.677018831912088e-12
C58_114 V58 V114 1.1298562903353017e-19

R58_115 V58 V115 8428.895575723627
L58_115 V58 V115 1.0753555342629354e-11
C58_115 V58 V115 8.526029255249672e-20

R58_116 V58 V116 -43382.15789585116
L58_116 V58 V116 -2.5986811433217418e-11
C58_116 V58 V116 1.914307654998754e-20

R58_117 V58 V117 4182.186273379088
L58_117 V58 V117 3.430340858376617e-11
C58_117 V58 V117 4.390370617317702e-20

R58_118 V58 V118 -313.2837771302824
L58_118 V58 V118 5.917199235038086e-12
C58_118 V58 V118 1.971262450885122e-19

R58_119 V58 V119 -1775.3927620901638
L58_119 V58 V119 1.5831300133456492e-11
C58_119 V58 V119 5.866956521098461e-20

R58_120 V58 V120 -1875.6786054410045
L58_120 V58 V120 4.35016652336796e-12
C58_120 V58 V120 1.3921899467227827e-19

R58_121 V58 V121 -1044.3179325514852
L58_121 V58 V121 5.8427901158345085e-12
C58_121 V58 V121 1.441554030814122e-19

R58_122 V58 V122 1088.4252818215261
L58_122 V58 V122 -5.34534680987904e-12
C58_122 V58 V122 -2.2967285960745575e-19

R58_123 V58 V123 -7975.113561254959
L58_123 V58 V123 -2.9931772536368724e-12
C58_123 V58 V123 -1.3447645335150862e-19

R58_124 V58 V124 59884.815286304685
L58_124 V58 V124 -2.0759371036806913e-12
C58_124 V58 V124 -2.334599543097827e-19

R58_125 V58 V125 -2086.039509138146
L58_125 V58 V125 6.383400799581139e-12
C58_125 V58 V125 5.050359661582103e-20

R58_126 V58 V126 379.9147439058455
L58_126 V58 V126 -3.9165806669850654e-11
C58_126 V58 V126 1.3032323591158983e-19

R58_127 V58 V127 766.6375927683825
L58_127 V58 V127 8.820772878781583e-12
C58_127 V58 V127 4.351548375741301e-21

R58_128 V58 V128 783.0900890431961
L58_128 V58 V128 4.5449187518877494e-12
C58_128 V58 V128 4.5612977815540674e-20

R58_129 V58 V129 537.9249079442077
L58_129 V58 V129 -1.3413940444091364e-11
C58_129 V58 V129 -2.6596684859946524e-19

R58_130 V58 V130 -617.1804457564878
L58_130 V58 V130 -2.1648109884517973e-11
C58_130 V58 V130 3.767503759513493e-20

R58_131 V58 V131 -683.7776093069995
L58_131 V58 V131 9.23851658511429e-12
C58_131 V58 V131 6.518568817766423e-20

R58_132 V58 V132 -515.9749268309941
L58_132 V58 V132 5.131841067399556e-12
C58_132 V58 V132 1.1242585892173185e-19

R58_133 V58 V133 13212.563436997409
L58_133 V58 V133 3.024074682932132e-11
C58_133 V58 V133 1.6213299679622985e-19

R58_134 V58 V134 -674.0127421652907
L58_134 V58 V134 -1.8046508104587035e-11
C58_134 V58 V134 -1.4803894170079132e-19

R58_135 V58 V135 -1567.7677632664231
L58_135 V58 V135 -5.213232027817485e-12
C58_135 V58 V135 -1.4411940364498362e-20

R58_136 V58 V136 -871.0939405807532
L58_136 V58 V136 -2.7775510714911098e-12
C58_136 V58 V136 -1.8915941646743651e-19

R58_137 V58 V137 -611.9014758494992
L58_137 V58 V137 -7.485357342027071e-12
C58_137 V58 V137 4.7006000344574136e-20

R58_138 V58 V138 490.5079289519149
L58_138 V58 V138 9.756956468783228e-12
C58_138 V58 V138 1.532338201446218e-19

R58_139 V58 V139 509.50346835478655
L58_139 V58 V139 3.369781379386647e-12
C58_139 V58 V139 7.032011930092234e-20

R58_140 V58 V140 379.98042200829514
L58_140 V58 V140 3.591149033590769e-12
C58_140 V58 V140 2.0031239392881548e-19

R58_141 V58 V141 -1083.9244241318956
L58_141 V58 V141 -5.66182150324925e-12
C58_141 V58 V141 -1.6589763269782296e-19

R58_142 V58 V142 792.7311242162023
L58_142 V58 V142 -2.8517086161365984e-12
C58_142 V58 V142 -5.944400027847101e-20

R58_143 V58 V143 -1162.7799459603366
L58_143 V58 V143 -7.705886931184931e-12
C58_143 V58 V143 -1.1790526136897738e-19

R58_144 V58 V144 -13000.698442450865
L58_144 V58 V144 8.046503762147613e-12
C58_144 V58 V144 -3.543675830393886e-20

R58_145 V58 V145 404.6496221177552
L58_145 V58 V145 4.543488873037779e-12
C58_145 V58 V145 -3.0056119421830747e-20

R58_146 V58 V146 -560.7443152539146
L58_146 V58 V146 1.6013941352327687e-11
C58_146 V58 V146 3.048774213465244e-20

R58_147 V58 V147 3502.324864253772
L58_147 V58 V147 -3.912163868992463e-12
C58_147 V58 V147 1.9683710531354175e-20

R58_148 V58 V148 -685.6525633769322
L58_148 V58 V148 -1.980300822495482e-12
C58_148 V58 V148 -7.614742744404772e-20

R58_149 V58 V149 14000.71821138807
L58_149 V58 V149 1.8822499490026233e-12
C58_149 V58 V149 2.9318043732222923e-19

R58_150 V58 V150 -320.3201783009399
L58_150 V58 V150 1.7122602596138275e-12
C58_150 V58 V150 -1.6016617199893677e-19

R58_151 V58 V151 -1882.7919827936864
L58_151 V58 V151 -2.6191286125605002e-11
C58_151 V58 V151 4.820797966301118e-20

R58_152 V58 V152 919.1199106839088
L58_152 V58 V152 -1.5319988090045403e-11
C58_152 V58 V152 6.849183603933577e-21

R58_153 V58 V153 -809.2933208001076
L58_153 V58 V153 -5.6163399701821805e-12
C58_153 V58 V153 -6.036080125088862e-20

R58_154 V58 V154 635.9315278120255
L58_154 V58 V154 -1.3848260087409925e-11
C58_154 V58 V154 9.584783592427913e-20

R58_155 V58 V155 474.6401260548217
L58_155 V58 V155 3.1998861707668647e-12
C58_155 V58 V155 9.668846957025016e-20

R58_156 V58 V156 -871.6180832335892
L58_156 V58 V156 6.8680233870001805e-12
C58_156 V58 V156 4.819749221360501e-20

R58_157 V58 V157 -993.0289033492271
L58_157 V58 V157 -1.7375144837386342e-12
C58_157 V58 V157 -3.3541998968785234e-19

R58_158 V58 V158 1326.1822332001082
L58_158 V58 V158 -9.183265437389223e-13
C58_158 V58 V158 -3.975647667065351e-20

R58_159 V58 V159 -478.4668553637014
L58_159 V58 V159 8.96164026399617e-12
C58_159 V58 V159 -6.524100149752819e-20

R58_160 V58 V160 -4544.2755515301815
L58_160 V58 V160 3.4633754073586956e-12
C58_160 V58 V160 1.0072471706073898e-20

R58_161 V58 V161 497.40733377113656
L58_161 V58 V161 5.302376884314198e-12
C58_161 V58 V161 4.124982821937723e-20

R58_162 V58 V162 2021.9044089039312
L58_162 V58 V162 3.558661138944366e-12
C58_162 V58 V162 6.410176320844937e-20

R58_163 V58 V163 1309.3561852800603
L58_163 V58 V163 -3.206582579315902e-12
C58_163 V58 V163 -7.489320444105638e-20

R58_164 V58 V164 1895.7363396680998
L58_164 V58 V164 -3.1144871618178454e-12
C58_164 V58 V164 3.0847533952746827e-20

R58_165 V58 V165 4938.2302999190815
L58_165 V58 V165 1.597506761681157e-12
C58_165 V58 V165 2.5009782425324665e-19

R58_166 V58 V166 -419.92168532719995
L58_166 V58 V166 8.138479126360806e-13
C58_166 V58 V166 -5.958976664510066e-20

R58_167 V58 V167 -1150369.226918837
L58_167 V58 V167 -2.8680762064421713e-12
C58_167 V58 V167 9.190903819209382e-21

R58_168 V58 V168 711.6727356685667
L58_168 V58 V168 -5.801759175532682e-12
C58_168 V58 V168 -1.1473636995853314e-20

R58_169 V58 V169 -406.1069930135016
L58_169 V58 V169 -4.0387463150567396e-12
C58_169 V58 V169 -1.3869989902304377e-19

R58_170 V58 V170 12174.662272151761
L58_170 V58 V170 -1.7288802248440905e-12
C58_170 V58 V170 1.2027270732814232e-19

R58_171 V58 V171 -13576.366328068649
L58_171 V58 V171 1.8059991048714034e-12
C58_171 V58 V171 1.5776514663960686e-19

R58_172 V58 V172 -1148.1997016203263
L58_172 V58 V172 4.627310637909589e-12
C58_172 V58 V172 8.044232456251734e-20

R58_173 V58 V173 660.2061481500233
L58_173 V58 V173 -1.9228972554085607e-12
C58_173 V58 V173 -1.0564574247824579e-19

R58_174 V58 V174 483.70426656972893
L58_174 V58 V174 -1.1218091007682387e-12
C58_174 V58 V174 -1.3445477675571022e-19

R58_175 V58 V175 -1366.045885265354
L58_175 V58 V175 1.528600042624103e-11
C58_175 V58 V175 -3.00170058649813e-21

R58_176 V58 V176 -2004.7742150642339
L58_176 V58 V176 6.774306193743013e-12
C58_176 V58 V176 1.7553803668030122e-20

R58_177 V58 V177 1599.3387333388937
L58_177 V58 V177 6.735171424485176e-12
C58_177 V58 V177 4.9981549191329586e-20

R58_178 V58 V178 -2897.248581759685
L58_178 V58 V178 2.8983175532280492e-12
C58_178 V58 V178 -6.567114352697878e-20

R58_179 V58 V179 1141.9845521258449
L58_179 V58 V179 -1.928086361400973e-12
C58_179 V58 V179 -1.7066306879742794e-19

R58_180 V58 V180 1627.2453106196465
L58_180 V58 V180 -1.958924938229192e-12
C58_180 V58 V180 -1.5682507170627598e-19

R58_181 V58 V181 -901.3039551207783
L58_181 V58 V181 1.9412936179585154e-12
C58_181 V58 V181 1.0648031132528993e-19

R58_182 V58 V182 -577.2320252872331
L58_182 V58 V182 2.2419064694095993e-12
C58_182 V58 V182 8.428367089653364e-20

R58_183 V58 V183 -2617.0886619673893
L58_183 V58 V183 -6.515204884143929e-12
C58_183 V58 V183 -3.124913757233964e-20

R58_184 V58 V184 -43740.96416627353
L58_184 V58 V184 -2.7170286653721696e-11
C58_184 V58 V184 5.425272741005101e-20

R58_185 V58 V185 22186.83675031486
L58_185 V58 V185 -3.0503313239432472e-12
C58_185 V58 V185 -8.580456802676322e-20

R58_186 V58 V186 7139.764352583438
L58_186 V58 V186 2.176519780372745e-12
C58_186 V58 V186 5.626758755475204e-20

R58_187 V58 V187 3967.4444562422973
L58_187 V58 V187 1.897779873980714e-12
C58_187 V58 V187 1.8308296254619287e-19

R58_188 V58 V188 1100.4213407090685
L58_188 V58 V188 1.3901914107161947e-12
C58_188 V58 V188 1.4010832901867211e-19

R58_189 V58 V189 -8957.682951984792
L58_189 V58 V189 -1.6178968190442267e-12
C58_189 V58 V189 6.977973033606722e-21

R58_190 V58 V190 1752.5092012505795
L58_190 V58 V190 -1.616769071858067e-12
C58_190 V58 V190 -1.2362852278540777e-19

R58_191 V58 V191 4813.535444546245
L58_191 V58 V191 -3.0311013026690003e-11
C58_191 V58 V191 3.609419595070967e-20

R58_192 V58 V192 -6869.5222520000125
L58_192 V58 V192 -2.0934118228436596e-12
C58_192 V58 V192 -6.313420612244785e-20

R58_193 V58 V193 1393.6724716676395
L58_193 V58 V193 2.301479208569823e-12
C58_193 V58 V193 -4.4612634380043766e-20

R58_194 V58 V194 -1165.7086795299517
L58_194 V58 V194 -2.167787425722744e-12
C58_194 V58 V194 -9.133708908747808e-20

R58_195 V58 V195 -1700.5771688688753
L58_195 V58 V195 -2.2502564080971305e-12
C58_195 V58 V195 -1.8401944925266197e-19

R58_196 V58 V196 -1045.619368199673
L58_196 V58 V196 -3.0029928766610642e-12
C58_196 V58 V196 -9.5550367929868e-20

R58_197 V58 V197 -16535.509041123412
L58_197 V58 V197 9.448678015009253e-12
C58_197 V58 V197 -9.718996590458823e-21

R58_198 V58 V198 -934.9714466078257
L58_198 V58 V198 1.2022605153494038e-12
C58_198 V58 V198 -4.9715192167677485e-21

R58_199 V58 V199 -2105.8952066519673
L58_199 V58 V199 3.54921471470027e-12
C58_199 V58 V199 -1.0859724943044037e-19

R58_200 V58 V200 791.9775471374651
L58_200 V58 V200 2.4162446106464834e-12
C58_200 V58 V200 4.9561774712814905e-20

R59_59 V59 0 -470.09632861649237
L59_59 V59 0 -6.52967889216548e-13
C59_59 V59 0 1.6202627594460116e-18

R59_60 V59 V60 -2087.703517919517
L59_60 V59 V60 -1.989160401867622e-12
C59_60 V59 V60 -2.9651482911163896e-19

R59_61 V59 V61 -11356.749182152804
L59_61 V59 V61 3.5550169249966644e-12
C59_61 V59 V61 1.9543291308490245e-19

R59_62 V59 V62 -5836.362604739407
L59_62 V59 V62 -6.544554628821522e-12
C59_62 V59 V62 -1.3823094756449098e-19

R59_63 V59 V63 4851.7035863040255
L59_63 V59 V63 1.6518063984017024e-12
C59_63 V59 V63 6.088034073243202e-19

R59_64 V59 V64 8486.583818971905
L59_64 V59 V64 5.0759110874356444e-12
C59_64 V59 V64 2.175599600353488e-19

R59_65 V59 V65 5432.902738758737
L59_65 V59 V65 7.351012149152801e-12
C59_65 V59 V65 -7.321780985999995e-20

R59_66 V59 V66 23633.587018272774
L59_66 V59 V66 -1.1007332474480794e-11
C59_66 V59 V66 -7.581236954978355e-20

R59_67 V59 V67 1880.6503181641874
L59_67 V59 V67 9.913117040727893e-13
C59_67 V59 V67 6.322550362218692e-19

R59_68 V59 V68 3508.385989387932
L59_68 V59 V68 5.859495325388984e-12
C59_68 V59 V68 8.220388558800543e-20

R59_69 V59 V69 2537.704302745194
L59_69 V59 V69 1.2511762328874476e-11
C59_69 V59 V69 4.653971850115648e-21

R59_70 V59 V70 187766.53650366951
L59_70 V59 V70 3.728787065877224e-12
C59_70 V59 V70 2.4233150581816395e-19

R59_71 V59 V71 -6444.899905852146
L59_71 V59 V71 -9.076493847972695e-13
C59_71 V59 V71 -9.042603579609663e-19

R59_72 V59 V72 -40708.537410170255
L59_72 V59 V72 -1.2005946712908714e-11
C59_72 V59 V72 -6.189276042099692e-20

R59_73 V59 V73 -176525.44945917197
L59_73 V59 V73 5.211868171492745e-11
C59_73 V59 V73 -4.7216577753189725e-20

R59_74 V59 V74 -8598.856094695253
L59_74 V59 V74 -1.2213147549841183e-11
C59_74 V59 V74 -1.563639434293856e-19

R59_75 V59 V75 -2087.718439396615
L59_75 V59 V75 4.565121775379996e-12
C59_75 V59 V75 2.192575472099656e-19

R59_76 V59 V76 -3228.010717893194
L59_76 V59 V76 1.6888915338241455e-11
C59_76 V59 V76 1.03513597911805e-19

R59_77 V59 V77 -2173.3361094821526
L59_77 V59 V77 -3.339122321072325e-12
C59_77 V59 V77 -1.5858776586597293e-19

R59_78 V59 V78 4186.978856488224
L59_78 V59 V78 5.072065916152959e-10
C59_78 V59 V78 4.486896028829655e-20

R59_79 V59 V79 2147.5099067722003
L59_79 V59 V79 4.23286515908208e-12
C59_79 V59 V79 1.7735437009549233e-19

R59_80 V59 V80 5745.404607568379
L59_80 V59 V80 -7.111119967874653e-12
C59_80 V59 V80 -1.0953669178012722e-19

R59_81 V59 V81 1152.067062289713
L59_81 V59 V81 2.826181593088985e-12
C59_81 V59 V81 7.43852194266065e-20

R59_82 V59 V82 -6388.212907905513
L59_82 V59 V82 -5.904413925314966e-12
C59_82 V59 V82 -1.4948225495277417e-19

R59_83 V59 V83 -4641.94666733436
L59_83 V59 V83 -3.492164107156408e-12
C59_83 V59 V83 -2.891547174294274e-19

R59_84 V59 V84 -17623.413406471624
L59_84 V59 V84 -5.357397056391862e-12
C59_84 V59 V84 -5.669193548512895e-20

R59_85 V59 V85 -16197.298803312806
L59_85 V59 V85 -6.508180817009287e-12
C59_85 V59 V85 -9.932872970190852e-20

R59_86 V59 V86 -2157.1546059728853
L59_86 V59 V86 -6.040507767239037e-12
C59_86 V59 V86 -1.105695259100272e-19

R59_87 V59 V87 -1444.722950148371
L59_87 V59 V87 1.8301695650038832e-12
C59_87 V59 V87 4.524811557154827e-19

R59_88 V59 V88 -3644.452079590154
L59_88 V59 V88 3.671529231159767e-12
C59_88 V59 V88 2.460708826845744e-19

R59_89 V59 V89 149606.56890126836
L59_89 V59 V89 1.7098221932738937e-12
C59_89 V59 V89 2.686125644370837e-19

R59_90 V59 V90 2531.647307527334
L59_90 V59 V90 1.6248121519429793e-12
C59_90 V59 V90 4.600350971766363e-19

R59_91 V59 V91 613.2142575045723
L59_91 V59 V91 -1.2209112612525749e-12
C59_91 V59 V91 -5.835807996664705e-19

R59_92 V59 V92 2694.006016499238
L59_92 V59 V92 -3.6286037221853776e-12
C59_92 V59 V92 -2.1007487325853724e-19

R59_93 V59 V93 3474.5022273718623
L59_93 V59 V93 -3.352944017099682e-11
C59_93 V59 V93 -3.8119593091222776e-20

R59_94 V59 V94 4941.45044652138
L59_94 V59 V94 -4.521589412472375e-12
C59_94 V59 V94 -2.222993775341564e-19

R59_95 V59 V95 -4959.794534913892
L59_95 V59 V95 -1.8104728481243567e-12
C59_95 V59 V95 -2.890785446562513e-19

R59_96 V59 V96 152538.32639489823
L59_96 V59 V96 -1.9429713542661136e-11
C59_96 V59 V96 -1.5015842697489628e-19

R59_97 V59 V97 -16419.733439158408
L59_97 V59 V97 -1.6636067056565501e-12
C59_97 V59 V97 -5.425486028636638e-19

R59_98 V59 V98 -2370.2965542683687
L59_98 V59 V98 -2.3756891108999195e-12
C59_98 V59 V98 -2.957818008726458e-19

R59_99 V59 V99 -657.3921445516193
L59_99 V59 V99 7.251625109694046e-13
C59_99 V59 V99 8.445639644609003e-19

R59_100 V59 V100 -2061.494912517072
L59_100 V59 V100 2.1175927389372473e-11
C59_100 V59 V100 3.5420898997872244e-19

R59_101 V59 V101 2188.0122056607975
L59_101 V59 V101 2.781610430227993e-12
C59_101 V59 V101 3.1103922390703747e-19

R59_102 V59 V102 -3869.383534629559
L59_102 V59 V102 3.916645537510829e-12
C59_102 V59 V102 2.4221553045190226e-19

R59_103 V59 V103 2005.622563871566
L59_103 V59 V103 -4.696970001654988e-12
C59_103 V59 V103 -2.62324202874873e-19

R59_104 V59 V104 -6638.936683303896
L59_104 V59 V104 -4.1481075502278474e-12
C59_104 V59 V104 -1.482179719082043e-19

R59_105 V59 V105 3562.6824149219683
L59_105 V59 V105 1.5951122114856164e-12
C59_105 V59 V105 2.4796862730715367e-19

R59_106 V59 V106 4552.639621306265
L59_106 V59 V106 2.8886116575004936e-12
C59_106 V59 V106 2.7215729856468214e-19

R59_107 V59 V107 947.6712029189631
L59_107 V59 V107 -1.0173281334835391e-12
C59_107 V59 V107 -3.8261368738045194e-19

R59_108 V59 V108 2156.3322258454755
L59_108 V59 V108 2.886015125273087e-12
C59_108 V59 V108 2.46567423909032e-20

R59_109 V59 V109 -1308.0049512193236
L59_109 V59 V109 -1.0407255329143878e-11
C59_109 V59 V109 -3.147484430033287e-19

R59_110 V59 V110 12054.590247938017
L59_110 V59 V110 -3.9797744568852635e-12
C59_110 V59 V110 -2.3034418212120415e-19

R59_111 V59 V111 -4818.224909997964
L59_111 V59 V111 2.0730749891740312e-12
C59_111 V59 V111 1.5625523967761088e-19

R59_112 V59 V112 28127.403634386774
L59_112 V59 V112 -8.848064572850394e-12
C59_112 V59 V112 -7.438488739179359e-20

R59_113 V59 V113 824.6128546986557
L59_113 V59 V113 -1.8400551962650564e-12
C59_113 V59 V113 -2.0486728624502296e-19

R59_114 V59 V114 -3803.7945578450167
L59_114 V59 V114 -3.3325600272386566e-12
C59_114 V59 V114 -2.5752596083311287e-19

R59_115 V59 V115 -688.7182355557175
L59_115 V59 V115 1.817909580053185e-12
C59_115 V59 V115 2.221025125050531e-19

R59_116 V59 V116 -1283.7330739215463
L59_116 V59 V116 -1.7755680420570224e-11
C59_116 V59 V116 -2.5534158728944803e-20

R59_117 V59 V117 2318.922062994998
L59_117 V59 V117 3.41036782737259e-11
C59_117 V59 V117 1.3428708446443215e-19

R59_118 V59 V118 54761.122528401895
L59_118 V59 V118 2.5054831685572814e-12
C59_118 V59 V118 3.9035935663080312e-19

R59_119 V59 V119 784.5522522391158
L59_119 V59 V119 -1.1314962188618812e-12
C59_119 V59 V119 1.188431679335998e-19

R59_120 V59 V120 1584.2263533173436
L59_120 V59 V120 4.712071886311212e-12
C59_120 V59 V120 2.9947200750780616e-19

R59_121 V59 V121 -909.0441636250114
L59_121 V59 V121 1.405447296024182e-12
C59_121 V59 V121 1.353905961631386e-19

R59_122 V59 V122 -34061.900966421286
L59_122 V59 V122 -1.1092182703109624e-11
C59_122 V59 V122 -8.626558825917452e-20

R59_123 V59 V123 -15454.626254452012
L59_123 V59 V123 4.80094940839927e-12
C59_123 V59 V123 -4.5833249582674335e-19

R59_124 V59 V124 24603.178309207604
L59_124 V59 V124 -2.5447641620600976e-12
C59_124 V59 V124 -4.134786501934145e-19

R59_125 V59 V125 2028.964757000891
L59_125 V59 V125 4.911777237612325e-12
C59_125 V59 V125 7.404733788764234e-20

R59_126 V59 V126 2288.3743235017114
L59_126 V59 V126 -4.660862588073007e-12
C59_126 V59 V126 -1.4946809986279835e-19

R59_127 V59 V127 -8955.714970673047
L59_127 V59 V127 2.096440400257377e-12
C59_127 V59 V127 1.0294055545397084e-19

R59_128 V59 V128 -2665.448143692549
L59_128 V59 V128 4.1784506718008235e-12
C59_128 V59 V128 4.760987615685721e-21

R59_129 V59 V129 1427.2684115898835
L59_129 V59 V129 -1.694485063289094e-12
C59_129 V59 V129 -3.780923353402696e-19

R59_130 V59 V130 -2787.3643585852533
L59_130 V59 V130 4.314154861375124e-12
C59_130 V59 V130 1.7524497139715928e-19

R59_131 V59 V131 -5131.22581877752
L59_131 V59 V131 -1.8418559327149896e-12
C59_131 V59 V131 2.467946308858885e-19

R59_132 V59 V132 4065.680262449577
L59_132 V59 V132 -5.1117260415739026e-11
C59_132 V59 V132 3.4571372447956446e-19

R59_133 V59 V133 -6030.999011653053
L59_133 V59 V133 -1.8059520837228754e-09
C59_133 V59 V133 1.7501525997446774e-19

R59_134 V59 V134 -5017.843337639038
L59_134 V59 V134 -2.8694024561803317e-12
C59_134 V59 V134 -5.373552584636916e-20

R59_135 V59 V135 -809.0954704006625
L59_135 V59 V135 1.7844544517838292e-12
C59_135 V59 V135 -3.4691712478228236e-19

R59_136 V59 V136 -3470.5009908350303
L59_136 V59 V136 -2.6935447992896766e-12
C59_136 V59 V136 -3.31512773684259e-19

R59_137 V59 V137 -1822.5500202543267
L59_137 V59 V137 2.5957400593161193e-12
C59_137 V59 V137 1.2984142573880877e-19

R59_138 V59 V138 3946.0091359698395
L59_138 V59 V138 4.63164421358532e-12
C59_138 V59 V138 -9.053268610386608e-20

R59_139 V59 V139 503.9303419525827
L59_139 V59 V139 -4.555050815448135e-12
C59_139 V59 V139 4.606453918102277e-19

R59_140 V59 V140 1769.9636867070353
L59_140 V59 V140 2.22863269924046e-12
C59_140 V59 V140 2.8490963308099726e-19

R59_141 V59 V141 -2562.324863942445
L59_141 V59 V141 -5.435144246240059e-12
C59_141 V59 V141 -2.8363213507977854e-19

R59_142 V59 V142 5847.846340296967
L59_142 V59 V142 2.9936606064380395e-12
C59_142 V59 V142 5.134868530621313e-20

R59_143 V59 V143 1646.8771016257595
L59_143 V59 V143 -8.523492629506501e-13
C59_143 V59 V143 -2.0471939076218683e-19

R59_144 V59 V144 3952.961757997929
L59_144 V59 V144 -1.4287701561608605e-11
C59_144 V59 V144 -2.009393825457876e-20

R59_145 V59 V145 699.9998605883624
L59_145 V59 V145 -3.9693733970272975e-12
C59_145 V59 V145 -1.0273532503960619e-19

R59_146 V59 V146 -1000069.2670575518
L59_146 V59 V146 -1.6228382759819793e-12
C59_146 V59 V146 7.04302665054911e-20

R59_147 V59 V147 -343.9541392544135
L59_147 V59 V147 8.203109618452622e-13
C59_147 V59 V147 -3.162940021456135e-19

R59_148 V59 V148 -2224.514119647387
L59_148 V59 V148 -1.5444271374734483e-12
C59_148 V59 V148 -1.924755421924557e-19

R59_149 V59 V149 -4638.6295980786435
L59_149 V59 V149 9.404202480707237e-13
C59_149 V59 V149 5.859104432282206e-19

R59_150 V59 V150 -2042.3717975530055
L59_150 V59 V150 6.502365733591047e-11
C59_150 V59 V150 -2.803120419183885e-19

R59_151 V59 V151 609.0766160664626
L59_151 V59 V151 9.036029580692102e-13
C59_151 V59 V151 2.3713266346031296e-19

R59_152 V59 V152 6178.42340331061
L59_152 V59 V152 5.580523423098135e-12
C59_152 V59 V152 1.4488316495158586e-20

R59_153 V59 V153 -1647.2726221226912
L59_153 V59 V153 -4.8982917218393274e-12
C59_153 V59 V153 -1.0153471607200192e-19

R59_154 V59 V154 -4772.31681532505
L59_154 V59 V154 4.578537061841577e-12
C59_154 V59 V154 1.0610407009324901e-19

R59_155 V59 V155 -324.16116972852853
L59_155 V59 V155 -1.5619738985668659e-12
C59_155 V59 V155 2.7341511456003967e-19

R59_156 V59 V156 171898.53107521552
L59_156 V59 V156 5.625212770120189e-12
C59_156 V59 V156 1.4443977036837553e-19

R59_157 V59 V157 -1528.500049065378
L59_157 V59 V157 -1.1598742324657517e-12
C59_157 V59 V157 -6.551472890665188e-19

R59_158 V59 V158 2072.4980411153724
L59_158 V59 V158 5.701497719800996e-12
C59_158 V59 V158 6.3516813334046e-20

R59_159 V59 V159 539.565810100134
L59_159 V59 V159 -6.747984105763345e-13
C59_159 V59 V159 -2.3682698778477674e-19

R59_160 V59 V160 -2860.8816323130022
L59_160 V59 V160 1.9145857048804014e-11
C59_160 V59 V160 -7.524370154412478e-21

R59_161 V59 V161 902.3300838156267
L59_161 V59 V161 2.0810078162232395e-12
C59_161 V59 V161 2.0615828552876702e-19

R59_162 V59 V162 2367.551772209705
L59_162 V59 V162 4.643554667762668e-12
C59_162 V59 V162 7.422053246943692e-20

R59_163 V59 V163 916.1907556837733
L59_163 V59 V163 1.2286453489014389e-12
C59_163 V59 V163 -6.838622199761053e-20

R59_164 V59 V164 905.7335398882204
L59_164 V59 V164 -1.5972783759539325e-11
C59_164 V59 V164 6.084548900536e-20

R59_165 V59 V165 858.8457529694246
L59_165 V59 V165 1.1122560228220273e-12
C59_165 V59 V165 2.803138691590218e-19

R59_166 V59 V166 -1230.2168717529962
L59_166 V59 V166 1.5166340769701504e-11
C59_166 V59 V166 -1.0116906595063467e-19

R59_167 V59 V167 -1388.3706827797341
L59_167 V59 V167 2.884554275579328e-12
C59_167 V59 V167 9.98727232413213e-20

R59_168 V59 V168 -2682.9100098499407
L59_168 V59 V168 6.229594449403131e-12
C59_168 V59 V168 2.4397052474729468e-20

R59_169 V59 V169 -1151.0172001178448
L59_169 V59 V169 -1.4953156292578842e-12
C59_169 V59 V169 -3.278460908706212e-19

R59_170 V59 V170 1401.5536156628455
L59_170 V59 V170 -1.522466122928491e-11
C59_170 V59 V170 1.5100192754475104e-19

R59_171 V59 V171 -595.7008792950663
L59_171 V59 V171 6.3911612688578e-12
C59_171 V59 V171 1.1543772243816131e-19

R59_172 V59 V172 -3326.427720300256
L59_172 V59 V172 -4.4708031174027783e-11
C59_172 V59 V172 5.358541956112008e-20

R59_173 V59 V173 -14687.472254563474
L59_173 V59 V173 -3.2878968702743406e-12
C59_173 V59 V173 -3.202605921613122e-20

R59_174 V59 V174 -2181.076083810575
L59_174 V59 V174 -4.5304563522195594e-12
C59_174 V59 V174 -2.1887468026599386e-19

R59_175 V59 V175 627.3546203727457
L59_175 V59 V175 -7.72535785347472e-12
C59_175 V59 V175 1.621380526779178e-19

R59_176 V59 V176 -3456.3095340917903
L59_176 V59 V176 -6.221525778390888e-12
C59_176 V59 V176 4.925597349039065e-20

R59_177 V59 V177 1024.3773918469788
L59_177 V59 V177 2.473087859847468e-12
C59_177 V59 V177 8.34669513036765e-20

R59_178 V59 V178 24266.940814276164
L59_178 V59 V178 -1.894859414205052e-11
C59_178 V59 V178 -8.685707627960825e-20

R59_179 V59 V179 -1950.6488322254233
L59_179 V59 V179 -1.8294283736035362e-12
C59_179 V59 V179 -3.6853994385112484e-19

R59_180 V59 V180 2280.4432176718697
L59_180 V59 V180 -4.433247245513304e-12
C59_180 V59 V180 -2.48004382375407e-19

R59_181 V59 V181 -1373.0375539089869
L59_181 V59 V181 1.190517938991967e-11
C59_181 V59 V181 7.13647825662951e-20

R59_182 V59 V182 -2243.143825555217
L59_182 V59 V182 2.2907713777423896e-12
C59_182 V59 V182 2.0542700180929938e-19

R59_183 V59 V183 4498.650433014529
L59_183 V59 V183 -1.9786209010472436e-11
C59_183 V59 V183 -6.55409683265185e-20

R59_184 V59 V184 3185.3714708219204
L59_184 V59 V184 -7.539098321848488e-12
C59_184 V59 V184 4.036929791684496e-20

R59_185 V59 V185 -9389.382248962376
L59_185 V59 V185 -4.758024541059579e-12
C59_185 V59 V185 -6.528843435917087e-20

R59_186 V59 V186 -127367.52958033426
L59_186 V59 V186 3.8428296941370035e-12
C59_186 V59 V186 2.672641178872464e-20

R59_187 V59 V187 14942.335954646485
L59_187 V59 V187 1.3819002333770335e-12
C59_187 V59 V187 3.7986592722080456e-19

R59_188 V59 V188 -1269.053200892033
L59_188 V59 V188 1.1551280965812993e-12
C59_188 V59 V188 2.513814787053889e-19

R59_189 V59 V189 49107.7741461846
L59_189 V59 V189 -3.889976962243477e-12
C59_189 V59 V189 -9.845076645582707e-21

R59_190 V59 V190 4614.477518405565
L59_190 V59 V190 -5.079892426946709e-12
C59_190 V59 V190 -1.8504383417296721e-19

R59_191 V59 V191 -30934.580101576485
L59_191 V59 V191 1.4992879830511933e-11
C59_191 V59 V191 -3.329938417782602e-20

R59_192 V59 V192 15605.166599896696
L59_192 V59 V192 -3.4157293598989294e-12
C59_192 V59 V192 -1.2406977611903484e-19

R59_193 V59 V193 3010.9671571629956
L59_193 V59 V193 5.7481702295731406e-12
C59_193 V59 V193 -1.0631942298688622e-19

R59_194 V59 V194 -2146.0710856969417
L59_194 V59 V194 -1.574050718510062e-12
C59_194 V59 V194 -2.48209565328472e-19

R59_195 V59 V195 16585.53476937439
L59_195 V59 V195 -1.8675113831173406e-12
C59_195 V59 V195 -6.403236713266517e-20

R59_196 V59 V196 1245.8938416330118
L59_196 V59 V196 -1.3673257211283997e-12
C59_196 V59 V196 -9.938111828020819e-20

R59_197 V59 V197 7875.226978792416
L59_197 V59 V197 -3.429141429192209e-11
C59_197 V59 V197 6.696451344661143e-20

R59_198 V59 V198 -27863.598576619483
L59_198 V59 V198 3.2350303758834087e-12
C59_198 V59 V198 2.4638553971740067e-20

R59_199 V59 V199 -2033.9178174086858
L59_199 V59 V199 4.338316455772392e-12
C59_199 V59 V199 -1.5388257367096714e-19

R59_200 V59 V200 -8021.787367487257
L59_200 V59 V200 2.1663345331007788e-12
C59_200 V59 V200 1.1503357661281105e-19

R60_60 V60 0 -232.9142117941365
L60_60 V60 0 -4.3875046900563056e-13
C60_60 V60 0 1.860884482806582e-18

R60_61 V60 V61 -11108.077642236834
L60_61 V60 V61 2.584896707858512e-12
C60_61 V60 V61 2.3473703382936785e-19

R60_62 V60 V62 -4666.986808032072
L60_62 V60 V62 -4.403136346687249e-12
C60_62 V60 V62 -1.823829423559629e-19

R60_63 V60 V63 14393.781278128872
L60_63 V60 V63 4.273572108530454e-12
C60_63 V60 V63 2.5517230068867473e-19

R60_64 V60 V64 2086.555403223862
L60_64 V60 V64 1.5313628028427054e-12
C60_64 V60 V64 6.316780506365438e-19

R60_65 V60 V65 3913.1567129335895
L60_65 V60 V65 6.341939869124823e-12
C60_65 V60 V65 -9.248760834363772e-20

R60_66 V60 V66 23263.85089859107
L60_66 V60 V66 -9.24521003319474e-12
C60_66 V60 V66 -9.261830725835063e-20

R60_67 V60 V67 5155.721388988175
L60_67 V60 V67 5.87881629463186e-12
C60_67 V60 V67 1.0068359476750744e-19

R60_68 V60 V68 1297.6748714509972
L60_68 V60 V68 9.184187729736023e-13
C60_68 V60 V68 6.598734482662057e-19

R60_69 V60 V69 2104.930033493496
L60_69 V60 V69 4.3958547070760305e-12
C60_69 V60 V69 1.9070537778179275e-20

R60_70 V60 V70 -37056.26511436585
L60_70 V60 V70 2.2818454300552374e-12
C60_70 V60 V70 3.3382678176127737e-19

R60_71 V60 V71 -26315.381412397026
L60_71 V60 V71 -6.3172038316744674e-12
C60_71 V60 V71 -1.7689408122345572e-19

R60_72 V60 V72 -3852.644947811713
L60_72 V60 V72 -9.051048758549322e-13
C60_72 V60 V72 -9.344377753883464e-19

R60_73 V60 V73 69202.41835427257
L60_73 V60 V73 -2.272554136155925e-11
C60_73 V60 V73 -7.567488053748406e-20

R60_74 V60 V74 -6006.35286807606
L60_74 V60 V74 -7.485984533699655e-12
C60_74 V60 V74 -1.8737996433395325e-19

R60_75 V60 V75 -5309.025398836079
L60_75 V60 V75 -4.152925623522819e-12
C60_75 V60 V75 -1.1319686621949786e-19

R60_76 V60 V76 -1110.2114188399516
L60_76 V60 V76 1.862276559780608e-12
C60_76 V60 V76 4.540533094405004e-19

R60_77 V60 V77 -1679.990858009211
L60_77 V60 V77 -2.1631585572016216e-12
C60_77 V60 V77 -1.8988967331798838e-19

R60_78 V60 V78 2368.1298085171097
L60_78 V60 V78 -2.5298845202217753e-11
C60_78 V60 V78 -4.933829628597516e-21

R60_79 V60 V79 12482.005542451217
L60_79 V60 V79 1.0870038328304254e-11
C60_79 V60 V79 5.183449815221804e-20

R60_80 V60 V80 1059.9408323157418
L60_80 V60 V80 -4.3564304866814795e-12
C60_80 V60 V80 -1.5690085341236126e-20

R60_81 V60 V81 797.9954021758164
L60_81 V60 V81 2.0931399032186143e-12
C60_81 V60 V81 1.060613840072711e-19

R60_82 V60 V82 -3574.455138054927
L60_82 V60 V82 -5.067000685060892e-12
C60_82 V60 V82 -1.421411515571306e-19

R60_83 V60 V83 -11916.707808286275
L60_83 V60 V83 -6.164795748693989e-12
C60_83 V60 V83 -5.614386373867652e-22

R60_84 V60 V84 -6622.339086276041
L60_84 V60 V84 -2.9524863733466287e-12
C60_84 V60 V84 -3.265398111429645e-19

R60_85 V60 V85 -18822.968194651115
L60_85 V60 V85 -5.7576147513501495e-12
C60_85 V60 V85 -1.0697095703224146e-19

R60_86 V60 V86 -1683.2607678504448
L60_86 V60 V86 -5.5041756332375415e-12
C60_86 V60 V86 -7.727755494830939e-20

R60_87 V60 V87 -2716.6478823457946
L60_87 V60 V87 6.372308893382605e-12
C60_87 V60 V87 1.6998063916887327e-19

R60_88 V60 V88 -818.9226455454036
L60_88 V60 V88 1.3056802535864783e-12
C60_88 V60 V88 5.823616218757179e-19

R60_89 V60 V89 -10712.810344774562
L60_89 V60 V89 1.196453150536101e-12
C60_89 V60 V89 3.5033465908983046e-19

R60_90 V60 V90 2127.0641849338026
L60_90 V60 V90 1.3705836778703312e-12
C60_90 V60 V90 4.9652272309974345e-19

R60_91 V60 V91 1311.9311914093967
L60_91 V60 V91 -3.1408234593670594e-12
C60_91 V60 V91 -3.1345602838840254e-19

R60_92 V60 V92 458.5452110800963
L60_92 V60 V92 -1.2062494062716978e-12
C60_92 V60 V92 -5.3978879232573465e-19

R60_93 V60 V93 2991.733142004116
L60_93 V60 V93 -8.292676625556616e-12
C60_93 V60 V93 -7.291210018188086e-20

R60_94 V60 V94 8964.045336907326
L60_94 V60 V94 -3.0437835677534372e-12
C60_94 V60 V94 -2.6552247681700227e-19

R60_95 V60 V95 -45117.61596925286
L60_95 V60 V95 -6.766570176488742e-12
C60_95 V60 V95 -1.3877187490540819e-19

R60_96 V60 V96 -4943.043412272029
L60_96 V60 V96 -2.0753170482479903e-12
C60_96 V60 V96 -2.946599072004673e-19

R60_97 V60 V97 52170.20655669185
L60_97 V60 V97 -1.2283390002331513e-12
C60_97 V60 V97 -6.0305909834992e-19

R60_98 V60 V98 -3206.821913534316
L60_98 V60 V98 -2.080144714413532e-12
C60_98 V60 V98 -3.053420523809348e-19

R60_99 V60 V99 -1147.25925037289
L60_99 V60 V99 2.868829505468458e-12
C60_99 V60 V99 4.693885090235171e-19

R60_100 V60 V100 -454.69213970752844
L60_100 V60 V100 1.065206847924873e-12
C60_100 V60 V100 7.283840482008696e-19

R60_101 V60 V101 1656.231673998345
L60_101 V60 V101 2.1093348091176563e-12
C60_101 V60 V101 3.7343589453392693e-19

R60_102 V60 V102 -3912.06539075207
L60_102 V60 V102 3.1442363941127765e-12
C60_102 V60 V102 2.886967040148341e-19

R60_103 V60 V103 69145.05441752907
L60_103 V60 V103 -4.014165341121694e-12
C60_103 V60 V103 -1.0728131226204343e-19

R60_104 V60 V104 2100.907075897392
L60_104 V60 V104 -4.379574256549993e-12
C60_104 V60 V104 -2.438999586185351e-19

R60_105 V60 V105 3927.850186369548
L60_105 V60 V105 1.2168026036689611e-12
C60_105 V60 V105 2.954953313803922e-19

R60_106 V60 V106 -9679.873598026761
L60_106 V60 V106 3.1094564054754545e-12
C60_106 V60 V106 2.3224034520299594e-19

R60_107 V60 V107 1573.6979237594192
L60_107 V60 V107 -4.258470789118841e-12
C60_107 V60 V107 -2.617958949945021e-19

R60_108 V60 V108 546.0674199990091
L60_108 V60 V108 -2.2871777090440695e-12
C60_108 V60 V108 -8.41626095472653e-20

R60_109 V60 V109 -1037.361635504414
L60_109 V60 V109 -5.634341686716741e-12
C60_109 V60 V109 -3.428723915558904e-19

R60_110 V60 V110 2622.757090926629
L60_110 V60 V110 -4.669758983085436e-12
C60_110 V60 V110 -2.368139163986122e-19

R60_111 V60 V111 14147.333438544954
L60_111 V60 V111 5.782147575679562e-12
C60_111 V60 V111 7.363649994971966e-20

R60_112 V60 V112 -1262.2136286365726
L60_112 V60 V112 6.2562368106510516e-12
C60_112 V60 V112 -4.7124185824151883e-20

R60_113 V60 V113 560.582246906917
L60_113 V60 V113 -1.622354990318005e-12
C60_113 V60 V113 -2.5996111491258757e-19

R60_114 V60 V114 -5940.2880091120305
L60_114 V60 V114 -3.912714667164533e-12
C60_114 V60 V114 -2.4259808767316715e-19

R60_115 V60 V115 -963.7264874864287
L60_115 V60 V115 3.168347452305579e-12
C60_115 V60 V115 1.5560590955019105e-19

R60_116 V60 V116 -449.32900403714086
L60_116 V60 V116 2.145154760252228e-12
C60_116 V60 V116 6.379772240879471e-20

R60_117 V60 V117 2680.4604685152763
L60_117 V60 V117 9.135174229353265e-12
C60_117 V60 V117 1.4871881099695467e-19

R60_118 V60 V118 -2149.4963344105627
L60_118 V60 V118 1.881593588782835e-12
C60_118 V60 V118 4.1738958382291506e-19

R60_119 V60 V119 1658.3244161414302
L60_119 V60 V119 1.6619462650415288e-11
C60_119 V60 V119 1.3249418300149882e-19

R60_120 V60 V120 327.89227836379814
L60_120 V60 V120 -1.4601561547843599e-12
C60_120 V60 V120 3.0024928447401835e-19

R60_121 V60 V121 -762.0313748152056
L60_121 V60 V121 1.244673669328235e-12
C60_121 V60 V121 2.079197747579793e-19

R60_122 V60 V122 3711.702051166571
L60_122 V60 V122 -3.987448858032679e-12
C60_122 V60 V122 -1.454729951335367e-19

R60_123 V60 V123 3564.5530087431766
L60_123 V60 V123 -2.2551246185820503e-12
C60_123 V60 V123 -2.8676771727512656e-19

R60_124 V60 V124 -839.3945782695552
L60_124 V60 V124 1.134228910737127e-11
C60_124 V60 V124 -5.697024821877458e-19

R60_125 V60 V125 1142.1074878419413
L60_125 V60 V125 5.065848521694244e-12
C60_125 V60 V125 7.361349874163584e-20

R60_126 V60 V126 1067.2193880520426
L60_126 V60 V126 -4.011918907904589e-12
C60_126 V60 V126 -1.3874628272754066e-19

R60_127 V60 V127 -5898.721627568227
L60_127 V60 V127 4.453269546941395e-11
C60_127 V60 V127 -4.3148120937906634e-20

R60_128 V60 V128 -1144.8220054607714
L60_128 V60 V128 1.8304490538185686e-12
C60_128 V60 V128 6.641530717187778e-20

R60_129 V60 V129 1654.7486832336758
L60_129 V60 V129 -1.5758357676243559e-12
C60_129 V60 V129 -4.69465465178177e-19

R60_130 V60 V130 -1221.7565022408762
L60_130 V60 V130 2.342001323284208e-12
C60_130 V60 V130 2.1012761376998039e-19

R60_131 V60 V131 14076.24065986143
L60_131 V60 V131 4.6860355106012836e-12
C60_131 V60 V131 2.0651851613245481e-19

R60_132 V60 V132 1109.4928831704412
L60_132 V60 V132 -1.6967198240322905e-12
C60_132 V60 V132 4.507820380680482e-19

R60_133 V60 V133 -78795.6291455997
L60_133 V60 V133 1.8990963597225023e-11
C60_133 V60 V133 2.2893962803118147e-19

R60_134 V60 V134 27855.927074069717
L60_134 V60 V134 -2.2928101664126696e-12
C60_134 V60 V134 -1.2269919101141813e-19

R60_135 V60 V135 -2460.5991350548475
L60_135 V60 V135 -1.0181874883889233e-11
C60_135 V60 V135 -1.0133120971881954e-19

R60_136 V60 V136 -549.8887953749199
L60_136 V60 V136 1.0048437143411031e-11
C60_136 V60 V136 -5.251906922870052e-19

R60_137 V60 V137 -1230.729994833843
L60_137 V60 V137 2.3444793216990616e-12
C60_137 V60 V137 1.6617609853111533e-19

R60_138 V60 V138 5119.5010716585075
L60_138 V60 V138 3.6376804274306546e-12
C60_138 V60 V138 -4.64367936869993e-20

R60_139 V60 V139 2564.986645972158
L60_139 V60 V139 1.9758770134280273e-12
C60_139 V60 V139 1.7685095560145294e-19

R60_140 V60 V140 329.7434293585412
L60_140 V60 V140 3.459140117149133e-12
C60_140 V60 V140 4.419115148236595e-19

R60_141 V60 V141 -1774.9739691848918
L60_141 V60 V141 -3.13634304718751e-12
C60_141 V60 V141 -3.5066016818359146e-19

R60_142 V60 V142 7625.854419845023
L60_142 V60 V142 2.7136842173783783e-12
C60_142 V60 V142 6.247576832067745e-20

R60_143 V60 V143 2385.8678895570974
L60_143 V60 V143 -1.955910700065803e-12
C60_143 V60 V143 -2.0625088556796647e-19

R60_144 V60 V144 -1681.6261341545303
L60_144 V60 V144 -1.4365157347874558e-12
C60_144 V60 V144 -2.9038055296663824e-20

R60_145 V60 V145 517.3454231263393
L60_145 V60 V145 -6.1646091509174065e-12
C60_145 V60 V145 -1.2309251543415102e-19

R60_146 V60 V146 -12938.828948161736
L60_146 V60 V146 -1.195906240599484e-12
C60_146 V60 V146 6.613744290113103e-20

R60_147 V60 V147 -841.7357943950287
L60_147 V60 V147 -4.586265984807067e-12
C60_147 V60 V147 -1.4551531958225149e-19

R60_148 V60 V148 -1609.1784962888148
L60_148 V60 V148 1.8429149772459177e-12
C60_148 V60 V148 -3.7687339886430424e-19

R60_149 V60 V149 -3639.2707245481442
L60_149 V60 V149 7.342965708704597e-13
C60_149 V60 V149 7.303308510899746e-19

R60_150 V60 V150 -1376.6735801505142
L60_150 V60 V150 4.6623679841942346e-12
C60_150 V60 V150 -3.3944781649611643e-19

R60_151 V60 V151 1795.7033659200824
L60_151 V60 V151 2.8223297276816695e-12
C60_151 V60 V151 1.8070880473885748e-19

R60_152 V60 V152 -951.7421333734017
L60_152 V60 V152 9.792330766167441e-13
C60_152 V60 V152 9.234077489655494e-20

R60_153 V60 V153 -927.823579829312
L60_153 V60 V153 -4.091001240491542e-12
C60_153 V60 V153 -1.1486691482207136e-19

R60_154 V60 V154 -1444.2959640338306
L60_154 V60 V154 5.530619002545297e-12
C60_154 V60 V154 1.6030677050317425e-19

R60_155 V60 V155 -599.0272658353243
L60_155 V60 V155 2.1526335815245966e-12
C60_155 V60 V155 2.148662741238085e-19

R60_156 V60 V156 555.386776993678
L60_156 V60 V156 -1.212598750272443e-12
C60_156 V60 V156 2.733733694472885e-19

R60_157 V60 V157 -2845.263082459415
L60_157 V60 V157 -7.937972694639477e-13
C60_157 V60 V157 -7.910906843602364e-19

R60_158 V60 V158 1062.0336894609704
L60_158 V60 V158 6.6004355110842165e-12
C60_158 V60 V158 6.097970186807249e-20

R60_159 V60 V159 1302.5885091363755
L60_159 V60 V159 -3.0320920924058287e-12
C60_159 V60 V159 -1.116263756005434e-19

R60_160 V60 V160 -3236.5743685039665
L60_160 V60 V160 -6.071671714106257e-13
C60_160 V60 V160 -1.4068662635434907e-19

R60_161 V60 V161 954.7908874213734
L60_161 V60 V161 1.5646143201383395e-12
C60_161 V60 V161 2.2719167424622255e-19

R60_162 V60 V162 1752.459156928259
L60_162 V60 V162 5.495615093358815e-12
C60_162 V60 V162 7.306832188121661e-20

R60_163 V60 V163 1184.8343138240257
L60_163 V60 V163 -2.2185581230373992e-12
C60_163 V60 V163 -1.3242972894670587e-19

R60_164 V60 V164 464.05809669346394
L60_164 V60 V164 8.549832287788239e-13
C60_164 V60 V164 1.2061237477433035e-19

R60_165 V60 V165 552.8847703826813
L60_165 V60 V165 7.846504716585612e-13
C60_165 V60 V165 3.8501608431040395e-19

R60_166 V60 V166 -1033.6725856874984
L60_166 V60 V166 9.490907926146898e-12
C60_166 V60 V166 -1.0575689699137463e-19

R60_167 V60 V167 2640.332211785916
L60_167 V60 V167 8.58421401336231e-12
C60_167 V60 V167 7.952697004538072e-20

R60_168 V60 V168 -428.95555801333353
L60_168 V60 V168 1.5505629999103001e-12
C60_168 V60 V168 1.8778805725754797e-20

R60_169 V60 V169 -754.5909805388453
L60_169 V60 V169 -1.1021280724600383e-12
C60_169 V60 V169 -3.3518686030652565e-19

R60_170 V60 V170 2400.0794025444334
L60_170 V60 V170 2.048460643248105e-11
C60_170 V60 V170 2.199772046478553e-19

R60_171 V60 V171 -861.8363669195811
L60_171 V60 V171 1.3014425703085319e-12
C60_171 V60 V171 2.6069301915892044e-19

R60_172 V60 V172 -1886.0659729851081
L60_172 V60 V172 -2.3837728631593204e-12
C60_172 V60 V172 5.3280912424417716e-20

R60_173 V60 V173 -15126.23106678937
L60_173 V60 V173 -2.111571294262556e-12
C60_173 V60 V173 -1.063177881086554e-19

R60_174 V60 V174 -4783.701976897945
L60_174 V60 V174 -1.858871616558157e-12
C60_174 V60 V174 -2.829669878524613e-19

R60_175 V60 V175 20778.350372729314
L60_175 V60 V175 -2.1645191109077513e-12
C60_175 V60 V175 -1.0021414352578153e-20

R60_176 V60 V176 827.8670856088632
L60_176 V60 V176 8.654734266699287e-12
C60_176 V60 V176 1.912132781107123e-19

R60_177 V60 V177 762.5878918279438
L60_177 V60 V177 1.6464429617181963e-12
C60_177 V60 V177 1.15283434367024e-19

R60_178 V60 V178 5056.258226096861
L60_178 V60 V178 -5.5490294392274995e-11
C60_178 V60 V178 -1.178258991517844e-19

R60_179 V60 V179 21038.712193632306
L60_179 V60 V179 -2.1466249124858454e-12
C60_179 V60 V179 -3.571879149277154e-19

R60_180 V60 V180 1033.7824285983143
L60_180 V60 V180 -1.2955491311333176e-12
C60_180 V60 V180 -3.903295232463506e-19

R60_181 V60 V181 -1005.7749987393746
L60_181 V60 V181 1.007857247689878e-11
C60_181 V60 V181 9.449061828172346e-20

R60_182 V60 V182 -972.0399921673167
L60_182 V60 V182 1.5175534310731385e-12
C60_182 V60 V182 2.2850565894944308e-19

R60_183 V60 V183 1314.1860102335968
L60_183 V60 V183 -2.740307616438184e-12
C60_183 V60 V183 -7.33943905711459e-20

R60_184 V60 V184 -3865.260210906962
L60_184 V60 V184 3.952891108063969e-12
C60_184 V60 V184 5.884747194944224e-20

R60_185 V60 V185 -7405.019172843737
L60_185 V60 V185 -3.5199530037782576e-12
C60_185 V60 V185 -9.11706561754673e-20

R60_186 V60 V186 2675.209818509317
L60_186 V60 V186 2.7430134514606002e-12
C60_186 V60 V186 8.105520287442493e-20

R60_187 V60 V187 9011.294606683836
L60_187 V60 V187 1.381046515489968e-12
C60_187 V60 V187 3.6729515670114607e-19

R60_188 V60 V188 -479.3482847275153
L60_188 V60 V188 7.554075950969457e-13
C60_188 V60 V188 3.135772573766388e-19

R60_189 V60 V189 -10515.650747446838
L60_189 V60 V189 -3.658810760045805e-12
C60_189 V60 V189 3.795944011602958e-20

R60_190 V60 V190 2151.1132170874384
L60_190 V60 V190 -3.5686164140664036e-12
C60_190 V60 V190 -2.1572473947686454e-19

R60_191 V60 V191 -1053.4317494150785
L60_191 V60 V191 1.8118983547069714e-12
C60_191 V60 V191 9.947801170607997e-20

R60_192 V60 V192 899.3362136965717
L60_192 V60 V192 -1.2287745862341504e-12
C60_192 V60 V192 -1.6683291733616972e-19

R60_193 V60 V193 2532.647583896819
L60_193 V60 V193 8.242982442014587e-12
C60_193 V60 V193 -1.6926223573316946e-19

R60_194 V60 V194 -1714.526816918597
L60_194 V60 V194 -1.0677242423104899e-12
C60_194 V60 V194 -2.7791493660332665e-19

R60_195 V60 V195 1516.0121222282542
L60_195 V60 V195 -8.855512267957332e-13
C60_195 V60 V195 -3.7828973499922483e-19

R60_196 V60 V196 1759.1737207849599
L60_196 V60 V196 -1.5109077632192917e-12
C60_196 V60 V196 5.0170567060470186e-20

R60_197 V60 V197 15476.649807011529
L60_197 V60 V197 -3.7152658644480305e-11
C60_197 V60 V197 7.021430958259895e-20

R60_198 V60 V198 -14181.774562262985
L60_198 V60 V198 2.112362189789569e-12
C60_198 V60 V198 2.9966845308077126e-20

R60_199 V60 V199 1243.2609569932456
L60_199 V60 V199 1.1757454463633705e-11
C60_199 V60 V199 -8.567755538749274e-20

R60_200 V60 V200 -792.1292890350676
L60_200 V60 V200 1.31628727305199e-12
C60_200 V60 V200 -1.905906397606945e-20

R61_61 V61 0 -681.4191253625814
L61_61 V61 0 2.811353713095094e-13
C61_61 V61 0 9.268012645393614e-19

R61_62 V61 V62 708359.3056850228
L61_62 V61 V62 -8.126848697177095e-12
C61_62 V61 V62 -1.025533507440884e-19

R61_63 V61 V63 -23963.002542324943
L61_63 V61 V63 -1.495920083869103e-11
C61_63 V61 V63 -1.0904445469589576e-19

R61_64 V61 V64 -7534.696636088361
L61_64 V61 V64 -4.19987606239595e-12
C61_64 V61 V64 -1.908420056045845e-19

R61_65 V61 V65 16244.15016746392
L61_65 V61 V65 -6.626181571797098e-12
C61_65 V61 V65 -1.199340261779642e-19

R61_66 V61 V66 32837.39334590149
L61_66 V61 V66 -7.06720062503367e-12
C61_66 V61 V66 -8.2502361436249e-20

R61_67 V61 V67 14002.197820606392
L61_67 V61 V67 -5.274124639853799e-12
C61_67 V61 V67 -1.2735477132907046e-19

R61_68 V61 V68 -391114.0181109343
L61_68 V61 V68 -2.219336751972494e-12
C61_68 V61 V68 -2.6065614127110457e-19

R61_69 V61 V69 1008.2027344959074
L61_69 V61 V69 2.8102589033655075e-12
C61_69 V61 V69 3.768182658832249e-19

R61_70 V61 V70 -4245.872326817577
L61_70 V61 V70 2.5240582119987173e-11
C61_70 V61 V70 -1.941036659749253e-20

R61_71 V61 V71 -2834.6465737141157
L61_71 V61 V71 -1.6619035174645326e-11
C61_71 V61 V71 3.055637233364154e-20

R61_72 V61 V72 -3025.1365257630264
L61_72 V61 V72 2.0093198035589727e-11
C61_72 V61 V72 1.1087708184186738e-19

R61_73 V61 V73 -1775.8627607665358
L61_73 V61 V73 -6.981579604554083e-12
C61_73 V61 V73 -4.648327265761565e-20

R61_74 V61 V74 44442.83447571144
L61_74 V61 V74 3.649535123021985e-12
C61_74 V61 V74 2.1938415950241096e-19

R61_75 V61 V75 8437.351023508809
L61_75 V61 V75 4.8125762351142345e-12
C61_75 V61 V75 9.356741571461573e-20

R61_76 V61 V76 3409.0107094059344
L61_76 V61 V76 1.82482139167094e-12
C61_76 V61 V76 2.314564758366104e-19

R61_77 V61 V77 -2037.7970627490738
L61_77 V61 V77 3.2753625868327966e-12
C61_77 V61 V77 2.279510413001709e-19

R61_78 V61 V78 2561.610155491437
L61_78 V61 V78 -1.9241486723106478e-11
C61_78 V61 V78 -1.5184520128724058e-20

R61_79 V61 V79 2032.7285145887674
L61_79 V61 V79 3.5570506855016734e-11
C61_79 V61 V79 7.98919428895992e-21

R61_80 V61 V80 2468.9525777879544
L61_80 V61 V80 -4.247068156127121e-12
C61_80 V61 V80 -9.689802257388332e-20

R61_81 V61 V81 668.5440994043493
L61_81 V61 V81 -2.828060266138656e-12
C61_81 V61 V81 -3.107905817064931e-19

R61_82 V61 V82 -4300.758605742686
L61_82 V61 V82 -3.792469268495052e-12
C61_82 V61 V82 -1.6720958451693965e-19

R61_83 V61 V83 -1855.1373862618213
L61_83 V61 V83 -2.1829222250598994e-11
C61_83 V61 V83 7.011249232054038e-21

R61_84 V61 V84 -1879.261612229526
L61_84 V61 V84 -3.3134070751133476e-12
C61_84 V61 V84 -1.5419542179731284e-19

R61_85 V61 V85 -1841.824812805788
L61_85 V61 V85 -1.0805250696761489e-11
C61_85 V61 V85 -1.9162520364226456e-19

R61_86 V61 V86 -812.8079029305671
L61_86 V61 V86 -9.582979148655363e-12
C61_86 V61 V86 -6.144242461204983e-20

R61_87 V61 V87 -3581.633625348864
L61_87 V61 V87 1.1508665849134324e-11
C61_87 V61 V87 1.7040083100221416e-20

R61_88 V61 V88 -3322.581298594696
L61_88 V61 V88 4.336024038542802e-12
C61_88 V61 V88 6.619969633064101e-20

R61_89 V61 V89 -1137.054525399552
L61_89 V61 V89 -9.682414469375464e-12
C61_89 V61 V89 2.1344143169407066e-20

R61_90 V61 V90 910.0486681638167
L61_90 V61 V90 1.851247566978068e-12
C61_90 V61 V90 2.5660796167257247e-19

R61_91 V61 V91 1690.6924222578616
L61_91 V61 V91 -2.485227523451225e-12
C61_91 V61 V91 -2.2297620815704494e-19

R61_92 V61 V92 2345.8564152930862
L61_92 V61 V92 -3.518914647795658e-12
C61_92 V61 V92 -7.30978774659975e-20

R61_93 V61 V93 551.8050493999197
L61_93 V61 V93 3.264699600117118e-12
C61_93 V61 V93 3.071493007032559e-19

R61_94 V61 V94 1666.0675021548097
L61_94 V61 V94 -1.0778075708084835e-11
C61_94 V61 V94 1.0270001682840744e-20

R61_95 V61 V95 8821.045483567013
L61_95 V61 V95 8.768173410971286e-12
C61_95 V61 V95 8.983710589125181e-20

R61_96 V61 V96 2872.077862955256
L61_96 V61 V96 6.043891570319429e-12
C61_96 V61 V96 7.481433861705984e-20

R61_97 V61 V97 -26080.654446160956
L61_97 V61 V97 -6.364185223589605e-12
C61_97 V61 V97 -3.858799230664831e-20

R61_98 V61 V98 -695.3431440772358
L61_98 V61 V98 -2.5898109835457273e-12
C61_98 V61 V98 -2.418539181800816e-19

R61_99 V61 V99 -1847.6748923148941
L61_99 V61 V99 2.0875781547019475e-12
C61_99 V61 V99 2.3779485758218694e-19

R61_100 V61 V100 -1754.9226659314218
L61_100 V61 V100 5.0951935625611195e-12
C61_100 V61 V100 6.583790174851546e-20

R61_101 V61 V101 -713.5241838590216
L61_101 V61 V101 9.876964374342681e-12
C61_101 V61 V101 -5.75972562926269e-20

R61_102 V61 V102 8560.260920917426
L61_102 V61 V102 3.791236791878529e-12
C61_102 V61 V102 1.571198582022823e-19

R61_103 V61 V103 -9566.29542683932
L61_103 V61 V103 -6.890917315386633e-12
C61_103 V61 V103 -4.37589885055865e-20

R61_104 V61 V104 -2903.3738908008295
L61_104 V61 V104 -5.311020317311154e-12
C61_104 V61 V104 -5.831151316608586e-20

R61_105 V61 V105 534.1391963293444
L61_105 V61 V105 -1.8709393691617537e-11
C61_105 V61 V105 -1.5008476351035162e-19

R61_106 V61 V106 2295.4728125670845
L61_106 V61 V106 4.077830155829506e-12
C61_106 V61 V106 8.527272338065258e-20

R61_107 V61 V107 -31769.92558952568
L61_107 V61 V107 -3.649777622263553e-12
C61_107 V61 V107 -2.1593172629585723e-19

R61_108 V61 V108 7894.530995647979
L61_108 V61 V108 -6.317826801236516e-11
C61_108 V61 V108 -9.254707837469125e-20

R61_109 V61 V109 3161.761893694758
L61_109 V61 V109 -2.3767981241452666e-12
C61_109 V61 V109 -1.6944714905723905e-19

R61_110 V61 V110 -3241.937519001176
L61_110 V61 V110 -4.677806125254696e-12
C61_110 V61 V110 -1.356528115720129e-19

R61_111 V61 V111 5308.761208246546
L61_111 V61 V111 -7.477022336361434e-12
C61_111 V61 V111 -2.128360899280899e-20

R61_112 V61 V112 4067.052691953393
L61_112 V61 V112 -7.10833606382555e-12
C61_112 V61 V112 2.013338573559797e-20

R61_113 V61 V113 -737.7661079962979
L61_113 V61 V113 6.910738553795719e-12
C61_113 V61 V113 3.5841390063499016e-19

R61_114 V61 V114 -22641.769311628166
L61_114 V61 V114 -4.122724235166105e-12
C61_114 V61 V114 -6.352650768499389e-20

R61_115 V61 V115 6011.253140643956
L61_115 V61 V115 2.581921096171284e-12
C61_115 V61 V115 2.103349268086838e-19

R61_116 V61 V116 10239.251665266675
L61_116 V61 V116 3.4113317390488448e-12
C61_116 V61 V116 1.6059484196128154e-19

R61_117 V61 V117 851.1425113771417
L61_117 V61 V117 2.000275023177119e-12
C61_117 V61 V117 1.6751533435109257e-19

R61_118 V61 V118 32069.932589290707
L61_118 V61 V118 2.890610904366358e-12
C61_118 V61 V118 1.2433621500796167e-19

R61_119 V61 V119 -2242.799352934814
L61_119 V61 V119 9.678864078907021e-12
C61_119 V61 V119 -4.2727309760023235e-20

R61_120 V61 V120 -1414.781309727233
L61_120 V61 V120 7.155533334897298e-12
C61_120 V61 V120 -1.9466856984085698e-20

R61_121 V61 V121 1876.4479833900548
L61_121 V61 V121 -2.93327194514474e-12
C61_121 V61 V121 -3.3462426987989974e-19

R61_122 V61 V122 -20990.96410561832
L61_122 V61 V122 -1.505303035383087e-11
C61_122 V61 V122 -8.721152706503709e-21

R61_123 V61 V123 6490.875584132621
L61_123 V61 V123 -2.976526643923541e-12
C61_123 V61 V123 -4.2777542020850655e-20

R61_124 V61 V124 2586.235611776974
L61_124 V61 V124 -2.0417987724470954e-12
C61_124 V61 V124 -1.377348451439966e-19

R61_125 V61 V125 -1283.0237881444295
L61_125 V61 V125 -2.8114627677965524e-12
C61_125 V61 V125 -1.5088857996326902e-19

R61_126 V61 V126 -4263.89949642549
L61_126 V61 V126 -2.4700294257781344e-12
C61_126 V61 V126 -1.8474139873672934e-19

R61_127 V61 V127 16206.225376472348
L61_127 V61 V127 -9.823924879028014e-12
C61_127 V61 V127 -7.747755693897228e-20

R61_128 V61 V128 3650.02637462676
L61_128 V61 V128 -2.0172200956869524e-11
C61_128 V61 V128 -7.340099579674732e-20

R61_129 V61 V129 1943.1274948294058
L61_129 V61 V129 7.393496012200289e-12
C61_129 V61 V129 5.432746281738705e-20

R61_130 V61 V130 7914.090718878007
L61_130 V61 V130 2.7215597860719804e-12
C61_130 V61 V130 1.367183240501347e-19

R61_131 V61 V131 -5343.826168246125
L61_131 V61 V131 4.415564072979705e-12
C61_131 V61 V131 8.653842834358212e-20

R61_132 V61 V132 -2053.364080401652
L61_132 V61 V132 2.178800574385084e-12
C61_132 V61 V132 2.288198891128175e-19

R61_133 V61 V133 2721.895961483807
L61_133 V61 V133 5.6732725330607446e-12
C61_133 V61 V133 2.3145466292651533e-19

R61_134 V61 V134 -9047.05137732459
L61_134 V61 V134 -1.171627196591855e-11
C61_134 V61 V134 -3.586584415718064e-20

R61_135 V61 V135 3507.604663833248
L61_135 V61 V135 -1.817933444402825e-11
C61_135 V61 V135 8.02474268615453e-21

R61_136 V61 V136 2737.844856659252
L61_136 V61 V136 -7.9938303598682e-12
C61_136 V61 V136 -2.3509539094760325e-20

R61_137 V61 V137 -2878.183721525228
L61_137 V61 V137 4.384058122659104e-12
C61_137 V61 V137 2.1591235885679164e-19

R61_138 V61 V138 13014.01664177767
L61_138 V61 V138 -4.678348030447604e-12
C61_138 V61 V138 -2.9518774352070734e-20

R61_139 V61 V139 -4785.766829021505
L61_139 V61 V139 1.0052832786362529e-11
C61_139 V61 V139 4.2918879286797834e-20

R61_140 V61 V140 -2259.7230309059237
L61_140 V61 V140 2.6394039517806414e-11
C61_140 V61 V140 1.2255316275956487e-19

R61_141 V61 V141 -10405.224772512765
L61_141 V61 V141 -2.7035062316973913e-12
C61_141 V61 V141 -4.749771611445679e-19

R61_142 V61 V142 11224.661832604916
L61_142 V61 V142 6.0224509444631e-12
C61_142 V61 V142 -1.0282125228782429e-20

R61_143 V61 V143 -4870.922488350268
L61_143 V61 V143 -3.960546915443806e-11
C61_143 V61 V143 -2.5547901101277145e-20

R61_144 V61 V144 85516.42507362035
L61_144 V61 V144 1.9869008051564938e-11
C61_144 V61 V144 -1.8006729855306853e-19

R61_145 V61 V145 1058.990564129483
L61_145 V61 V145 -2.512126565432429e-12
C61_145 V61 V145 -2.5535496790187523e-19

R61_146 V61 V146 -11135.941084159205
L61_146 V61 V146 4.531718700109397e-12
C61_146 V61 V146 5.069633580429347e-20

R61_147 V61 V147 2458.2796754935343
L61_147 V61 V147 -4.094033634334592e-12
C61_147 V61 V147 -2.4257812374245307e-19

R61_148 V61 V148 6346.109342263874
L61_148 V61 V148 -2.3768057548774578e-12
C61_148 V61 V148 -1.4900268712079532e-19

R61_149 V61 V149 -912.1006779157801
L61_149 V61 V149 1.4732220828099983e-12
C61_149 V61 V149 4.391205169579359e-19

R61_150 V61 V150 -2744.473796803313
L61_150 V61 V150 -2.1369476630776245e-12
C61_150 V61 V150 -2.1895403652739385e-19

R61_151 V61 V151 6572.487010215366
L61_151 V61 V151 -7.89292783693813e-12
C61_151 V61 V151 7.024900703914619e-20

R61_152 V61 V152 6652.364189089107
L61_152 V61 V152 2.062290352019199e-11
C61_152 V61 V152 8.990268710667916e-20

R61_153 V61 V153 2622.974807932513
L61_153 V61 V153 3.145376844467743e-12
C61_153 V61 V153 3.0784645846116667e-19

R61_154 V61 V154 6223.539572496438
L61_154 V61 V154 6.083140011468601e-12
C61_154 V61 V154 1.897684079040043e-19

R61_155 V61 V155 -64754.261281807216
L61_155 V61 V155 1.8650307270017167e-12
C61_155 V61 V155 2.6209435575518126e-20

R61_156 V61 V156 -1908.0447624789288
L61_156 V61 V156 5.341714854010809e-12
C61_156 V61 V156 1.9886342427242167e-19

R61_157 V61 V157 1036.8893507553605
L61_157 V61 V157 -1.9687890759920577e-12
C61_157 V61 V157 -2.197845330968134e-19

R61_158 V61 V158 20606.55034334261
L61_158 V61 V158 3.5709399587357976e-12
C61_158 V61 V158 7.453192503236869e-20

R61_159 V61 V159 -2683.416169845479
L61_159 V61 V159 8.49988508188545e-12
C61_159 V61 V159 1.9131097533712148e-19

R61_160 V61 V160 18736.37732165642
L61_160 V61 V160 2.8646676225547943e-12
C61_160 V61 V160 1.392180721272274e-20

R61_161 V61 V161 -2900.3211071678998
L61_161 V61 V161 -2.7882172973253463e-12
C61_161 V61 V161 -2.690807280216949e-19

R61_162 V61 V162 -5425.132798879673
L61_162 V61 V162 1.091461543954457e-11
C61_162 V61 V162 1.200243734795935e-19

R61_163 V61 V163 -2663.7349071058693
L61_163 V61 V163 -3.130288935228111e-12
C61_163 V61 V163 1.4808370972384035e-20

R61_164 V61 V164 -2939.2912646309933
L61_164 V61 V164 -1.971136012373383e-12
C61_164 V61 V164 -1.2101584975844318e-20

R61_165 V61 V165 1263.2405308817567
L61_165 V61 V165 -1.4104044082374145e-11
C61_165 V61 V165 -2.5387923223339165e-21

R61_166 V61 V166 -3356.599398991123
L61_166 V61 V166 -1.7047661872415746e-12
C61_166 V61 V166 -2.310180899594196e-19

R61_167 V61 V167 -22363.168021815916
L61_167 V61 V167 -1.1257444042856608e-11
C61_167 V61 V167 -1.2631563764611584e-19

R61_168 V61 V168 -6423.973534548513
L61_168 V61 V168 -1.5239459898667375e-11
C61_168 V61 V168 -2.9482541738207045e-19

R61_169 V61 V169 5818.331470758271
L61_169 V61 V169 1.7247307157010648e-12
C61_169 V61 V169 3.3094580738971715e-19

R61_170 V61 V170 2882.6167476794517
L61_170 V61 V170 3.0813381356718707e-12
C61_170 V61 V170 6.804246116713039e-20

R61_171 V61 V171 1595.8616533197862
L61_171 V61 V171 4.001828162056196e-12
C61_171 V61 V171 -2.555685335189852e-20

R61_172 V61 V172 2705.7828746418945
L61_172 V61 V172 9.870738183099999e-12
C61_172 V61 V172 1.0806375017734214e-19

R61_173 V61 V173 -1984.2503697694028
L61_173 V61 V173 2.8766753381976747e-11
C61_173 V61 V173 4.684995330819892e-20

R61_174 V61 V174 6090.952145779112
L61_174 V61 V174 1.7509460036028684e-12
C61_174 V61 V174 2.30414364217558e-19

R61_175 V61 V175 -5230.478185229957
L61_175 V61 V175 3.00201171117499e-12
C61_175 V61 V175 2.728209798200017e-19

R61_176 V61 V176 -35876.85026432764
L61_176 V61 V176 2.075997953949326e-12
C61_176 V61 V176 3.4182338322049684e-19

R61_177 V61 V177 1386.4558213084065
L61_177 V61 V177 -1.6297820905241107e-12
C61_177 V61 V177 -2.1036140954285941e-19

R61_178 V61 V178 -3211.4669160835006
L61_178 V61 V178 -2.091519407301364e-12
C61_178 V61 V178 -1.0341616209089421e-19

R61_179 V61 V179 -2879.37411565275
L61_179 V61 V179 -2.713125507622759e-12
C61_179 V61 V179 -1.7250536348088678e-19

R61_180 V61 V180 -2591.168830615605
L61_180 V61 V180 -2.4506275630581872e-12
C61_180 V61 V180 -2.3082096195327023e-19

R61_181 V61 V181 -1011.4856774264169
L61_181 V61 V181 8.387211380282428e-12
C61_181 V61 V181 -2.626899950265554e-19

R61_182 V61 V182 3461.4808571067783
L61_182 V61 V182 6.7584954499828474e-12
C61_182 V61 V182 3.6327407609832943e-20

R61_183 V61 V183 40188.08145657928
L61_183 V61 V183 -3.5037638176771795e-12
C61_183 V61 V183 -8.540821195737353e-21

R61_184 V61 V184 8092.464835872626
L61_184 V61 V184 -2.8457162767440602e-12
C61_184 V61 V184 -6.038736965657612e-20

R61_185 V61 V185 2748.1945248955412
L61_185 V61 V185 4.804637079574043e-12
C61_185 V61 V185 3.381980555634817e-19

R61_186 V61 V186 5388.97154413269
L61_186 V61 V186 -4.694467554077498e-12
C61_186 V61 V186 -1.8352135749286098e-19

R61_187 V61 V187 2299.4636511754297
L61_187 V61 V187 4.193598050791072e-12
C61_187 V61 V187 6.192112550927725e-20

R61_188 V61 V188 1414.5028215534803
L61_188 V61 V188 2.1827066517668265e-12
C61_188 V61 V188 8.179324302123786e-21

R61_189 V61 V189 -41503.10713543309
L61_189 V61 V189 3.946532150358681e-12
C61_189 V61 V189 7.63376686245635e-20

R61_190 V61 V190 -2850.765544297541
L61_190 V61 V190 4.753802718354401e-11
C61_190 V61 V190 -1.748535147288984e-20

R61_191 V61 V191 9214.572047428563
L61_191 V61 V191 2.851397408244973e-12
C61_191 V61 V191 9.812374745511844e-21

R61_192 V61 V192 -5236.050055817624
L61_192 V61 V192 6.71571253430839e-12
C61_192 V61 V192 1.2357193461644081e-19

R61_193 V61 V193 -3818.6678927525795
L61_193 V61 V193 -7.234818963406504e-12
C61_193 V61 V193 1.4077741315172982e-20

R61_194 V61 V194 -18407.240709512185
L61_194 V61 V194 2.104870136060959e-12
C61_194 V61 V194 2.3187596345716393e-19

R61_195 V61 V195 -3625.6055166770134
L61_195 V61 V195 -2.787139013305102e-12
C61_195 V61 V195 -5.727190834795111e-20

R61_196 V61 V196 -4162.054937403379
L61_196 V61 V196 3.646206977684846e-11
C61_196 V61 V196 7.528684684638241e-20

R61_197 V61 V197 5660.427428466282
L61_197 V61 V197 -2.573999423378903e-12
C61_197 V61 V197 -2.831004853695403e-19

R61_198 V61 V198 5049.968185261463
L61_198 V61 V198 -3.717465101388802e-12
C61_198 V61 V198 -3.026421867754938e-20

R61_199 V61 V199 -15519.81101000374
L61_199 V61 V199 -2.9111624848160373e-12
C61_199 V61 V199 1.0208497814525234e-19

R61_200 V61 V200 5015.178534160183
L61_200 V61 V200 -1.9400420472992043e-12
C61_200 V61 V200 -1.876571256067441e-19

R62_62 V62 0 -338.5620297070609
L62_62 V62 0 6.941117014994514e-13
C62_62 V62 0 1.3387460148802454e-18

R62_63 V62 V63 55909.356476577595
L62_63 V62 V63 1.542677612369033e-11
C62_63 V62 V63 4.70661324065378e-20

R62_64 V62 V64 10612.293941466303
L62_64 V62 V64 -2.525805548134491e-11
C62_64 V62 V64 4.992010471213703e-21

R62_65 V62 V65 142060.3451144707
L62_65 V62 V65 -1.2709562739340642e-11
C62_65 V62 V65 -6.609058139682644e-20

R62_66 V62 V66 3370.3771027609746
L62_66 V62 V66 1.5765552370757698e-12
C62_66 V62 V66 3.329976579642094e-19

R62_67 V62 V67 7902.828531577218
L62_67 V62 V67 8.730991705702165e-12
C62_67 V62 V67 1.1589408025085543e-19

R62_68 V62 V68 5386.321935768783
L62_68 V62 V68 -5.553484019369235e-11
C62_68 V62 V68 7.333906018787832e-20

R62_69 V62 V69 -36349.517066735716
L62_69 V62 V69 3.1213647416557254e-12
C62_69 V62 V69 1.9290714086364035e-19

R62_70 V62 V70 2135.216217580452
L62_70 V62 V70 9.040263697166308e-13
C62_70 V62 V70 6.781084086237999e-19

R62_71 V62 V71 14985.882714578502
L62_71 V62 V71 -5.551926585855004e-12
C62_71 V62 V71 -1.3466943903653627e-19

R62_72 V62 V72 8914.214469865672
L62_72 V62 V72 -3.086140067945911e-11
C62_72 V62 V72 -6.141337142053862e-20

R62_73 V62 V73 3799.9257848138323
L62_73 V62 V73 5.765416036285644e-11
C62_73 V62 V73 -3.246730652785272e-20

R62_74 V62 V74 -2296.704248165552
L62_74 V62 V74 -1.2360100652159663e-12
C62_74 V62 V74 -4.6784254582881e-19

R62_75 V62 V75 -23746.409257518728
L62_75 V62 V75 1.4549798592796838e-11
C62_75 V62 V75 -6.43311805284491e-21

R62_76 V62 V76 -4107.813820237215
L62_76 V62 V76 2.6522275823796782e-12
C62_76 V62 V76 2.0294881928916127e-19

R62_77 V62 V77 -6580.733146971089
L62_77 V62 V77 -6.201182336449495e-12
C62_77 V62 V77 -1.0110415860388237e-19

R62_78 V62 V78 -10718.388159952625
L62_78 V62 V78 -1.051816148297222e-11
C62_78 V62 V78 6.229533249967066e-20

R62_79 V62 V79 -3980.096505733713
L62_79 V62 V79 2.7157682976401258e-11
C62_79 V62 V79 7.257950361721366e-20

R62_80 V62 V80 -5360.953096145022
L62_80 V62 V80 -3.640576319480208e-12
C62_80 V62 V80 -7.795851282913347e-20

R62_81 V62 V81 -27945.791692421015
L62_81 V62 V81 -1.551938426912632e-11
C62_81 V62 V81 -8.376792729078717e-20

R62_82 V62 V82 7645.9392060189875
L62_82 V62 V82 1.2662039780422499e-11
C62_82 V62 V82 -6.81073960440766e-20

R62_83 V62 V83 6687.748552303808
L62_83 V62 V83 -2.4836289843105108e-11
C62_83 V62 V83 -5.459166886875207e-20

R62_84 V62 V84 5139.805626903801
L62_84 V62 V84 -3.3117976964302225e-12
C62_84 V62 V84 -1.9815801534217227e-19

R62_85 V62 V85 -18359.702286378884
L62_85 V62 V85 -8.622418445749733e-12
C62_85 V62 V85 -3.764247723580807e-20

R62_86 V62 V86 1240.937425255975
L62_86 V62 V86 -2.6655797605870077e-11
C62_86 V62 V86 -2.5242527847460046e-19

R62_87 V62 V87 5959.127197980745
L62_87 V62 V87 4.524099001752457e-12
C62_87 V62 V87 1.7384407254616896e-19

R62_88 V62 V88 5830.569605473116
L62_88 V62 V88 2.1402043891815025e-12
C62_88 V62 V88 3.0343059948722046e-19

R62_89 V62 V89 5662.827026560409
L62_89 V62 V89 2.008132457777139e-12
C62_89 V62 V89 2.641800025257466e-19

R62_90 V62 V90 -1386.638023554208
L62_90 V62 V90 1.5722843174768557e-12
C62_90 V62 V90 6.803163372133487e-19

R62_91 V62 V91 -6834.224149146493
L62_91 V62 V91 -2.0842866426556745e-12
C62_91 V62 V91 -2.73622981023102e-19

R62_92 V62 V92 -5338.213970623699
L62_92 V62 V92 -2.5602878855809904e-12
C62_92 V62 V92 -1.555794288129814e-19

R62_93 V62 V93 -23573.609885560323
L62_93 V62 V93 -1.9093086515747057e-11
C62_93 V62 V93 -5.724034247810079e-20

R62_94 V62 V94 -3921.6402925051357
L62_94 V62 V94 -3.1775141733981303e-12
C62_94 V62 V94 -2.4195918461700934e-19

R62_95 V62 V95 -5688.246979584987
L62_95 V62 V95 -6.4223297211472645e-12
C62_95 V62 V95 -1.7060134061826855e-19

R62_96 V62 V96 -3607.5535662123198
L62_96 V62 V96 -5.069649604670846e-12
C62_96 V62 V96 -2.3790989781921136e-19

R62_97 V62 V97 -2502.18946510788
L62_97 V62 V97 -1.6882223852313602e-12
C62_97 V62 V97 -4.1844371471256786e-19

R62_98 V62 V98 1720.9480391040033
L62_98 V62 V98 -1.839835164337183e-12
C62_98 V62 V98 -3.8927294758805787e-19

R62_99 V62 V99 11284.101725417597
L62_99 V62 V99 1.2435324654294772e-12
C62_99 V62 V99 5.202230412901803e-19

R62_100 V62 V100 5246.994463721561
L62_100 V62 V100 2.1274384421476697e-12
C62_100 V62 V100 3.9035455111956743e-19

R62_101 V62 V101 3035.646244564604
L62_101 V62 V101 2.9053116362957506e-12
C62_101 V62 V101 2.7669132343598927e-19

R62_102 V62 V102 -2002.5677739379016
L62_102 V62 V102 2.031669994851157e-12
C62_102 V62 V102 3.3893653961177e-19

R62_103 V62 V103 5873.947746406712
L62_103 V62 V103 -6.1479144887280994e-12
C62_103 V62 V103 -6.933090409676308e-20

R62_104 V62 V104 5052.50810380652
L62_104 V62 V104 -4.913868259708248e-12
C62_104 V62 V104 -9.408820764798128e-20

R62_105 V62 V105 5534.238081232643
L62_105 V62 V105 2.2073074539683836e-12
C62_105 V62 V105 1.5879447155594208e-19

R62_106 V62 V106 738.7679498047391
L62_106 V62 V106 2.6907215944341975e-12
C62_106 V62 V106 6.087076967662889e-20

R62_107 V62 V107 -10940.752225983371
L62_107 V62 V107 -1.8044353576186908e-12
C62_107 V62 V107 -3.4658531232861953e-19

R62_108 V62 V108 -8726.07718004734
L62_108 V62 V108 -3.198627592012385e-11
C62_108 V62 V108 -4.8437460062842974e-20

R62_109 V62 V109 -1774.7355772525084
L62_109 V62 V109 -2.5625727321208796e-12
C62_109 V62 V109 -3.080258963821178e-19

R62_110 V62 V110 -1022.4067978252178
L62_110 V62 V110 -4.362297724807964e-12
C62_110 V62 V110 7.171182794499746e-20

R62_111 V62 V111 2698.906128498818
L62_111 V62 V111 6.7247840509075305e-12
C62_111 V62 V111 2.953516909434563e-20

R62_112 V62 V112 4493.87729342982
L62_112 V62 V112 -1.9994727583428056e-11
C62_112 V62 V112 -1.0558657470589536e-19

R62_113 V62 V113 -173466.43027294357
L62_113 V62 V113 -2.3873605399409994e-12
C62_113 V62 V113 -1.0088902690251021e-19

R62_114 V62 V114 -929.6165515335618
L62_114 V62 V114 -1.5442486610193867e-12
C62_114 V62 V114 -4.468585805714411e-19

R62_115 V62 V115 -1953.9712011367003
L62_115 V62 V115 2.1566398758920064e-12
C62_115 V62 V115 2.498041419333737e-19

R62_116 V62 V116 -2530.0038543039436
L62_116 V62 V116 4.3781324977204185e-12
C62_116 V62 V116 6.38585099415413e-20

R62_117 V62 V117 3571.98398049555
L62_117 V62 V117 2.4823571543282895e-12
C62_117 V62 V117 1.7153585973461802e-19

R62_118 V62 V118 480.8774010477893
L62_118 V62 V118 1.2207582760244454e-12
C62_118 V62 V118 3.65734765116971e-19

R62_119 V62 V119 2940.016081595685
L62_119 V62 V119 -1.690302970095331e-11
C62_119 V62 V119 6.931027182039891e-20

R62_120 V62 V120 2767.203271703305
L62_120 V62 V120 1.0702885069484405e-11
C62_120 V62 V120 2.665582573560742e-19

R62_121 V62 V121 -6658.917917734452
L62_121 V62 V121 3.422356262807321e-12
C62_121 V62 V121 5.494362935341691e-20

R62_122 V62 V122 -4505.120400534904
L62_122 V62 V122 -4.4244925188749814e-11
C62_122 V62 V122 5.594475664650139e-20

R62_123 V62 V123 2300.4965724475005
L62_123 V62 V123 -3.289257164440283e-12
C62_123 V62 V123 -2.624174342725735e-19

R62_124 V62 V124 3551.5321397304842
L62_124 V62 V124 -2.134099268207023e-12
C62_124 V62 V124 -4.375917838494082e-19

R62_125 V62 V125 7013.820972357809
L62_125 V62 V125 -6.511053157559828e-12
C62_125 V62 V125 -5.1701623053064885e-21

R62_126 V62 V126 -712.8292769179149
L62_126 V62 V126 -9.483166813067217e-13
C62_126 V62 V126 -4.485893870796008e-19

R62_127 V62 V127 -1178.117821892884
L62_127 V62 V127 -7.068616066560509e-12
C62_127 V62 V127 -5.779018804214713e-20

R62_128 V62 V128 -1360.6693494878623
L62_128 V62 V128 1.4206633687387088e-11
C62_128 V62 V128 -4.0607762586381863e-20

R62_129 V62 V129 -2816.765066319294
L62_129 V62 V129 -1.926378633629267e-12
C62_129 V62 V129 -3.64009092865984e-19

R62_130 V62 V130 1644.874417189316
L62_130 V62 V130 1.2021500729038942e-12
C62_130 V62 V130 4.031422210648104e-19

R62_131 V62 V131 1366.2376685152578
L62_131 V62 V131 2.662856423947232e-12
C62_131 V62 V131 2.3186183718909473e-19

R62_132 V62 V132 1129.5087956901275
L62_132 V62 V132 2.0810785249055372e-12
C62_132 V62 V132 4.2961705840666727e-19

R62_133 V62 V133 -75679.04394174344
L62_133 V62 V133 2.228810706686231e-12
C62_133 V62 V133 2.7308347612758294e-19

R62_134 V62 V134 1503.3245169134223
L62_134 V62 V134 -5.596228487280441e-12
C62_134 V62 V134 -1.8619133515765904e-19

R62_135 V62 V135 3437.505328221848
L62_135 V62 V135 2.582525071084085e-11
C62_135 V62 V135 -1.256446243982432e-19

R62_136 V62 V136 2103.6245190204827
L62_136 V62 V136 -7.656402883934253e-12
C62_136 V62 V136 -3.130086350743384e-19

R62_137 V62 V137 2204.997168706392
L62_137 V62 V137 3.1882478179906474e-12
C62_137 V62 V137 2.262461663498869e-19

R62_138 V62 V138 -1215.516188310068
L62_138 V62 V138 -2.577359497446859e-12
C62_138 V62 V138 -1.0327144434579181e-19

R62_139 V62 V139 -1013.7910670502544
L62_139 V62 V139 -1.0402063390811732e-11
C62_139 V62 V139 1.8952241944973438e-19

R62_140 V62 V140 -900.6685759583565
L62_140 V62 V140 -3.52110634869134e-12
C62_140 V62 V140 2.2165563876536187e-19

R62_141 V62 V141 7836.933757826193
L62_141 V62 V141 -1.6877169551196206e-12
C62_141 V62 V141 -4.990089182348564e-19

R62_142 V62 V142 -1084.6144441060044
L62_142 V62 V142 2.458967671743695e-12
C62_142 V62 V142 2.1610873545247246e-19

R62_143 V62 V143 1399.2278535552978
L62_143 V62 V143 -7.598228650589877e-12
C62_143 V62 V143 -1.6622483418729116e-19

R62_144 V62 V144 8830.31523696652
L62_144 V62 V144 4.554779427797072e-12
C62_144 V62 V144 -5.663497484805236e-20

R62_145 V62 V145 -2362.8143190331834
L62_145 V62 V145 -4.089208721517403e-12
C62_145 V62 V145 -1.8728773959738368e-19

R62_146 V62 V146 426.5836166244988
L62_146 V62 V146 -3.5641856161573075e-12
C62_146 V62 V146 -4.9047295536912395e-20

R62_147 V62 V147 -2940.9217205047344
L62_147 V62 V147 -6.590905027889434e-11
C62_147 V62 V147 -2.42556394422768e-19

R62_148 V62 V148 919.6188479134032
L62_148 V62 V148 -3.0596751750980126e-12
C62_148 V62 V148 -2.207106105239134e-19

R62_149 V62 V149 5431.93540399119
L62_149 V62 V149 7.689295943099726e-13
C62_149 V62 V149 8.311376852045434e-19

R62_150 V62 V150 -10952.305958956618
L62_150 V62 V150 4.498194800277522e-12
C62_150 V62 V150 -4.418472135444765e-19

R62_151 V62 V151 4187.597099502444
L62_151 V62 V151 -1.703726720479404e-11
C62_151 V62 V151 2.163988085295223e-19

R62_152 V62 V152 -705.0378491611989
L62_152 V62 V152 -1.5444732441764674e-11
C62_152 V62 V152 4.031045383241736e-20

R62_153 V62 V153 -12554.204204476557
L62_153 V62 V153 -1.98301601550679e-11
C62_153 V62 V153 2.3466477524385175e-20

R62_154 V62 V154 -888.0080841033861
L62_154 V62 V154 7.43699273145457e-11
C62_154 V62 V154 2.9572460612886597e-19

R62_155 V62 V155 -581.2379505793392
L62_155 V62 V155 2.6236989944896326e-12
C62_155 V62 V155 1.935085013991561e-19

R62_156 V62 V156 777.158052182377
L62_156 V62 V156 -1.753572510833953e-11
C62_156 V62 V156 2.4430739036261304e-19

R62_157 V62 V157 -4825.02616964941
L62_157 V62 V157 -8.221821423166531e-13
C62_157 V62 V157 -8.294240690750504e-19

R62_158 V62 V158 2435.3910262906024
L62_158 V62 V158 -8.110761010223707e-12
C62_158 V62 V158 8.962484561865864e-20

R62_159 V62 V159 513.7292850957402
L62_159 V62 V159 8.437268745063975e-12
C62_159 V62 V159 -6.485095318260569e-20

R62_160 V62 V160 2063.712902940042
L62_160 V62 V160 1.9558718117292846e-12
C62_160 V62 V160 -4.061206999245962e-20

R62_161 V62 V161 -2247.230650299691
L62_161 V62 V161 -1.123647263984215e-11
C62_161 V62 V161 9.50791542656554e-20

R62_162 V62 V162 1284.6485393542198
L62_162 V62 V162 -4.879809702070389e-12
C62_162 V62 V162 2.123060337309393e-20

R62_163 V62 V163 -2375.227288819677
L62_163 V62 V163 -2.3561106471650914e-12
C62_163 V62 V163 -1.132745183036304e-19

R62_164 V62 V164 -15541.607516489283
L62_164 V62 V164 -2.4111837755623334e-12
C62_164 V62 V164 4.030640398705213e-20

R62_165 V62 V165 1134.9729300752456
L62_165 V62 V165 1.3676345067699768e-12
C62_165 V62 V165 3.416995104578728e-19

R62_166 V62 V166 13944.875894304254
L62_166 V62 V166 1.952639910769721e-12
C62_166 V62 V166 -1.2538697158284831e-19

R62_167 V62 V167 7619.8365764757955
L62_167 V62 V167 -2.442646236706191e-12
C62_167 V62 V167 4.1885018007084535e-20

R62_168 V62 V168 -965.4999674989423
L62_168 V62 V168 -2.154327577877613e-12
C62_168 V62 V168 -7.850862957123814e-20

R62_169 V62 V169 2186.819830255
L62_169 V62 V169 8.703332492498539e-12
C62_169 V62 V169 -1.7321000173302052e-19

R62_170 V62 V170 -5295.616018021458
L62_170 V62 V170 1.4865025606769265e-12
C62_170 V62 V170 2.4852992693923286e-19

R62_171 V62 V171 -9658.485873791675
L62_171 V62 V171 1.0439296687968466e-12
C62_171 V62 V171 2.0842127696442413e-19

R62_172 V62 V172 1528.3585023215874
L62_172 V62 V172 1.8653220952990982e-12
C62_172 V62 V172 1.129806398267922e-19

R62_173 V62 V173 -1529.3710320921084
L62_173 V62 V173 -2.320488618152912e-12
C62_173 V62 V173 -5.0263760155135867e-20

R62_174 V62 V174 -1884.6618651011258
L62_174 V62 V174 -7.563082908598617e-13
C62_174 V62 V174 -2.6624815318786187e-19

R62_175 V62 V175 3827.4424612894227
L62_175 V62 V175 1.0695029488448611e-11
C62_175 V62 V175 9.914164535651213e-20

R62_176 V62 V176 8283.370582912286
L62_176 V62 V176 3.639940391574732e-12
C62_176 V62 V176 1.4198883916757874e-19

R62_177 V62 V177 1860.7196690455023
L62_177 V62 V177 -3.957934235736119e-11
C62_177 V62 V177 6.615930378628179e-20

R62_178 V62 V178 2261.5580777642062
L62_178 V62 V178 -1.1434906646429467e-11
C62_178 V62 V178 -6.219005543104276e-20

R62_179 V62 V179 -1789.4139017166697
L62_179 V62 V179 -1.398833752888565e-12
C62_179 V62 V179 -3.752752303798996e-19

R62_180 V62 V180 -6257.71353104918
L62_180 V62 V180 -1.3625315329508357e-12
C62_180 V62 V180 -3.1547345796867516e-19

R62_181 V62 V181 52321.336926979566
L62_181 V62 V181 1.620122260126344e-11
C62_181 V62 V181 -8.359628496336662e-20

R62_182 V62 V182 -16382.890573567904
L62_182 V62 V182 6.764570592056858e-13
C62_182 V62 V182 2.0513048061829296e-19

R62_183 V62 V183 1440.3448701291193
L62_183 V62 V183 -4.0878262924568926e-12
C62_183 V62 V183 -4.521272810747274e-20

R62_184 V62 V184 3001.5778283727022
L62_184 V62 V184 -6.6483388480480614e-12
C62_184 V62 V184 2.8392042895464286e-20

R62_185 V62 V185 -2661.769593981042
L62_185 V62 V185 1.1715807014965895e-11
C62_185 V62 V185 4.2590312410005174e-20

R62_186 V62 V186 -5069.736139126896
L62_186 V62 V186 -1.5870908607520332e-12
C62_186 V62 V186 -1.0821834415285443e-19

R62_187 V62 V187 -5991.755262483696
L62_187 V62 V187 2.953470645675231e-12
C62_187 V62 V187 3.16728688981269e-19

R62_188 V62 V188 -1037.8626382740251
L62_188 V62 V188 1.3565615433622548e-12
C62_188 V62 V188 2.729699819693003e-19

R62_189 V62 V189 2500.7922803296815
L62_189 V62 V189 5.300301175993834e-12
C62_189 V62 V189 1.4587436570243825e-19

R62_190 V62 V190 3165.7212823384853
L62_190 V62 V190 -2.7936497845581267e-12
C62_190 V62 V190 -1.347932656726424e-19

R62_191 V62 V191 -1906.4797367007454
L62_191 V62 V191 1.6870188745534083e-12
C62_191 V62 V191 1.162460255658907e-19

R62_192 V62 V192 11862.325554947249
L62_192 V62 V192 2.802165702071651e-11
C62_192 V62 V192 -3.6744629095242224e-20

R62_193 V62 V193 -7212.438307895659
L62_193 V62 V193 -4.9053599131514116e-12
C62_193 V62 V193 -1.5491530439221386e-19

R62_194 V62 V194 -3930.0834952282803
L62_194 V62 V194 -7.694311019698696e-12
C62_194 V62 V194 -1.9576812025362017e-19

R62_195 V62 V195 1919.5703570877
L62_195 V62 V195 -1.3233856663725749e-12
C62_195 V62 V195 -3.11788833004032e-19

R62_196 V62 V196 1300.3738834757173
L62_196 V62 V196 -1.7696351006873155e-12
C62_196 V62 V196 -8.765070724474698e-20

R62_197 V62 V197 -4094.624982507198
L62_197 V62 V197 -1.104673031304076e-11
C62_197 V62 V197 -5.0888649419433526e-20

R62_198 V62 V198 -58920.00728133265
L62_198 V62 V198 2.8973409553038332e-12
C62_198 V62 V198 7.295711529647453e-20

R62_199 V62 V199 2209.001791477626
L62_199 V62 V199 -4.8658463031190515e-12
C62_199 V62 V199 -6.57017068341488e-20

R62_200 V62 V200 -2442.4298289857848
L62_200 V62 V200 -7.604147395316324e-12
C62_200 V62 V200 -3.428190517114204e-21

R63_63 V63 0 -3477.05111564273
L63_63 V63 0 -8.770626576604855e-13
C63_63 V63 0 -5.058426944966197e-19

R63_64 V63 V64 -9273.677086731717
L63_64 V63 V64 -1.459545500244817e-11
C63_64 V63 V64 -1.0585484315887292e-19

R63_65 V63 V65 33489.45247509936
L63_65 V63 V65 4.41233894505191e-12
C63_65 V63 V65 1.7125280929086538e-19

R63_66 V63 V66 -174610.63657606606
L63_66 V63 V66 -1.2493415488035942e-11
C63_66 V63 V66 -8.269615167024531e-21

R63_67 V63 V67 -35297.92848987641
L63_67 V63 V67 1.702214600120596e-12
C63_67 V63 V67 3.267929691652725e-19

R63_68 V63 V68 -14912.986792103226
L63_68 V63 V68 5.799901270315675e-11
C63_68 V63 V68 2.122409695679839e-20

R63_69 V63 V69 -38542.509552642456
L63_69 V63 V69 6.6735508030408e-12
C63_69 V63 V69 8.479308083667013e-20

R63_70 V63 V70 -48919.86828044892
L63_70 V63 V70 -8.620383575022952e-12
C63_70 V63 V70 -1.3966746061018527e-19

R63_71 V63 V71 4598.219116503032
L63_71 V63 V71 6.754278790698185e-13
C63_71 V63 V71 1.056170398052824e-18

R63_72 V63 V72 -159501.65823355794
L63_72 V63 V72 -2.944358163969148e-11
C63_72 V63 V72 -3.4123964460363114e-20

R63_73 V63 V73 7174.742070589123
L63_73 V63 V73 -4.162462668830755e-12
C63_73 V63 V73 -2.094444661551269e-19

R63_74 V63 V74 14091.438734975101
L63_74 V63 V74 9.026271821785559e-12
C63_74 V63 V74 8.48524027415114e-20

R63_75 V63 V75 -196541.24661310264
L63_75 V63 V75 -7.12996443724378e-13
C63_75 V63 V75 -9.61405235464033e-19

R63_76 V63 V76 6040.832857540848
L63_76 V63 V76 2.3714595352813335e-11
C63_76 V63 V76 1.2251313827625105e-20

R63_77 V63 V77 9856.804199807379
L63_77 V63 V77 1.4460612945817188e-11
C63_77 V63 V77 1.1650210426021119e-19

R63_78 V63 V78 -14046.342193891518
L63_78 V63 V78 1.323853514731027e-11
C63_78 V63 V78 1.125684389918509e-19

R63_79 V63 V79 -2774.1174818914947
L63_79 V63 V79 -4.0271813239792e-12
C63_79 V63 V79 -1.5535714924262793e-19

R63_80 V63 V80 -5253.786465434727
L63_80 V63 V80 -7.929124842432807e-11
C63_80 V63 V80 7.417624616906895e-20

R63_81 V63 V81 -3433.958791853616
L63_81 V63 V81 6.696396009541585e-12
C63_81 V63 V81 6.128878793617359e-20

R63_82 V63 V82 55651.7855075843
L63_82 V63 V82 -1.7127606922598543e-11
C63_82 V63 V82 -6.281734041597898e-20

R63_83 V63 V83 4913.824805978839
L63_83 V63 V83 9.719387106196836e-13
C63_83 V63 V83 7.029085789825475e-19

R63_84 V63 V84 41103.01763427227
L63_84 V63 V84 1.7486859719671194e-11
C63_84 V63 V84 1.593106692073395e-21

R63_85 V63 V85 17183.958531091226
L63_85 V63 V85 -2.3509593587801203e-09
C63_85 V63 V85 -1.1961393286171762e-20

R63_86 V63 V86 6706.592476107634
L63_86 V63 V86 8.270557952529988e-12
C63_86 V63 V86 2.04287272201158e-20

R63_87 V63 V87 1990.0462135307448
L63_87 V63 V87 -1.6267766492419087e-12
C63_87 V63 V87 -4.400069516105323e-19

R63_88 V63 V88 9363.454562825544
L63_88 V63 V88 3.4316678488387124e-11
C63_88 V63 V88 -2.122915817418925e-20

R63_89 V63 V89 3828.948443232701
L63_89 V63 V89 2.398579812327432e-11
C63_89 V63 V89 -3.093898902999853e-20

R63_90 V63 V90 -15761.178469198558
L63_90 V63 V90 -6.5310114165996825e-12
C63_90 V63 V90 -3.962753988256917e-20

R63_91 V63 V91 -969.7257655524387
L63_91 V63 V91 2.15274359833339e-12
C63_91 V63 V91 2.7454497480987657e-19

R63_92 V63 V92 -4399.694156427841
L63_92 V63 V92 9.361907374367074e-11
C63_92 V63 V92 4.42096798323235e-20

R63_93 V63 V93 -4356.015979829793
L63_93 V63 V93 -1.3051537786443336e-11
C63_93 V63 V93 -2.6177213512407585e-20

R63_94 V63 V94 -16069.895604951349
L63_94 V63 V94 -1.0611174042622951e-11
C63_94 V63 V94 -1.1925595442336914e-20

R63_95 V63 V95 -16491.105498882684
L63_95 V63 V95 4.05094598116848e-12
C63_95 V63 V95 2.41616558087464e-19

R63_96 V63 V96 8709.723591161835
L63_96 V63 V96 -1.0151120677589744e-11
C63_96 V63 V96 -1.5237593002194245e-20

R63_97 V63 V97 13516.716326565625
L63_97 V63 V97 4.1623206625297087e-11
C63_97 V63 V97 7.897402403484724e-20

R63_98 V63 V98 12663.30042795734
L63_98 V63 V98 3.795049571886427e-12
C63_98 V63 V98 9.970798182523895e-20

R63_99 V63 V99 895.4390442802902
L63_99 V63 V99 -1.0466137334201512e-12
C63_99 V63 V99 -5.581236437794994e-19

R63_100 V63 V100 15633.662586077227
L63_100 V63 V100 2.2475919220537627e-11
C63_100 V63 V100 -3.155594307457418e-20

R63_101 V63 V101 -4472354.33052082
L63_101 V63 V101 2.359050294397686e-10
C63_101 V63 V101 -6.598252580084559e-21

R63_102 V63 V102 11508.67532994355
L63_102 V63 V102 -1.3789297838353223e-11
C63_102 V63 V102 -3.8209166614009434e-20

R63_103 V63 V103 -1571.6490117104393
L63_103 V63 V103 1.6238482642873386e-12
C63_103 V63 V103 2.4529656155649395e-19

R63_104 V63 V104 -10821.146249278227
L63_104 V63 V104 1.0004644033171035e-11
C63_104 V63 V104 5.736053442075047e-20

R63_105 V63 V105 -27241.64032386338
L63_105 V63 V105 8.694050053284412e-12
C63_105 V63 V105 -5.187523892559793e-20

R63_106 V63 V106 -12452.177609519515
L63_106 V63 V106 -3.8426094879364864e-12
C63_106 V63 V106 -1.4149100595771925e-19

R63_107 V63 V107 -2155.3272726037108
L63_107 V63 V107 2.4203904071415048e-12
C63_107 V63 V107 1.895004256064946e-19

R63_108 V63 V108 -15784.058672140658
L63_108 V63 V108 -7.889364624736947e-12
C63_108 V63 V108 -3.8496203616267163e-20

R63_109 V63 V109 5341.095785250687
L63_109 V63 V109 7.10641154205577e-11
C63_109 V63 V109 4.618628323455183e-20

R63_110 V63 V110 9630.638466588007
L63_110 V63 V110 9.01150635456751e-12
C63_110 V63 V110 6.657624802342492e-20

R63_111 V63 V111 1322.7249212612294
L63_111 V63 V111 -1.7262124213849353e-12
C63_111 V63 V111 -1.184204418724054e-19

R63_112 V63 V112 6794.818764807365
L63_112 V63 V112 -2.6392332657028896e-11
C63_112 V63 V112 -3.976225327960467e-20

R63_113 V63 V113 -2604.7299101919634
L63_113 V63 V113 -8.988874393690267e-12
C63_113 V63 V113 3.642304217084038e-20

R63_114 V63 V114 -42306.35483151981
L63_114 V63 V114 8.37375551363463e-12
C63_114 V63 V114 9.69273371847599e-20

R63_115 V63 V115 6082.819765067229
L63_115 V63 V115 -5.0906620436748855e-12
C63_115 V63 V115 -1.0716702103942389e-19

R63_116 V63 V116 5131.501508215243
L63_116 V63 V116 6.1618481417100866e-12
C63_116 V63 V116 6.674357710134219e-20

R63_117 V63 V117 6341.514029091615
L63_117 V63 V117 -1.4214502097647984e-11
C63_117 V63 V117 -7.342017208255279e-20

R63_118 V63 V118 -10359.262387532459
L63_118 V63 V118 8.39683772696196e-12
C63_118 V63 V118 -4.263569032054838e-20

R63_119 V63 V119 -1744.547558044999
L63_119 V63 V119 1.2474545809987353e-12
C63_119 V63 V119 -5.979853477598086e-20

R63_120 V63 V120 -1726.683482556583
L63_120 V63 V120 -1.456109438282436e-11
C63_120 V63 V120 -4.83545020243046e-20

R63_121 V63 V121 5678.444067566011
L63_121 V63 V121 4.227499039683107e-12
C63_121 V63 V121 8.636174820145681e-20

R63_122 V63 V122 12208.11793233151
L63_122 V63 V122 -4.248122306226306e-12
C63_122 V63 V122 -7.006420966057402e-20

R63_123 V63 V123 2717.0948961982035
L63_123 V63 V123 -3.3366853764462204e-12
C63_123 V63 V123 3.268530368860176e-19

R63_124 V63 V124 3021.8570674794328
L63_124 V63 V124 -8.510586573086928e-12
C63_124 V63 V124 -4.947691800407657e-21

R63_125 V63 V125 -2393.8445546827033
L63_125 V63 V125 8.094521009136911e-12
C63_125 V63 V125 -1.930164009885714e-21

R63_126 V63 V126 -24094.808659175353
L63_126 V63 V126 -1.4099577676514108e-11
C63_126 V63 V126 3.7991041026341084e-20

R63_127 V63 V127 -4629.668264581667
L63_127 V63 V127 -1.04182485163307e-12
C63_127 V63 V127 -1.2882302781727684e-19

R63_128 V63 V128 2443.5698045742106
L63_128 V63 V128 -2.2624571531968625e-11
C63_128 V63 V128 3.540163007654457e-20

R63_129 V63 V129 4180.014557412066
L63_129 V63 V129 -2.900854942167543e-12
C63_129 V63 V129 -3.0545124032715504e-20

R63_130 V63 V130 28111.99737801079
L63_130 V63 V130 5.110728367225922e-12
C63_130 V63 V130 4.0352608965202907e-20

R63_131 V63 V131 4059.797761742634
L63_131 V63 V131 1.0568619641471322e-12
C63_131 V63 V131 -1.41833466053296e-19

R63_132 V63 V132 -1912.6340218404102
L63_132 V63 V132 2.5562318345143107e-12
C63_132 V63 V132 -8.40123569352958e-20

R63_133 V63 V133 8528.286971766236
L63_133 V63 V133 7.2124692238362415e-12
C63_133 V63 V133 1.705912069641031e-20

R63_134 V63 V134 -2710.3597312922498
L63_134 V63 V134 1.9810432680021897e-11
C63_134 V63 V134 -8.814261538129053e-20

R63_135 V63 V135 2051.9334315255846
L63_135 V63 V135 5.55912618220812e-12
C63_135 V63 V135 3.4527679179684013e-19

R63_136 V63 V136 177164.8895939102
L63_136 V63 V136 6.33109378645356e-12
C63_136 V63 V136 -6.485551325944276e-21

R63_137 V63 V137 -2608.8144441776594
L63_137 V63 V137 8.300563560694108e-12
C63_137 V63 V137 -7.460991958185763e-21

R63_138 V63 V138 3900.5169716958344
L63_138 V63 V138 -7.087575563648649e-12
C63_138 V63 V138 9.895101895635072e-20

R63_139 V63 V139 -927.0353926874946
L63_139 V63 V139 -3.040596569030138e-12
C63_139 V63 V139 -3.7875346177160605e-19

R63_140 V63 V140 -4364.099531117366
L63_140 V63 V140 -1.610061631718393e-12
C63_140 V63 V140 3.1195771171766005e-20

R63_141 V63 V141 6405.515067347805
L63_141 V63 V141 3.108750837848775e-11
C63_141 V63 V141 3.8408816752654836e-20

R63_142 V63 V142 2386.4708948722086
L63_142 V63 V142 -3.3588229842938566e-12
C63_142 V63 V142 1.8183197944022182e-20

R63_143 V63 V143 3088.76470659254
L63_143 V63 V143 -4.7394578673138616e-11
C63_143 V63 V143 2.4722967580122053e-20

R63_144 V63 V144 2528.799393879789
L63_144 V63 V144 3.0941742572659246e-12
C63_144 V63 V144 -2.835863220207157e-20

R63_145 V63 V145 2247.1523881955964
L63_145 V63 V145 -2.704165809097424e-11
C63_145 V63 V145 3.8031451180671245e-20

R63_146 V63 V146 209455.84165930745
L63_146 V63 V146 1.9223621955663216e-12
C63_146 V63 V146 -7.855460165382922e-20

R63_147 V63 V147 1071.546563742165
L63_147 V63 V147 -4.279013455055137e-12
C63_147 V63 V147 2.8064102927450887e-19

R63_148 V63 V148 -5793.7053806001895
L63_148 V63 V148 2.2534834176511202e-11
C63_148 V63 V148 6.746490612888484e-21

R63_149 V63 V149 -3713.064029561174
L63_149 V63 V149 -1.8144510358828446e-11
C63_149 V63 V149 -6.975993646405417e-20

R63_150 V63 V150 -1314.1500721178754
L63_150 V63 V150 7.57127169384401e-12
C63_150 V63 V150 -1.8662121513770932e-20

R63_151 V63 V151 -1939.0272707166407
L63_151 V63 V151 3.053793049503789e-12
C63_151 V63 V151 -1.0925381114782044e-19

R63_152 V63 V152 -51770.38833987797
L63_152 V63 V152 -3.0599347908680026e-12
C63_152 V63 V152 1.0975812834653164e-20

R63_153 V63 V153 -1924.1943877636445
L63_153 V63 V153 1.473168798666241e-11
C63_153 V63 V153 9.760539533763399e-21

R63_154 V63 V154 8362.962460184252
L63_154 V63 V154 -4.061355908385838e-12
C63_154 V63 V154 7.341310261451316e-20

R63_155 V63 V155 -11021.462786971093
L63_155 V63 V155 3.2926375556581006e-12
C63_155 V63 V155 -1.0415007409257696e-19

R63_156 V63 V156 -3313.2713551176257
L63_156 V63 V156 -8.194511328356562e-12
C63_156 V63 V156 2.6922408671122075e-20

R63_157 V63 V157 5970.781215644222
L63_157 V63 V157 1.7397718656931808e-11
C63_157 V63 V157 -7.6284633549614e-21

R63_158 V63 V158 3294.123497380667
L63_158 V63 V158 -6.537831716005176e-11
C63_158 V63 V158 -3.487240151828805e-20

R63_159 V63 V159 6705.678820188368
L63_159 V63 V159 -1.949485525127072e-12
C63_159 V63 V159 1.400302714627227e-19

R63_160 V63 V160 2244.251559891687
L63_160 V63 V160 1.5343977428186517e-12
C63_160 V63 V160 -3.3263198999615764e-20

R63_161 V63 V161 12835.911231190317
L63_161 V63 V161 -3.026723028079109e-12
C63_161 V63 V161 3.2206719379041994e-21

R63_162 V63 V162 654987.4696664163
L63_162 V63 V162 -5.845597786565244e-11
C63_162 V63 V162 -8.348813422479035e-20

R63_163 V63 V163 -6047.749294749222
L63_163 V63 V163 -9.690771349956894e-13
C63_163 V63 V163 -1.157722890937337e-19

R63_164 V63 V164 -2220.2516410463754
L63_164 V63 V164 -2.0138120115874298e-12
C63_164 V63 V164 -2.765816164412314e-20

R63_165 V63 V165 -8152.6155727442865
L63_165 V63 V165 3.969235186368503e-12
C63_165 V63 V165 8.350852055352855e-20

R63_166 V63 V166 -2185.430781595952
L63_166 V63 V166 -4.053367127799572e-12
C63_166 V63 V166 6.338003791127354e-20

R63_167 V63 V167 -3410.6514567626605
L63_167 V63 V167 5.916466536900451e-13
C63_167 V63 V167 -1.9153089621874174e-21

R63_168 V63 V168 4938.686379157937
L63_168 V63 V168 -2.274788732789856e-12
C63_168 V63 V168 -9.579686498027746e-22

R63_169 V63 V169 -30084.36737155314
L63_169 V63 V169 4.882110552401965e-12
C63_169 V63 V169 5.3095410909285077e-20

R63_170 V63 V170 2815.3732431825592
L63_170 V63 V170 4.533166226561631e-12
C63_170 V63 V170 1.7980751345134466e-20

R63_171 V63 V171 1458.3989091929425
L63_171 V63 V171 -2.9848669498156037e-11
C63_171 V63 V171 1.296838108910678e-19

R63_172 V63 V172 3415.077922749019
L63_172 V63 V172 2.469524642647295e-12
C63_172 V63 V172 4.382105249543439e-20

R63_173 V63 V173 9326.725183175055
L63_173 V63 V173 -2.742256242092028e-12
C63_173 V63 V173 -1.3057902927496027e-19

R63_174 V63 V174 3884.2522416911775
L63_174 V63 V174 4.7466123853102375e-12
C63_174 V63 V174 -4.365209594804988e-20

R63_175 V63 V175 -3240.09534993597
L63_175 V63 V175 -6.740934713196526e-13
C63_175 V63 V175 -2.3474066506427086e-19

R63_176 V63 V176 -5520.04386706316
L63_176 V63 V176 -1.1080123276897757e-11
C63_176 V63 V176 -2.574084032213376e-20

R63_177 V63 V177 -10856.40356766026
L63_177 V63 V177 1.2879388458377752e-11
C63_177 V63 V177 5.135263546407813e-20

R63_178 V63 V178 -2802.1845966254223
L63_178 V63 V178 -3.2908446925808196e-12
C63_178 V63 V178 3.4943392021966763e-22

R63_179 V63 V179 -2974.250225128337
L63_179 V63 V179 1.3017377786609794e-12
C63_179 V63 V179 1.4654680688794084e-19

R63_180 V63 V180 -4035.8266493885067
L63_180 V63 V180 -1.1390509132574867e-11
C63_180 V63 V180 -3.6815851201400106e-22

R63_181 V63 V181 -66097.95607465498
L63_181 V63 V181 7.678292337568336e-12
C63_181 V63 V181 4.3858416189155535e-20

R63_182 V63 V182 14286.647413573082
L63_182 V63 V182 2.2444052130553908e-11
C63_182 V63 V182 -3.8024458396696647e-22

R63_183 V63 V183 3160.2411822083714
L63_183 V63 V183 2.9361562871063967e-12
C63_183 V63 V183 -2.9213368842967984e-20

R63_184 V63 V184 7392.197117690388
L63_184 V63 V184 4.71031042794582e-12
C63_184 V63 V184 3.9717564520339195e-20

R63_185 V63 V185 10270.866991717146
L63_185 V63 V185 -1.2335896397494118e-10
C63_185 V63 V185 -4.94266434812052e-20

R63_186 V63 V186 4349.441331312304
L63_186 V63 V186 2.732486959062575e-12
C63_186 V63 V186 6.749487649538522e-20

R63_187 V63 V187 29859.84189082342
L63_187 V63 V187 -1.3507708425341382e-12
C63_187 V63 V187 -1.3921370519517326e-19

R63_188 V63 V188 2465.1170908887516
L63_188 V63 V188 -1.1514648246253816e-11
C63_188 V63 V188 -5.127277472418801e-21

R63_189 V63 V189 -9230.311836829025
L63_189 V63 V189 -7.720663476336452e-12
C63_189 V63 V189 5.970406680773862e-20

R63_190 V63 V190 -4619.676592850207
L63_190 V63 V190 -8.167234277641574e-12
C63_190 V63 V190 -2.709275290905162e-20

R63_191 V63 V191 -3755.592678494504
L63_191 V63 V191 5.121287235906511e-11
C63_191 V63 V191 1.9023930654099006e-19

R63_192 V63 V192 -3440.120490178767
L63_192 V63 V192 -4.744879224862961e-12
C63_192 V63 V192 -1.5942651215084377e-21

R63_193 V63 V193 112912.07075579598
L63_193 V63 V193 3.3026654218745705e-11
C63_193 V63 V193 -3.600815830232472e-20

R63_194 V63 V194 -5508.300222159766
L63_194 V63 V194 -1.2098794889800643e-11
C63_194 V63 V194 3.9702522248184756e-20

R63_195 V63 V195 6695.950551184784
L63_195 V63 V195 -1.210054684600184e-10
C63_195 V63 V195 -2.748402917770093e-19

R63_196 V63 V196 -6103.383945955348
L63_196 V63 V196 4.695379189283958e-12
C63_196 V63 V196 4.627447514586665e-20

R63_197 V63 V197 15855.738928919378
L63_197 V63 V197 2.8109975569813678e-11
C63_197 V63 V197 -1.55843903591068e-20

R63_198 V63 V198 6871.529170315842
L63_198 V63 V198 2.3781571567703127e-11
C63_198 V63 V198 -5.953173077632245e-21

R63_199 V63 V199 8710.602562021137
L63_199 V63 V199 6.05384970722735e-12
C63_199 V63 V199 -2.615128520462393e-21

R63_200 V63 V200 2080.466129553291
L63_200 V63 V200 -2.4399448774432535e-11
C63_200 V63 V200 -6.787569954611618e-20

R64_64 V64 0 773.4911455717157
L64_64 V64 0 -1.5625951845534523e-12
C64_64 V64 0 -3.4874479890910383e-20

R64_65 V64 V65 -25311.162284580434
L64_65 V64 V65 6.717727845238975e-12
C64_65 V64 V65 1.3676406390563825e-19

R64_66 V64 V66 -15610.500915373714
L64_66 V64 V66 -3.1342004861508296e-11
C64_66 V64 V66 7.128486279483033e-21

R64_67 V64 V67 -31142.035120635876
L64_67 V64 V67 -3.7429385116161414e-11
C64_67 V64 V67 -2.2318784046485955e-20

R64_68 V64 V68 -3312.5002484304555
L64_68 V64 V68 2.30101241607744e-12
C64_68 V64 V68 3.351922645922506e-19

R64_69 V64 V69 94384.75182761202
L64_69 V64 V69 3.359310574812082e-12
C64_69 V64 V69 1.6841365383651042e-19

R64_70 V64 V70 -18446.705387713093
L64_70 V64 V70 -7.651740417821161e-12
C64_70 V64 V70 -1.9152220121453503e-19

R64_71 V64 V71 -16618.689690775605
L64_71 V64 V71 -1.489130092389999e-11
C64_71 V64 V71 2.375284282094394e-21

R64_72 V64 V72 4075.6974262871026
L64_72 V64 V72 6.088888764179166e-13
C64_72 V64 V72 1.1997977617550293e-18

R64_73 V64 V73 9150.870153105474
L64_73 V64 V73 -4.567674374705615e-12
C64_73 V64 V73 -1.8351345094713794e-19

R64_74 V64 V74 5311.803367264723
L64_74 V64 V74 4.5517645829217114e-12
C64_74 V64 V74 1.7432999333820312e-19

R64_75 V64 V75 12207.482696885592
L64_75 V64 V75 1.2640347525713588e-11
C64_75 V64 V75 2.720686726833532e-20

R64_76 V64 V76 2152.4476413970565
L64_76 V64 V76 -7.976129145553283e-13
C64_76 V64 V76 -1.0401274764977269e-18

R64_77 V64 V77 4258.954293079278
L64_77 V64 V77 7.143649556485944e-12
C64_77 V64 V77 1.4342728279774338e-19

R64_78 V64 V78 -5389.673346904267
L64_78 V64 V78 1.3854335685571797e-11
C64_78 V64 V78 1.302431256892e-19

R64_79 V64 V79 37609.37074835058
L64_79 V64 V79 2.6544973572496837e-11
C64_79 V64 V79 4.483383542034824e-20

R64_80 V64 V80 -1467.7052563505586
L64_80 V64 V80 -4.421999555891402e-12
C64_80 V64 V80 -6.730146994936347e-20

R64_81 V64 V81 -1735.4410987051847
L64_81 V64 V81 -1.754225269062196e-11
C64_81 V64 V81 -4.8806890372884734e-20

R64_82 V64 V82 11222.333419467222
L64_82 V64 V82 -4.471100113364265e-12
C64_82 V64 V82 -1.7198997350614097e-19

R64_83 V64 V83 19856.439774944654
L64_83 V64 V83 1.2930362417387443e-11
C64_83 V64 V83 3.445947919638638e-20

R64_84 V64 V84 11990.486431547424
L64_84 V64 V84 1.4732913505751561e-12
C64_84 V64 V84 6.013022035945671e-19

R64_85 V64 V85 20375.8535433863
L64_85 V64 V85 -8.855890159235762e-12
C64_85 V64 V85 -6.23955199508415e-20

R64_86 V64 V86 24873.984671415248
L64_86 V64 V86 2.3953500137432407e-11
C64_86 V64 V86 4.389740303797757e-22

R64_87 V64 V87 7311.099925242762
L64_87 V64 V87 4.445085531480009e-11
C64_87 V64 V87 -3.174022833155906e-20

R64_88 V64 V88 1211.5876213465892
L64_88 V64 V88 -5.161063534936292e-12
C64_88 V64 V88 -3.6992379993293534e-19

R64_89 V64 V89 2459.5730276081463
L64_89 V64 V89 4.945748009103573e-12
C64_89 V64 V89 2.13157098738303e-20

R64_90 V64 V90 46160.688687160095
L64_90 V64 V90 3.864423572037148e-12
C64_90 V64 V90 1.2094115068233784e-19

R64_91 V64 V91 -1858.9778528135012
L64_91 V64 V91 -4.593163393898287e-12
C64_91 V64 V91 -1.928811570192527e-20

R64_92 V64 V92 -598.1451888339997
L64_92 V64 V92 4.0338280696532025e-11
C64_92 V64 V92 2.3862609845744497e-19

R64_93 V64 V93 -3244.4367135488496
L64_93 V64 V93 5.2725380792308065e-11
C64_93 V64 V93 1.457920424730126e-20

R64_94 V64 V94 5620.8380141977
L64_94 V64 V94 -5.377608145744143e-12
C64_94 V64 V94 -6.945099216161254e-20

R64_95 V64 V95 6854.00874283206
L64_95 V64 V95 -9.505475340802494e-11
C64_95 V64 V95 6.488482189148283e-21

R64_96 V64 V96 3371.267816425189
L64_96 V64 V96 1.5462952522154852e-11
C64_96 V64 V96 1.0756047159535993e-19

R64_97 V64 V97 7002.49406863562
L64_97 V64 V97 -4.4142048603161926e-12
C64_97 V64 V97 -1.7476001936514983e-20

R64_98 V64 V98 -4052.184461329686
L64_98 V64 V98 -2.707262347484706e-11
C64_98 V64 V98 -1.724068714017224e-21

R64_99 V64 V99 1608.9475254910817
L64_99 V64 V99 2.820817118608163e-12
C64_99 V64 V99 6.738299952667762e-20

R64_100 V64 V100 615.1005148458627
L64_100 V64 V100 -2.355154304124838e-12
C64_100 V64 V100 -4.0196202116225894e-19

R64_101 V64 V101 -13738.122665001976
L64_101 V64 V101 1.3209652214416784e-11
C64_101 V64 V101 1.70232928196749e-20

R64_102 V64 V102 10359.555532720307
L64_102 V64 V102 8.991204105229014e-12
C64_102 V64 V102 4.101663422331285e-20

R64_103 V64 V103 -2882.0566835542195
L64_103 V64 V103 -1.9633840733719948e-11
C64_103 V64 V103 1.4258739386186498e-20

R64_104 V64 V104 -934.2680801779102
L64_104 V64 V104 2.9360651284925767e-12
C64_104 V64 V104 2.4505023913731804e-19

R64_105 V64 V105 -7265.123366968732
L64_105 V64 V105 3.923590345822908e-12
C64_105 V64 V105 -2.744172724740203e-20

R64_106 V64 V106 7688.967966961046
L64_106 V64 V106 4.533596235728392e-11
C64_106 V64 V106 -5.569979621999095e-20

R64_107 V64 V107 -3020.1680693241274
L64_107 V64 V107 -3.925226550237356e-12
C64_107 V64 V107 -8.371322702749524e-20

R64_108 V64 V108 -1185.7556996376204
L64_108 V64 V108 2.7122308908399568e-12
C64_108 V64 V108 1.021209730806002e-19

R64_109 V64 V109 3316.037778284935
L64_109 V64 V109 -7.737229144495031e-12
C64_109 V64 V109 -1.6827035810765126e-20

R64_110 V64 V110 -177787.0689724696
L64_110 V64 V110 -1.0343495777075008e-11
C64_110 V64 V110 -1.9313637986783625e-20

R64_111 V64 V111 3066.2144593451826
L64_111 V64 V111 -2.387197998128406e-11
C64_111 V64 V111 -2.651720491297817e-20

R64_112 V64 V112 905.9798962764328
L64_112 V64 V112 -1.6759125808634243e-12
C64_112 V64 V112 -1.219732731334608e-19

R64_113 V64 V113 -1481.82515968006
L64_113 V64 V113 -4.042466795521915e-12
C64_113 V64 V113 2.3870697152960474e-20

R64_114 V64 V114 -29735.34774329552
L64_114 V64 V114 -6.248219065052297e-12
C64_114 V64 V114 1.6708160741180986e-20

R64_115 V64 V115 2506.5481650829106
L64_115 V64 V115 2.9435904378899307e-12
C64_115 V64 V115 1.0607269626699099e-19

R64_116 V64 V116 1035.8362465707726
L64_116 V64 V116 1.3913094052566988e-11
C64_116 V64 V116 -3.0224641748119275e-20

R64_117 V64 V117 2192.450713571945
L64_117 V64 V117 9.392719423164156e-12
C64_117 V64 V117 -1.8113275367867372e-20

R64_118 V64 V118 -19953.33767755275
L64_118 V64 V118 2.3266852403559583e-12
C64_118 V64 V118 6.102844032574323e-20

R64_119 V64 V119 -1372.1588518192025
L64_119 V64 V119 -8.294100712916541e-11
C64_119 V64 V119 -5.164382501433357e-20

R64_120 V64 V120 -435.50586647253465
L64_120 V64 V120 1.3727716277500368e-12
C64_120 V64 V120 -6.444226697803435e-20

R64_121 V64 V121 14466.507429878764
L64_121 V64 V121 3.0130735193957894e-12
C64_121 V64 V121 5.831348546919784e-20

R64_122 V64 V122 -12080.943577394723
L64_122 V64 V122 -4.653226816107027e-12
C64_122 V64 V122 -9.08946333405454e-20

R64_123 V64 V123 5732.453107884139
L64_123 V64 V123 -3.7604357244792806e-12
C64_123 V64 V123 -4.311778104553085e-20

R64_124 V64 V124 844.2238324076122
L64_124 V64 V124 -1.4942946316638225e-12
C64_124 V64 V124 2.297528002877612e-19

R64_125 V64 V125 -878.4706847456143
L64_125 V64 V125 1.548567875197312e-11
C64_125 V64 V125 -9.355919975656304e-21

R64_126 V64 V126 -3679.870489011637
L64_126 V64 V126 -2.5500187647162157e-12
C64_126 V64 V126 -5.210874093203113e-20

R64_127 V64 V127 3173.617108094366
L64_127 V64 V127 5.550364413138393e-11
C64_127 V64 V127 4.032285266309642e-20

R64_128 V64 V128 1120.139586622293
L64_128 V64 V128 -1.4470547524791028e-12
C64_128 V64 V128 -6.276030540173482e-20

R64_129 V64 V129 1067.0031104814686
L64_129 V64 V129 -1.6386839395044362e-12
C64_129 V64 V129 -1.1325916796523357e-19

R64_130 V64 V130 2374.193415222178
L64_130 V64 V130 2.6914245133196666e-12
C64_130 V64 V130 1.2618189455633655e-19

R64_131 V64 V131 -2454.2208853491725
L64_131 V64 V131 3.729934225522619e-12
C64_131 V64 V131 -4.537945559017651e-21

R64_132 V64 V132 -915.2759238324317
L64_132 V64 V132 7.707441079047382e-13
C64_132 V64 V132 -1.5183620550411802e-19

R64_133 V64 V133 3815.2967967234636
L64_133 V64 V133 2.976359244149256e-12
C64_133 V64 V133 7.808133084200021e-20

R64_134 V64 V134 -1131.1543073946377
L64_134 V64 V134 -1.526529725402977e-10
C64_134 V64 V134 -1.9341016513702788e-19

R64_135 V64 V135 -78249.34105725582
L64_135 V64 V135 -3.938726258617152e-11
C64_135 V64 V135 -6.890584917058953e-20

R64_136 V64 V136 1203.8734975014515
L64_136 V64 V136 7.723739914883571e-12
C64_136 V64 V136 2.512821733176962e-19

R64_137 V64 V137 -1021.2028048863257
L64_137 V64 V137 2.9943965966581167e-12
C64_137 V64 V137 1.1491806199552394e-19

R64_138 V64 V138 1951.0400025274757
L64_138 V64 V138 -3.23816236199303e-12
C64_138 V64 V138 1.1234846573079344e-19

R64_139 V64 V139 12811.341150905842
L64_139 V64 V139 -4.393399419619379e-12
C64_139 V64 V139 1.3743892660466617e-19

R64_140 V64 V140 -548.0860048229018
L64_140 V64 V140 -1.609389903474158e-12
C64_140 V64 V140 -2.1905439395838347e-19

R64_141 V64 V141 8189.637603618602
L64_141 V64 V141 -3.4169182944055923e-12
C64_141 V64 V141 -1.402276364390041e-19

R64_142 V64 V142 1073.7563669242754
L64_142 V64 V142 -5.631280657604459e-12
C64_142 V64 V142 7.610609663965414e-20

R64_143 V64 V143 182461.27848350196
L64_143 V64 V143 9.728996397835728e-12
C64_143 V64 V143 -6.862384202666024e-20

R64_144 V64 V144 804.5208678632647
L64_144 V64 V144 5.141696800915866e-11
C64_144 V64 V144 -1.8702316379173485e-20

R64_145 V64 V145 1043.779631809807
L64_145 V64 V145 -4.112188561041792e-12
C64_145 V64 V145 -8.896744519702166e-20

R64_146 V64 V146 -8531.787086921775
L64_146 V64 V146 1.6975365343134182e-12
C64_146 V64 V146 -9.011689297676568e-20

R64_147 V64 V147 1016.2169405377848
L64_147 V64 V147 -9.68232827195983e-11
C64_147 V64 V147 -4.83420876811532e-20

R64_148 V64 V148 4332.570277398767
L64_148 V64 V148 -1.9651832130553553e-11
C64_148 V64 V148 2.0283040392948738e-19

R64_149 V64 V149 -9638.171062930032
L64_149 V64 V149 2.240162294344563e-12
C64_149 V64 V149 2.4231864546877214e-19

R64_150 V64 V150 -653.4715152171041
L64_150 V64 V150 -6.560074721488977e-11
C64_150 V64 V150 -1.4905180216167633e-19

R64_151 V64 V151 -1173.3212620738868
L64_151 V64 V151 -4.485475943011212e-12
C64_151 V64 V151 6.714337922529624e-20

R64_152 V64 V152 318596.5352124488
L64_152 V64 V152 -8.867273237496454e-12
C64_152 V64 V152 -9.032705748117695e-20

R64_153 V64 V153 -895.4992250032872
L64_153 V64 V153 4.181567704031138e-12
C64_153 V64 V153 1.761252268053538e-20

R64_154 V64 V154 3530.2074426483573
L64_154 V64 V154 -4.8772989284304925e-12
C64_154 V64 V154 1.7294766570202973e-19

R64_155 V64 V155 752.9571261360185
L64_155 V64 V155 3.0215481027240603e-12
C64_155 V64 V155 5.822322350587567e-20

R64_156 V64 V156 -490.00515075992405
L64_156 V64 V156 1.1985140520802948e-12
C64_156 V64 V156 -9.120423474322338e-20

R64_157 V64 V157 -6253.896390912865
L64_157 V64 V157 -2.896212520982824e-12
C64_157 V64 V157 -1.7294252137258974e-19

R64_158 V64 V158 1899.3590310102052
L64_158 V64 V158 1.1322362595828731e-11
C64_158 V64 V158 -1.7372129543583454e-20

R64_159 V64 V159 -1185.7574376826117
L64_159 V64 V159 1.79243666600431e-12
C64_159 V64 V159 -3.075044862102407e-20

R64_160 V64 V160 672.7277635235483
L64_160 V64 V160 -2.7000498067541622e-12
C64_160 V64 V160 1.5860657258188286e-19

R64_161 V64 V161 2714.8698762974536
L64_161 V64 V161 -2.6145946618417185e-12
C64_161 V64 V161 -7.04773377154922e-20

R64_162 V64 V162 17177.467358958205
L64_162 V64 V162 5.688414269998791e-12
C64_162 V64 V162 -3.160703030018235e-20

R64_163 V64 V163 -3256.569165315933
L64_163 V64 V163 -1.9227177636391222e-12
C64_163 V64 V163 -4.273354941814408e-20

R64_164 V64 V164 -1655.7392876244917
L64_164 V64 V164 -8.007866949982407e-13
C64_164 V64 V164 -1.286658845124074e-19

R64_165 V64 V165 -3739.7623096960833
L64_165 V64 V165 2.3974022084554405e-12
C64_165 V64 V165 1.7274235339033275e-19

R64_166 V64 V166 -1059.5497368799827
L64_166 V64 V166 -2.670623635665684e-12
C64_166 V64 V166 3.1393835810510175e-20

R64_167 V64 V167 -9989.56643756113
L64_167 V64 V167 -2.279656342612533e-12
C64_167 V64 V167 -3.133620082977679e-20

R64_168 V64 V168 16249.275639481439
L64_168 V64 V168 6.197333137917841e-13
C64_168 V64 V168 -2.5703213629823597e-20

R64_169 V64 V169 -4238.68792003482
L64_169 V64 V169 3.395979225538265e-12
C64_169 V64 V169 5.787988285615759e-20

R64_170 V64 V170 1519.084589981939
L64_170 V64 V170 2.451106076560071e-12
C64_170 V64 V170 4.806495068281664e-20

R64_171 V64 V171 982.1896747910334
L64_171 V64 V171 1.4549616166633765e-12
C64_171 V64 V171 9.372792375140096e-20

R64_172 V64 V172 1731.1714668064055
L64_172 V64 V172 5.713529692396069e-12
C64_172 V64 V172 1.1401872827669966e-19

R64_173 V64 V173 5461.5004138406375
L64_173 V64 V173 -2.98936334210699e-12
C64_173 V64 V173 -1.0628072560969368e-19

R64_174 V64 V174 1666.4263930399468
L64_174 V64 V174 2.3374027185329744e-12
C64_174 V64 V174 -4.3651784945468974e-20

R64_175 V64 V175 -1674.3709855385766
L64_175 V64 V175 4.526022205264492e-12
C64_175 V64 V175 6.29325951927695e-20

R64_176 V64 V176 -24810.612004564115
L64_176 V64 V176 -6.810391294510255e-13
C64_176 V64 V176 -1.6616288580009908e-19

R64_177 V64 V177 -4621.634699245379
L64_177 V64 V177 -5.94998036916427e-12
C64_177 V64 V177 2.3149929544187e-20

R64_178 V64 V178 -1218.7144506807979
L64_178 V64 V178 -1.3565226848037904e-12
C64_178 V64 V178 -4.8601159699363366e-20

R64_179 V64 V179 14567.80823799306
L64_179 V64 V179 -1.6132977870230845e-12
C64_179 V64 V179 -1.2246372350590004e-19

R64_180 V64 V180 -911.2490220832428
L64_180 V64 V180 1.6595105489176683e-12
C64_180 V64 V180 8.077384152677046e-20

R64_181 V64 V181 14150.224410896184
L64_181 V64 V181 3.701829126689271e-12
C64_181 V64 V181 -1.4238519365828584e-20

R64_182 V64 V182 2493.1622516477114
L64_182 V64 V182 2.47186429960182e-12
C64_182 V64 V182 9.911113778904762e-20

R64_183 V64 V183 -3115.91304957606
L64_183 V64 V183 7.387847363142762e-11
C64_183 V64 V183 2.815007650274949e-20

R64_184 V64 V184 2961.200973983889
L64_184 V64 V184 8.94588706579904e-12
C64_184 V64 V184 -6.674352986542512e-20

R64_185 V64 V185 69113.23177094916
L64_185 V64 V185 2.3236143355550072e-11
C64_185 V64 V185 1.0951089984485992e-20

R64_186 V64 V186 3376.164432785245
L64_186 V64 V186 2.4395732515169726e-12
C64_186 V64 V186 -4.0839321187564305e-20

R64_187 V64 V187 10050.931012454785
L64_187 V64 V187 2.292700881620917e-12
C64_187 V64 V187 4.718728370238065e-20

R64_188 V64 V188 620.9028076109195
L64_188 V64 V188 -2.981823533138426e-12
C64_188 V64 V188 3.080133423451161e-20

R64_189 V64 V189 -7422.000682383784
L64_189 V64 V189 -6.298620953933995e-12
C64_189 V64 V189 7.846599095135914e-20

R64_190 V64 V190 -1721.3649536923847
L64_190 V64 V190 -3.4208201853372386e-12
C64_190 V64 V190 -7.817415306560439e-20

R64_191 V64 V191 4006.3431345610466
L64_191 V64 V191 4.9086154365760854e-11
C64_191 V64 V191 1.6749644104282786e-20

R64_192 V64 V192 -1021.4503610953851
L64_192 V64 V192 -8.696731117988026e-11
C64_192 V64 V192 1.547614641747358e-19

R64_193 V64 V193 5147.321066487674
L64_193 V64 V193 1.6188314267484132e-11
C64_193 V64 V193 -1.7521025070124405e-20

R64_194 V64 V194 -4516.6893822869715
L64_194 V64 V194 -3.5143995185538925e-11
C64_194 V64 V194 9.070587198433334e-20

R64_195 V64 V195 -2125.589261728432
L64_195 V64 V195 -4.600828567187171e-12
C64_195 V64 V195 2.6721090776675663e-20

R64_196 V64 V196 -1888.9546078547216
L64_196 V64 V196 -3.1268375047308032e-12
C64_196 V64 V196 -3.556055256685968e-19

R64_197 V64 V197 -19327.30916598071
L64_197 V64 V197 -1.0898603517362596e-11
C64_197 V64 V197 -1.1161508319961837e-19

R64_198 V64 V198 3865.6431364537884
L64_198 V64 V198 9.180228016299655e-12
C64_198 V64 V198 1.4479313718897156e-20

R64_199 V64 V199 -169397.57977495398
L64_199 V64 V199 -5.783690091615483e-12
C64_199 V64 V199 -1.0766780097258579e-19

R64_200 V64 V200 813.6235911062101
L64_200 V64 V200 3.446421864386154e-12
C64_200 V64 V200 6.975377775415261e-20

R65_65 V65 0 181.4218444430396
L65_65 V65 0 2.8230814574189815e-13
C65_65 V65 0 1.2447618722498356e-18

R65_66 V65 V66 77021.5879462157
L65_66 V65 V66 -3.5844490932632052e-12
C65_66 V65 V66 -1.2874015213284165e-19

R65_67 V65 V67 14321.97763652643
L65_67 V65 V67 -2.767067807774595e-12
C65_67 V65 V67 -1.3135444105819075e-19

R65_68 V65 V68 -125962.5489931745
L65_68 V65 V68 -1.838784148503935e-12
C65_68 V65 V68 -2.159553928623312e-19

R65_69 V65 V69 162758.6254598831
L65_69 V65 V69 1.7270221815224473e-12
C65_69 V65 V69 3.6572000568471933e-19

R65_70 V65 V70 24577.5883699817
L65_70 V65 V70 1.0817432754596488e-11
C65_70 V65 V70 8.866195836408627e-20

R65_71 V65 V71 -22457.907270670097
L65_71 V65 V71 -4.332673028906333e-12
C65_71 V65 V71 -1.7927291931593463e-19

R65_72 V65 V72 -51317.2221442674
L65_72 V65 V72 -5.078200466314354e-12
C65_72 V65 V72 -1.5696487978084921e-19

R65_73 V65 V73 -22838.699064627242
L65_73 V65 V73 3.694405240263999e-12
C65_73 V65 V73 1.7624468853333392e-19

R65_74 V65 V74 -21020.151432350576
L65_74 V65 V74 3.4031591471302654e-12
C65_74 V65 V74 1.4870655122706115e-19

R65_75 V65 V75 -5667.294744408043
L65_75 V65 V75 2.3962813743814676e-12
C65_75 V65 V75 2.2339621003956604e-19

R65_76 V65 V76 397528.21553205285
L65_76 V65 V76 1.4482092306917233e-12
C65_76 V65 V76 4.1125870133646035e-19

R65_77 V65 V77 6547.277406467606
L65_77 V65 V77 1.1053851089057586e-11
C65_77 V65 V77 -1.1170784551857008e-19

R65_78 V65 V78 -102732.20725366923
L65_78 V65 V78 -2.057355713511653e-11
C65_78 V65 V78 -5.993184170009937e-20

R65_79 V65 V79 4206.535683060626
L65_79 V65 V79 1.4002942985794872e-11
C65_79 V65 V79 1.1633233758703057e-20

R65_80 V65 V80 4010.150870527443
L65_80 V65 V80 -7.989720741988715e-12
C65_80 V65 V80 -1.2298217527601876e-19

R65_81 V65 V81 -914.9415174440416
L65_81 V65 V81 -1.7113906604443538e-12
C65_81 V65 V81 -1.705590781140496e-19

R65_82 V65 V82 6952.812980063795
L65_82 V65 V82 -3.242498704688418e-12
C65_82 V65 V82 -1.6242426990840327e-19

R65_83 V65 V83 3585.0725477900646
L65_83 V65 V83 -4.062969567334082e-12
C65_83 V65 V83 -1.3418693458429445e-19

R65_84 V65 V84 6204.459901333284
L65_84 V65 V84 -2.258387776729341e-12
C65_84 V65 V84 -2.39880257929797e-19

R65_85 V65 V85 -3614.5231949387257
L65_85 V65 V85 -6.582498514042623e-12
C65_85 V65 V85 -1.49539269182723e-19

R65_86 V65 V86 4237.3531844322515
L65_86 V65 V86 2.4246674350724835e-11
C65_86 V65 V86 -3.2338154921727604e-20

R65_87 V65 V87 -27693.124321966156
L65_87 V65 V87 4.0415564424482675e-12
C65_87 V65 V87 1.3149974149512655e-19

R65_88 V65 V88 -12362.443837501769
L65_88 V65 V88 2.6477838719559916e-12
C65_88 V65 V88 2.188417102173932e-19

R65_89 V65 V89 -5007.665311623095
L65_89 V65 V89 -7.084009510822406e-12
C65_89 V65 V89 1.3463186610751405e-19

R65_90 V65 V90 -6114.449299693582
L65_90 V65 V90 2.4797900231357174e-12
C65_90 V65 V90 3.078300989420543e-19

R65_91 V65 V91 -12468.667437992315
L65_91 V65 V91 -2.58549462809537e-12
C65_91 V65 V91 -2.2170147681543065e-19

R65_92 V65 V92 3573.4970845877015
L65_92 V65 V92 -4.022821224452523e-12
C65_92 V65 V92 -1.452659977346237e-19

R65_93 V65 V93 -3660.502003552733
L65_93 V65 V93 4.851779106567522e-12
C65_93 V65 V93 8.655233336818863e-20

R65_94 V65 V94 -6620.234717469077
L65_94 V65 V94 -4.6313617665874726e-12
C65_94 V65 V94 -1.0215241676974726e-19

R65_95 V65 V95 -67660.15242702472
L65_95 V65 V95 -3.079168549906874e-11
C65_95 V65 V95 -1.399548848442757e-20

R65_96 V65 V96 -24910.522775112848
L65_96 V65 V96 -2.086532828691131e-11
C65_96 V65 V96 -4.043162187487993e-20

R65_97 V65 V97 -2709.712333092268
L65_97 V65 V97 -3.7044688114953746e-12
C65_97 V65 V97 -1.0988267046936788e-19

R65_98 V65 V98 2091.145072265554
L65_98 V65 V98 -3.773649223208759e-12
C65_98 V65 V98 -2.3495230244153786e-19

R65_99 V65 V99 1930.769430708528
L65_99 V65 V99 2.1207817889176515e-12
C65_99 V65 V99 2.740739459618773e-19

R65_100 V65 V100 3379.7625189457262
L65_100 V65 V100 2.867278625848287e-12
C65_100 V65 V100 2.3113422385462206e-19

R65_101 V65 V101 -15894.19976497641
L65_101 V65 V101 6.8821010747329274e-12
C65_101 V65 V101 -5.096148966604706e-21

R65_102 V65 V102 12766.71719413187
L65_102 V65 V102 1.9641069694862225e-12
C65_102 V65 V102 2.3719334128569767e-19

R65_103 V65 V103 -75968.34751841986
L65_103 V65 V103 2.086328858272677e-11
C65_103 V65 V103 -4.305997122182052e-20

R65_104 V65 V104 17019.20219097842
L65_104 V65 V104 1.1591315754773404e-10
C65_104 V65 V104 -9.890515115487263e-20

R65_105 V65 V105 -749.0313729757348
L65_105 V65 V105 -3.017719386723913e-12
C65_105 V65 V105 -4.434721809533248e-20

R65_106 V65 V106 21108.676779631718
L65_106 V65 V106 3.4219866002249213e-11
C65_106 V65 V106 8.158284864687418e-20

R65_107 V65 V107 -33800.57947667482
L65_107 V65 V107 -3.107805044412669e-12
C65_107 V65 V107 -1.9589226888035762e-19

R65_108 V65 V108 7074.504898878592
L65_108 V65 V108 -5.2473939095873765e-12
C65_108 V65 V108 -6.364801504830889e-20

R65_109 V65 V109 2786.3861647918884
L65_109 V65 V109 -4.674536688647466e-12
C65_109 V65 V109 -1.6427478240761616e-19

R65_110 V65 V110 57013.96155173688
L65_110 V65 V110 -3.420725884194278e-12
C65_110 V65 V110 -1.6921421557322187e-19

R65_111 V65 V111 -18784.398207364356
L65_111 V65 V111 -9.696802153905921e-12
C65_111 V65 V111 -9.105109581167808e-21

R65_112 V65 V112 -13205.765037813098
L65_112 V65 V112 -1.1423305072918657e-11
C65_112 V65 V112 -3.7234369368892566e-20

R65_113 V65 V113 -8045.345398961037
L65_113 V65 V113 1.5790493972212126e-11
C65_113 V65 V113 9.381845817858724e-20

R65_114 V65 V114 5899.31633424984
L65_114 V65 V114 3.180053726907787e-11
C65_114 V65 V114 -5.345273926508371e-20

R65_115 V65 V115 4391.430888455659
L65_115 V65 V115 2.6008636382068525e-12
C65_115 V65 V115 1.8371921704464437e-19

R65_116 V65 V116 -25656.802633009556
L65_116 V65 V116 2.702889568371748e-12
C65_116 V65 V116 1.2152785359393362e-19

R65_117 V65 V117 -2079.8194636602075
L65_117 V65 V117 2.8228634431633434e-11
C65_117 V65 V117 1.7471197670988686e-19

R65_118 V65 V118 -4015.966205694314
L65_118 V65 V118 5.646919309961401e-12
C65_118 V65 V118 1.7550775458435975e-19

R65_119 V65 V119 4883.995358629836
L65_119 V65 V119 -1.6816402822254045e-11
C65_119 V65 V119 2.1416413269336258e-20

R65_120 V65 V120 1735.5492947889138
L65_120 V65 V120 -3.896702214168346e-11
C65_120 V65 V120 9.712597057475683e-20

R65_121 V65 V121 -17086.525694031872
L65_121 V65 V121 -7.198017606873278e-12
C65_121 V65 V121 -2.420854838421799e-19

R65_122 V65 V122 3700.6709817538517
L65_122 V65 V122 4.533659912341429e-11
C65_122 V65 V122 -2.7275501129157836e-20

R65_123 V65 V123 -4005.028820144113
L65_123 V65 V123 -9.906244805998147e-12
C65_123 V65 V123 -9.160110558678862e-20

R65_124 V65 V124 -2082.256741128182
L65_124 V65 V124 -4.566973192392453e-12
C65_124 V65 V124 -2.459421200942337e-19

R65_125 V65 V125 -828.2765376107071
L65_125 V65 V125 -8.785460269289289e-12
C65_125 V65 V125 -4.126635719366785e-20

R65_126 V65 V126 9423.34503641878
L65_126 V65 V126 -4.2900521452646696e-12
C65_126 V65 V126 -1.66459606316894e-19

R65_127 V65 V127 28792.80871631048
L65_127 V65 V127 -2.083096308886383e-11
C65_127 V65 V127 -8.085940163136156e-20

R65_128 V65 V128 -4410.939123631936
L65_128 V65 V128 -1.9190624256879898e-11
C65_128 V65 V128 -5.313638672213784e-20

R65_129 V65 V129 1965.412962336236
L65_129 V65 V129 -4.835230907842186e-12
C65_129 V65 V129 -1.0869657560037577e-19

R65_130 V65 V130 -8986.743088765841
L65_130 V65 V130 6.1784110813252195e-12
C65_130 V65 V130 1.314600259461588e-19

R65_131 V65 V131 24669.169335285194
L65_131 V65 V131 2.6369237575807524e-11
C65_131 V65 V131 1.1139269048035227e-19

R65_132 V65 V132 1790.203017945262
L65_132 V65 V132 5.902050483594692e-12
C65_132 V65 V132 2.3515778823907175e-19

R65_133 V65 V133 1283.477221305846
L65_133 V65 V133 5.169195389646797e-12
C65_133 V65 V133 3.1244665222544396e-19

R65_134 V65 V134 2279.563374217802
L65_134 V65 V134 1.3858828329486895e-11
C65_134 V65 V134 3.8130566689333534e-20

R65_135 V65 V135 -6010.842590385137
L65_135 V65 V135 9.129182339710316e-12
C65_135 V65 V135 1.5767732191891737e-20

R65_136 V65 V136 -2271.7493627487042
L65_136 V65 V136 -1.655558541483307e-10
C65_136 V65 V136 -1.0603700485301795e-19

R65_137 V65 V137 -749.7491322536632
L65_137 V65 V137 2.0450215573548427e-12
C65_137 V65 V137 7.605678439663798e-20

R65_138 V65 V138 -1443.9556023566734
L65_138 V65 V138 -1.3391262730012656e-11
C65_138 V65 V138 -5.867989221271053e-20

R65_139 V65 V139 1957.2871089607186
L65_139 V65 V139 7.209174808589133e-12
C65_139 V65 V139 6.79116344564883e-20

R65_140 V65 V140 1719.4734079718369
L65_140 V65 V140 2.7216510894221763e-12
C65_140 V65 V140 1.9764388786904852e-19

R65_141 V65 V141 2093.8739443050886
L65_141 V65 V141 -1.7935904457153746e-12
C65_141 V65 V141 -4.080274447513354e-19

R65_142 V65 V142 1722.719190889628
L65_142 V65 V142 -1.1504174344938805e-11
C65_142 V65 V142 -4.834662680692143e-20

R65_143 V65 V143 25005.172958930787
L65_143 V65 V143 -5.019920352558615e-12
C65_143 V65 V143 -6.826530737310762e-20

R65_144 V65 V144 2842.006152675484
L65_144 V65 V144 -2.9954460006803006e-12
C65_144 V65 V144 -1.2691701298841734e-19

R65_145 V65 V145 -1256.039706499998
L65_145 V65 V145 -1.7198888178690868e-12
C65_145 V65 V145 -4.549327776368106e-20

R65_146 V65 V146 3072.2934363621025
L65_146 V65 V146 -7.203512857763777e-12
C65_146 V65 V146 6.836163861474127e-20

R65_147 V65 V147 -2439.878659691084
L65_147 V65 V147 -5.738047718216734e-12
C65_147 V65 V147 -1.5518002614960378e-19

R65_148 V65 V148 -940.5903532131151
L65_148 V65 V148 -3.309917973721975e-12
C65_148 V65 V148 -1.7909042850614884e-19

R65_149 V65 V149 462.17898837840704
L65_149 V65 V149 1.7661388457728568e-12
C65_149 V65 V149 2.79831849902497e-19

R65_150 V65 V150 -1111.6062797494758
L65_150 V65 V150 8.564262816533882e-12
C65_150 V65 V150 -1.885160595312794e-19

R65_151 V65 V151 -2973.158836169881
L65_151 V65 V151 6.907137565802936e-11
C65_151 V65 V151 4.30605046695997e-20

R65_152 V65 V152 2062.6655810337274
L65_152 V65 V152 2.9250060589458085e-12
C65_152 V65 V152 7.811041517499644e-20

R65_153 V65 V153 -570.6763934606905
L65_153 V65 V153 2.1863034358261512e-12
C65_153 V65 V153 8.717843196677947e-20

R65_154 V65 V154 5990.885856019045
L65_154 V65 V154 3.529512945865788e-12
C65_154 V65 V154 1.251980151170526e-19

R65_155 V65 V155 997.7406208000067
L65_155 V65 V155 3.589896680124765e-12
C65_155 V65 V155 1.093877964155068e-19

R65_156 V65 V156 20159.752616131413
L65_156 V65 V156 1.9500632711264598e-11
C65_156 V65 V156 1.634352143411011e-19

R65_157 V65 V157 -914.6545383671842
L65_157 V65 V157 -1.7449283315500698e-12
C65_157 V65 V157 -2.1262779260412664e-19

R65_158 V65 V158 3278.1563098801967
L65_158 V65 V158 -6.468332412566664e-12
C65_158 V65 V158 3.2041621346791986e-20

R65_159 V65 V159 -2123.7475194256917
L65_159 V65 V159 4.96954044178023e-11
C65_159 V65 V159 4.164376942688305e-20

R65_160 V65 V160 5405.465367009569
L65_160 V65 V160 -1.6466644162242747e-11
C65_160 V65 V160 4.331115392418155e-21

R65_161 V65 V161 -3040.192736615298
L65_161 V65 V161 1.980322028016742e-11
C65_161 V65 V161 -7.369820844787771e-20

R65_162 V65 V162 3286.362941840795
L65_162 V65 V162 1.969545178929685e-11
C65_162 V65 V162 9.085852113553327e-20

R65_163 V65 V163 1552.0975227695974
L65_163 V65 V163 4.4214986290893484e-12
C65_163 V65 V163 1.2905614177552653e-20

R65_164 V65 V164 10095.819164465038
L65_164 V65 V164 6.850918174874416e-12
C65_164 V65 V164 2.1133986330710574e-20

R65_165 V65 V165 -2228.7767127362954
L65_165 V65 V165 -1.675167375343621e-12
C65_165 V65 V165 -3.7441469835010326e-21

R65_166 V65 V166 4773.828504881823
L65_166 V65 V166 7.893418583396998e-12
C65_166 V65 V166 -1.5424010319162377e-19

R65_167 V65 V167 -19631.08103197225
L65_167 V65 V167 -3.908744593704242e-12
C65_167 V65 V167 -8.264722219042475e-20

R65_168 V65 V168 1324.7538051007114
L65_168 V65 V168 -4.848372050686772e-12
C65_168 V65 V168 -1.519577100068305e-19

R65_169 V65 V169 -3568.9556005050836
L65_169 V65 V169 2.464141470891582e-12
C65_169 V65 V169 2.4901754760625963e-20

R65_170 V65 V170 -997.1400730589492
L65_170 V65 V170 -4.327455815888798e-12
C65_170 V65 V170 5.453137583066336e-20

R65_171 V65 V171 -1282.294838344604
L65_171 V65 V171 -1.0143377232584925e-11
C65_171 V65 V171 1.3751889837542676e-20

R65_172 V65 V172 -1580.798847174206
L65_172 V65 V172 -6.3023023307435815e-12
C65_172 V65 V172 6.082070975847682e-20

R65_173 V65 V173 -1112.623295159248
L65_173 V65 V173 2.836844359503299e-12
C65_173 V65 V173 1.0097062089415568e-19

R65_174 V65 V174 1040.6696422383152
L65_174 V65 V174 1.6025579908981336e-11
C65_174 V65 V174 6.886632342381818e-20

R65_175 V65 V175 1330.0563194792244
L65_175 V65 V175 2.4665859514999676e-12
C65_175 V65 V175 1.7343868625659316e-19

R65_176 V65 V176 2137.07094328044
L65_176 V65 V176 1.7563773536274658e-12
C65_176 V65 V176 2.5272325671151883e-19

R65_177 V65 V177 1829.5075185881783
L65_177 V65 V177 -1.1407076850346225e-12
C65_177 V65 V177 -1.2104146381450785e-19

R65_178 V65 V178 -3338.156089605531
L65_178 V65 V178 4.408606197984118e-12
C65_178 V65 V178 -4.7727099778526276e-20

R65_179 V65 V179 20894.59770169482
L65_179 V65 V179 -5.133697833904429e-12
C65_179 V65 V179 -1.36674711502913e-19

R65_180 V65 V180 -7935.349635444602
L65_180 V65 V180 -3.9751284632973324e-12
C65_180 V65 V180 -1.8792771645213124e-19

R65_181 V65 V181 2243.228810873971
L65_181 V65 V181 1.5169856020865982e-11
C65_181 V65 V181 -1.5977405078096614e-19

R65_182 V65 V182 -2478.9849167517505
L65_182 V65 V182 -2.8328713355281124e-11
C65_182 V65 V182 3.832053582924471e-20

R65_183 V65 V183 -3255.090529114735
L65_183 V65 V183 -4.197837051593573e-12
C65_183 V65 V183 -4.50360795756613e-20

R65_184 V65 V184 -6272.017802073064
L65_184 V65 V184 -3.358740721719599e-12
C65_184 V65 V184 -2.9623924451960396e-20

R65_185 V65 V185 -509.7024448746084
L65_185 V65 V185 1.6518734914332492e-12
C65_185 V65 V185 2.1016202643410745e-19

R65_186 V65 V186 873.2376153254202
L65_186 V65 V186 -2.1418034628712114e-12
C65_186 V65 V186 -1.238344684069517e-19

R65_187 V65 V187 2888.6742609100784
L65_187 V65 V187 1.2007692596426599e-11
C65_187 V65 V187 1.2050901304442023e-19

R65_188 V65 V188 6013.753562377988
L65_188 V65 V188 4.1047096892844095e-12
C65_188 V65 V188 6.957776853940983e-20

R65_189 V65 V189 467.98591059340373
L65_189 V65 V189 2.9459311945523065e-12
C65_189 V65 V189 5.0432545174428986e-20

R65_190 V65 V190 -3650.8731593239486
L65_190 V65 V190 5.7464440474202064e-12
C65_190 V65 V190 -4.0359013879916e-20

R65_191 V65 V191 -1346.9225671628856
L65_191 V65 V191 2.6713450882242e-12
C65_191 V65 V191 1.4313574850725304e-20

R65_192 V65 V192 -2102.4051631914176
L65_192 V65 V192 3.892782422873576e-12
C65_192 V65 V192 2.8600593610313575e-20

R65_193 V65 V193 2073.0483306460906
L65_193 V65 V193 -2.4304011516659673e-12
C65_193 V65 V193 -1.9696076842722062e-20

R65_194 V65 V194 -903.1981826122944
L65_194 V65 V194 2.1911569242558e-12
C65_194 V65 V194 2.7344799493809115e-20

R65_195 V65 V195 -19467.114405239845
L65_195 V65 V195 -3.681633360643596e-12
C65_195 V65 V195 -1.1535099172017845e-19

R65_196 V65 V196 -5440.77873942538
L65_196 V65 V196 -4.4147748044836546e-11
C65_196 V65 V196 5.2910541158352065e-20

R65_197 V65 V197 -608.7570578205728
L65_197 V65 V197 -3.153365727158925e-12
C65_197 V65 V197 -1.6480462767889904e-19

R65_198 V65 V198 1333.394619310764
L65_198 V65 V198 -3.030270507332275e-12
C65_198 V65 V198 -3.66497569269638e-20

R65_199 V65 V199 904.1961566775299
L65_199 V65 V199 -2.6539819639689535e-12
C65_199 V65 V199 2.0470111639985443e-20

R65_200 V65 V200 968.7009811347235
L65_200 V65 V200 -1.9838206995154946e-12
C65_200 V65 V200 -6.166738261412723e-20

R66_66 V66 0 -2246.2051934010055
L66_66 V66 0 6.035307717199742e-12
C66_66 V66 0 4.3099820402547124e-19

R66_67 V66 V67 -6424.459203222266
L66_67 V66 V67 -1.0976629440935575e-11
C66_67 V66 V67 -3.510740809828735e-20

R66_68 V66 V68 -5344.736432801419
L66_68 V66 V68 -1.64034847939323e-11
C66_68 V66 V68 -5.0855073176713175e-20

R66_69 V66 V69 -35427.68996216859
L66_69 V66 V69 5.110972293795243e-12
C66_69 V66 V69 1.617154110080251e-19

R66_70 V66 V70 2570.2267850605217
L66_70 V66 V70 3.3344664003327338e-12
C66_70 V66 V70 1.7504191330253972e-19

R66_71 V66 V71 11788.683079309485
L66_71 V66 V71 6.573887754291524e-11
C66_71 V66 V71 -3.8833968380144405e-20

R66_72 V66 V72 6247.566661552511
L66_72 V66 V72 -1.2922371160370915e-11
C66_72 V66 V72 -8.044663893368725e-20

R66_73 V66 V73 13728.098298647807
L66_73 V66 V73 5.749979847869153e-12
C66_73 V66 V73 1.0474448030723249e-19

R66_74 V66 V74 1071.336173235915
L66_74 V66 V74 1.3156620426220017e-12
C66_74 V66 V74 3.485942992035514e-19

R66_75 V66 V75 16620.87915177299
L66_75 V66 V75 1.7029857868168436e-11
C66_75 V66 V75 7.925597950579547e-20

R66_76 V66 V76 7501.398413259045
L66_76 V66 V76 1.2957290364268062e-11
C66_76 V66 V76 1.646082774028714e-19

R66_77 V66 V77 3203.1420023795686
L66_77 V66 V77 -4.628693610028228e-12
C66_77 V66 V77 -1.8044615533592422e-19

R66_78 V66 V78 -647.6268967523287
L66_78 V66 V78 -2.7320356142741247e-12
C66_78 V66 V78 -1.8479938019585637e-19

R66_79 V66 V79 -3873.539947913475
L66_79 V66 V79 -2.1531930025676182e-11
C66_79 V66 V79 -2.2322074869229917e-20

R66_80 V66 V80 -2180.2304848913545
L66_80 V66 V80 -2.796765574097164e-11
C66_80 V66 V80 -7.076178019042153e-20

R66_81 V66 V81 -1725.9837106515663
L66_81 V66 V81 -5.810872374734204e-12
C66_81 V66 V81 -3.073509578911698e-20

R66_82 V66 V82 1641.2888438672942
L66_82 V66 V82 -2.4663196209632032e-12
C66_82 V66 V82 -2.3323885950119392e-19

R66_83 V66 V83 5428.302418069095
L66_83 V66 V83 -1.1617975251629268e-11
C66_83 V66 V83 -6.630778408456008e-20

R66_84 V66 V84 16293.05105521252
L66_84 V66 V84 -9.068196664047453e-12
C66_84 V66 V84 -1.174211598404305e-19

R66_85 V66 V85 4619.665374469264
L66_85 V66 V85 4.445877166129293e-12
C66_85 V66 V85 9.04727800066532e-20

R66_86 V66 V86 1324.1995859058252
L66_86 V66 V86 9.344648131661679e-12
C66_86 V66 V86 9.538789623876358e-20

R66_87 V66 V87 4131.04636408161
L66_87 V66 V87 2.4871355398554354e-11
C66_87 V66 V87 1.8555288189539574e-20

R66_88 V66 V88 2357.7719314976516
L66_88 V66 V88 1.5132894534131954e-11
C66_88 V66 V88 7.528201706085017e-20

R66_89 V66 V89 3339.7745665753373
L66_89 V66 V89 -6.673820100473708e-12
C66_89 V66 V89 4.962915499673377e-21

R66_90 V66 V90 -916.8477172963425
L66_90 V66 V90 3.7902972258911394e-12
C66_90 V66 V90 2.353138830551811e-19

R66_91 V66 V91 -2082.062234127101
L66_91 V66 V91 1.0165634941073536e-11
C66_91 V66 V91 4.4049534579989905e-20

R66_92 V66 V92 -3703.038381643754
L66_92 V66 V92 7.48131994831632e-12
C66_92 V66 V92 2.9405829376606033e-20

R66_93 V66 V93 -3601.045444922046
L66_93 V66 V93 -7.169452881079209e-12
C66_93 V66 V93 -7.686896886457913e-20

R66_94 V66 V94 3444.9363897159315
L66_94 V66 V94 -4.697299467082767e-12
C66_94 V66 V94 -1.9804703037338779e-19

R66_95 V66 V95 -11135.327183570049
L66_95 V66 V95 -6.167710677426018e-12
C66_95 V66 V95 -4.388695703150838e-20

R66_96 V66 V96 -3589.291051882317
L66_96 V66 V96 -4.027778791776732e-12
C66_96 V66 V96 -6.678426749239846e-20

R66_97 V66 V97 3878.718660875361
L66_97 V66 V97 3.4484023527076497e-11
C66_97 V66 V97 -3.646363396333692e-21

R66_98 V66 V98 2312.4350046144036
L66_98 V66 V98 4.169212005949687e-12
C66_98 V66 V98 1.6612202628959787e-20

R66_99 V66 V99 2246.391312375218
L66_99 V66 V99 -1.1623251168573176e-11
C66_99 V66 V99 -2.4868503551178954e-20

R66_100 V66 V100 3417.277098101645
L66_100 V66 V100 6.117453614727462e-10
C66_100 V66 V100 -4.37228155967665e-21

R66_101 V66 V101 -1642.0096846826598
L66_101 V66 V101 9.59695737526476e-12
C66_101 V66 V101 6.57140941467295e-20

R66_102 V66 V102 -4129.368918815225
L66_102 V66 V102 -7.696459557130558e-11
C66_102 V66 V102 7.147952850112527e-20

R66_103 V66 V103 3695.7390778657514
L66_103 V66 V103 3.431180847114582e-12
C66_103 V66 V103 9.837718608486523e-20

R66_104 V66 V104 2565.47410795594
L66_104 V66 V104 3.024074735006052e-12
C66_104 V66 V104 7.607440975060686e-20

R66_105 V66 V105 1313.1966773009735
L66_105 V66 V105 -1.2031221170781355e-11
C66_105 V66 V105 -1.4679954374524102e-21

R66_106 V66 V106 -10078.95225430031
L66_106 V66 V106 -8.842697736459039e-12
C66_106 V66 V106 -8.168383098680732e-20

R66_107 V66 V107 -1476.9864227313371
L66_107 V66 V107 -7.947664985402062e-12
C66_107 V66 V107 -6.03722974716385e-20

R66_108 V66 V108 -2248.8658152084977
L66_108 V66 V108 -5.187018069858618e-12
C66_108 V66 V108 -3.17851339115938e-20

R66_109 V66 V109 2992.924332589202
L66_109 V66 V109 -1.5381797909949403e-11
C66_109 V66 V109 -8.368783542739477e-20

R66_110 V66 V110 -2267.74827881255
L66_110 V66 V110 4.78645210110316e-12
C66_110 V66 V110 6.912815551727832e-20

R66_111 V66 V111 -3417.2134808492397
L66_111 V66 V111 -1.290021309664509e-11
C66_111 V66 V111 -3.5556187290081473e-20

R66_112 V66 V112 -3421.9175950501844
L66_112 V66 V112 4.5607773298824985e-11
C66_112 V66 V112 -2.2331551042281534e-20

R66_113 V66 V113 -678.9589186851568
L66_113 V66 V113 -1.1715694823053064e-11
C66_113 V66 V113 -4.219416489880422e-20

R66_114 V66 V114 -12474.33055427741
L66_114 V66 V114 1.3005950809775751e-09
C66_114 V66 V114 -1.3733786888795535e-20

R66_115 V66 V115 1113.7355510415073
L66_115 V66 V115 1.751980319520063e-11
C66_115 V66 V115 4.257326070951238e-20

R66_116 V66 V116 1592.6881711364517
L66_116 V66 V116 1.8094597227122648e-11
C66_116 V66 V116 -2.682484189645572e-21

R66_117 V66 V117 4723.685655523626
L66_117 V66 V117 4.682393103845e-11
C66_117 V66 V117 1.1900982020029283e-19

R66_118 V66 V118 487.69163011927213
L66_118 V66 V118 1.2548402323262868e-11
C66_118 V66 V118 5.577916051046452e-21

R66_119 V66 V119 19126.310606625237
L66_119 V66 V119 -2.9012137736060982e-11
C66_119 V66 V119 -4.436806293545825e-21

R66_120 V66 V120 9814.890041725781
L66_120 V66 V120 -1.0989263730495725e-11
C66_120 V66 V120 1.0649627931533162e-20

R66_121 V66 V121 909.3095002718537
L66_121 V66 V121 8.781994462230255e-12
C66_121 V66 V121 -6.270576560698217e-21

R66_122 V66 V122 -739.3975377064476
L66_122 V66 V122 -9.565057694833962e-12
C66_122 V66 V122 -6.194067266509768e-20

R66_123 V66 V123 -1668.6522199340316
L66_123 V66 V123 4.47233101870492e-12
C66_123 V66 V123 6.559919860600387e-20

R66_124 V66 V124 -1480.1849506121412
L66_124 V66 V124 2.9411676866979167e-12
C66_124 V66 V124 6.108247609196436e-20

R66_125 V66 V125 21646.78480758983
L66_125 V66 V125 -4.078905928543297e-11
C66_125 V66 V125 -8.521451685503563e-20

R66_126 V66 V126 -422.29739768694924
L66_126 V66 V126 3.691933957491445e-12
C66_126 V66 V126 3.205215757652272e-20

R66_127 V66 V127 -2108.833062178421
L66_127 V66 V127 -1.0540979668878357e-11
C66_127 V66 V127 -7.764309067198593e-20

R66_128 V66 V128 -2388.2752325880065
L66_128 V66 V128 -7.125367451875425e-12
C66_128 V66 V128 -8.259045901157578e-20

R66_129 V66 V129 -721.1392682822835
L66_129 V66 V129 -4.9118586001442615e-12
C66_129 V66 V129 -6.740097807830045e-20

R66_130 V66 V130 407.9307871760776
L66_130 V66 V130 9.416038095802731e-12
C66_130 V66 V130 8.327595740647579e-20

R66_131 V66 V131 949.7812129428191
L66_131 V66 V131 -1.1838117355099247e-11
C66_131 V66 V131 -1.2369337634504713e-20

R66_132 V66 V132 685.0246290245528
L66_132 V66 V132 -7.031534227103432e-12
C66_132 V66 V132 4.8163854925806604e-21

R66_133 V66 V133 2496.6077919598542
L66_133 V66 V133 8.682553183041831e-12
C66_133 V66 V133 1.5801224593607468e-19

R66_134 V66 V134 4131.43050734997
L66_134 V66 V134 -2.3879785472665583e-12
C66_134 V66 V134 -1.289745240254061e-19

R66_135 V66 V135 3903.29761307651
L66_135 V66 V135 3.094137009861374e-12
C66_135 V66 V135 1.3841359687254188e-19

R66_136 V66 V136 2043.5972354880344
L66_136 V66 V136 3.10201830111347e-12
C66_136 V66 V136 6.988553614286597e-20

R66_137 V66 V137 1590.208846121897
L66_137 V66 V137 4.156002529991831e-12
C66_137 V66 V137 5.729410461807354e-20

R66_138 V66 V138 -621.8561492764004
L66_138 V66 V138 4.211740015819323e-12
C66_138 V66 V138 5.13506498911411e-20

R66_139 V66 V139 -844.6130975883017
L66_139 V66 V139 -5.651892930615025e-12
C66_139 V66 V139 -8.924993998375901e-20

R66_140 V66 V140 -474.6410416459916
L66_140 V66 V140 -2.258700428794301e-11
C66_140 V66 V140 -2.1885822997823167e-20

R66_141 V66 V141 1521.98353275695
L66_141 V66 V141 -1.60223688865255e-11
C66_141 V66 V141 -1.8719268381824295e-19

R66_142 V66 V142 1417.690881580762
L66_142 V66 V142 3.2616984689474537e-12
C66_142 V66 V142 5.421298351512246e-20

R66_143 V66 V143 3077.3010166095632
L66_143 V66 V143 -6.589472890763202e-12
C66_143 V66 V143 -5.624660214341513e-20

R66_144 V66 V144 1256.2850932294516
L66_144 V66 V144 -4.339223170846893e-12
C66_144 V66 V144 -3.855938962133104e-20

R66_145 V66 V145 -1157.46114290367
L66_145 V66 V145 -4.787074832894122e-12
C66_145 V66 V145 -2.3164459556920352e-20

R66_146 V66 V146 -944.5953018850424
L66_146 V66 V146 -4.0569813892119435e-12
C66_146 V66 V146 -2.1451537027236406e-20

R66_147 V66 V147 2867.4098974271956
L66_147 V66 V147 4.103284638567641e-12
C66_147 V66 V147 7.926757813760155e-20

R66_148 V66 V148 -2231.9623167591108
L66_148 V66 V148 3.822809771991035e-12
C66_148 V66 V148 -1.0190018340308363e-20

R66_149 V66 V149 -1121.960033946426
L66_149 V66 V149 4.3820054830551234e-11
C66_149 V66 V149 1.8544226071907623e-19

R66_150 V66 V150 333.6632442376525
L66_150 V66 V150 -3.951294605341021e-12
C66_150 V66 V150 -1.737764877113426e-19

R66_151 V66 V151 -3485.1757009770326
L66_151 V66 V151 4.1702529365061235e-12
C66_151 V66 V151 -1.608162110988527e-20

R66_152 V66 V152 2272.2493854751506
L66_152 V66 V152 5.0526919352374735e-12
C66_152 V66 V152 -1.30392588024423e-22

R66_153 V66 V153 1378.4150871542447
L66_153 V66 V153 7.620271641275195e-12
C66_153 V66 V153 2.499487056681559e-20

R66_154 V66 V154 -1117.3829705753199
L66_154 V66 V154 -1.0134026543614798e-11
C66_154 V66 V154 1.2802715646327546e-19

R66_155 V66 V155 2161.177801640317
L66_155 V66 V155 -4.78553754011188e-12
C66_155 V66 V155 3.737570571845303e-20

R66_156 V66 V156 -1236.270428888478
L66_156 V66 V156 -8.495982543606303e-12
C66_156 V66 V156 3.489502436340687e-20

R66_157 V66 V157 602.2137447527289
L66_157 V66 V157 -1.1433764511072559e-11
C66_157 V66 V157 -1.8276956476223459e-19

R66_158 V66 V158 -1743.9318558559053
L66_158 V66 V158 1.4293373404053218e-12
C66_158 V66 V158 -1.6032880587565065e-20

R66_159 V66 V159 -2667.9741818780635
L66_159 V66 V159 -3.994802499974103e-12
C66_159 V66 V159 3.878984965569701e-20

R66_160 V66 V160 1786.755911060095
L66_160 V66 V160 -2.461384449157667e-12
C66_160 V66 V160 5.005823350815665e-20

R66_161 V66 V161 -672.2929897461079
L66_161 V66 V161 -1.7984724884694534e-11
C66_161 V66 V161 -2.2160666716629366e-20

R66_162 V66 V162 -602.1857432871285
L66_162 V66 V162 -1.1387911369907751e-11
C66_162 V66 V162 -1.7485115008717868e-20

R66_163 V66 V163 -1230.6181636981548
L66_163 V66 V163 8.007741519414672e-12
C66_163 V66 V163 -7.960442008786256e-20

R66_164 V66 V164 -692.1505535833347
L66_164 V66 V164 3.502607097837443e-12
C66_164 V66 V164 -4.722278871913282e-20

R66_165 V66 V165 -1052.819019450392
L66_165 V66 V165 4.9631860007316085e-11
C66_165 V66 V165 9.320664656191608e-20

R66_166 V66 V166 800.2959789616599
L66_166 V66 V166 -1.3918589951264507e-12
C66_166 V66 V166 2.488683397222896e-20

R66_167 V66 V167 -2154.0644247594655
L66_167 V66 V167 3.6096653418527428e-12
C66_167 V66 V167 -4.090864601823129e-20

R66_168 V66 V168 -6280.502707343386
L66_168 V66 V168 5.2449053124428464e-12
C66_168 V66 V168 -5.798122145968283e-20

R66_169 V66 V169 460.4521591875134
L66_169 V66 V169 5.355890342964925e-11
C66_169 V66 V169 -1.497237470714934e-20

R66_170 V66 V170 490.4321991719752
L66_170 V66 V170 6.098057676200439e-12
C66_170 V66 V170 3.2803235444542394e-22

R66_171 V66 V171 753.6421839098463
L66_171 V66 V171 -4.878346419186802e-12
C66_171 V66 V171 1.1692060618464972e-19

R66_172 V66 V172 1097.1458256022333
L66_172 V66 V172 -5.59925421987389e-12
C66_172 V66 V172 9.07499159098499e-20

R66_173 V66 V173 -1034.1306539091388
L66_173 V66 V173 7.714152445610326e-11
C66_173 V66 V173 -2.488191078541921e-21

R66_174 V66 V174 -652.8595923436479
L66_174 V66 V174 1.430197702339538e-12
C66_174 V66 V174 -4.194120723697293e-20

R66_175 V66 V175 15971.06283895846
L66_175 V66 V175 -4.887505261345949e-12
C66_175 V66 V175 -1.606965119225868e-20

R66_176 V66 V176 -8763.069323597645
L66_176 V66 V176 -4.02985609834405e-12
C66_176 V66 V176 2.053249596059473e-20

R66_177 V66 V177 -583.4155989085132
L66_177 V66 V177 -9.335364319003598e-12
C66_177 V66 V177 1.664221751396937e-20

R66_178 V66 V178 -520.8345017511986
L66_178 V66 V178 -6.879980773537224e-12
C66_178 V66 V178 -2.329798116742972e-20

R66_179 V66 V179 -1784.2175509803503
L66_179 V66 V179 9.440586114342615e-12
C66_179 V66 V179 -5.999766325177347e-20

R66_180 V66 V180 -1106.0021309894464
L66_180 V66 V180 5.714553216592621e-12
C66_180 V66 V180 -6.064952976155886e-20

R66_181 V66 V181 714.7173470420545
L66_181 V66 V181 -3.815927184136576e-12
C66_181 V66 V181 -7.716420890230049e-20

R66_182 V66 V182 290.2232868557624
L66_182 V66 V182 -2.8462071418422138e-12
C66_182 V66 V182 7.593238352452508e-20

R66_183 V66 V183 -1893.9020688471894
L66_183 V66 V183 -2.4989861449723985e-11
C66_183 V66 V183 -2.810014850668525e-20

R66_184 V66 V184 -6109.738308836602
L66_184 V66 V184 1.949240052963632e-11
C66_184 V66 V184 4.837429691425058e-21

R66_185 V66 V185 1038.0120395565016
L66_185 V66 V185 3.3617851851042378e-12
C66_185 V66 V185 2.9200055356873934e-20

R66_186 V66 V186 1127.8235456429916
L66_186 V66 V186 7.998935417747403e-12
C66_186 V66 V186 2.50240612206053e-21

R66_187 V66 V187 3820.5635429189415
L66_187 V66 V187 -1.7277687292320507e-11
C66_187 V66 V187 4.041126103583266e-20

R66_188 V66 V188 1496.6666940508903
L66_188 V66 V188 -3.5645226822579224e-12
C66_188 V66 V188 1.0174521470090311e-20

R66_189 V66 V189 -694.3862589195406
L66_189 V66 V189 3.0026667828991927e-12
C66_189 V66 V189 1.2140174903712706e-19

R66_190 V66 V190 -436.4593212429696
L66_190 V66 V190 2.937335147912197e-12
C66_190 V66 V190 -9.651175721568229e-20

R66_191 V66 V191 2406.748768648775
L66_191 V66 V191 5.722801846490316e-12
C66_191 V66 V191 9.262997953996798e-20

R66_192 V66 V192 -4431.887210332914
L66_192 V66 V192 5.361160332597508e-12
C66_192 V66 V192 9.40154469674955e-20

R66_193 V66 V193 -3038.9658084895686
L66_193 V66 V193 -2.075144291737246e-12
C66_193 V66 V193 -5.263587970555773e-20

R66_194 V66 V194 635.8616702001339
L66_194 V66 V194 5.923152208286679e-12
C66_194 V66 V194 1.9480290861235665e-20

R66_195 V66 V195 -2759.805162507494
L66_195 V66 V195 -6.445474512716536e-12
C66_195 V66 V195 -1.564877774315e-19

R66_196 V66 V196 -1982.5895435166397
L66_196 V66 V196 -6.585311944404635e-12
C66_196 V66 V196 -1.306138090609164e-19

R66_197 V66 V197 1148.1800013262637
L66_197 V66 V197 -4.5671044876166e-12
C66_197 V66 V197 -1.0281308539321958e-19

R66_198 V66 V198 510.6475425689059
L66_198 V66 V198 -2.608615291711338e-12
C66_198 V66 V198 -3.7930390501148785e-21

R66_199 V66 V199 -69600.53624554319
L66_199 V66 V199 -2.4553485735605454e-12
C66_199 V66 V199 -8.903100258462789e-20

R66_200 V66 V200 -2524.3002416614854
L66_200 V66 V200 -3.1771922482657167e-12
C66_200 V66 V200 -3.0258820615055544e-20

R67_67 V67 0 -516.925632945206
L67_67 V67 0 3.368268182140376e-12
C67_67 V67 0 -7.94009558373896e-19

R67_68 V67 V68 -3433.4496581002195
L67_68 V67 V68 -5.010223706391831e-12
C67_68 V67 V68 -1.7832507961563558e-19

R67_69 V67 V69 -4213.010985608379
L67_69 V67 V69 7.803157344734655e-12
C67_69 V67 V69 9.6079087404608e-20

R67_70 V67 V70 7138.198138359881
L67_70 V67 V70 -1.1659752429163837e-11
C67_70 V67 V70 -6.886362214205644e-20

R67_71 V67 V71 3399.3118150649116
L67_71 V67 V71 2.355109532743534e-12
C67_71 V67 V71 2.3621085714309767e-19

R67_72 V67 V72 6334.597609275506
L67_72 V67 V72 4.008821996857162e-11
C67_72 V67 V72 -6.978992829709156e-21

R67_73 V67 V73 5198.556443859522
L67_73 V67 V73 5.2294536977415706e-12
C67_73 V67 V73 1.5632784539741305e-19

R67_74 V67 V74 4521.005999852605
L67_74 V67 V74 8.268585202711865e-12
C67_74 V67 V74 1.1017763611644134e-19

R67_75 V67 V75 1317.674214856262
L67_75 V67 V75 1.1789854427473814e-12
C67_75 V67 V75 4.436346562645177e-19

R67_76 V67 V76 7586.579033432668
L67_76 V67 V76 -3.330163927262659e-11
C67_76 V67 V76 1.0263378159576135e-19

R67_77 V67 V77 2219.0307986610715
L67_77 V67 V77 -1.0659649095327137e-11
C67_77 V67 V77 -6.344076241952452e-20

R67_78 V67 V78 -2280.353648248979
L67_78 V67 V78 -5.906364172304305e-11
C67_78 V67 V78 -3.056334669407083e-20

R67_79 V67 V79 -1453.9778864335221
L67_79 V67 V79 -2.512069598538279e-12
C67_79 V67 V79 -2.3289373099750246e-19

R67_80 V67 V80 -4421.840472563458
L67_80 V67 V80 6.047776279048641e-12
C67_80 V67 V80 4.1825066767610805e-21

R67_81 V67 V81 -2200.2832815628717
L67_81 V67 V81 -4.785150119993738e-12
C67_81 V67 V81 -2.6252480990397446e-20

R67_82 V67 V82 7274.407609628306
L67_82 V67 V82 -3.578531671911788e-11
C67_82 V67 V82 4.15208484846133e-20

R67_83 V67 V83 17842.50453985603
L67_83 V67 V83 -2.2660351470946722e-12
C67_83 V67 V83 -1.6251206328520825e-19

R67_84 V67 V84 -11721.377240491269
L67_84 V67 V84 -1.1096414380634297e-11
C67_84 V67 V84 -7.332842031409469e-20

R67_85 V67 V85 17440.5908091973
L67_85 V67 V85 5.68853049210888e-12
C67_85 V67 V85 6.692211234930501e-20

R67_86 V67 V86 1621.1318434556613
L67_86 V67 V86 2.1296783708207475e-11
C67_86 V67 V86 9.237822383194768e-21

R67_87 V67 V87 1489.1687921282594
L67_87 V67 V87 4.068194307486867e-12
C67_87 V67 V87 7.366176016225247e-20

R67_88 V67 V88 2644.8477176816073
L67_88 V67 V88 -6.543253543029259e-12
C67_88 V67 V88 -6.824796923919375e-20

R67_89 V67 V89 8685.078360801841
L67_89 V67 V89 -2.505321278118165e-12
C67_89 V67 V89 -1.4400692162785781e-19

R67_90 V67 V90 -1762.889645119756
L67_90 V67 V90 -5.384705418540552e-12
C67_90 V67 V90 -1.3362142429128348e-19

R67_91 V67 V91 -661.4981598544637
L67_91 V67 V91 -1.4124376016077337e-11
C67_91 V67 V91 6.938060806162657e-20

R67_92 V67 V92 -2961.053494405563
L67_92 V67 V92 2.7473649118087627e-12
C67_92 V67 V92 1.0466071340017313e-19

R67_93 V67 V93 18007.664990235124
L67_93 V67 V93 2.576895518280919e-10
C67_93 V67 V93 4.5140476318995285e-20

R67_94 V67 V94 -3582.604738290243
L67_94 V67 V94 8.94442551093713e-12
C67_94 V67 V94 1.106756635151349e-19

R67_95 V67 V95 15155.70959252199
L67_95 V67 V95 4.849632269645626e-12
C67_95 V67 V95 4.7322956349480717e-20

R67_96 V67 V96 -2916.8814984998057
L67_96 V67 V96 -7.872009679935692e-12
C67_96 V67 V96 6.364053422956603e-20

R67_97 V67 V97 4803.3143702021025
L67_97 V67 V97 5.216495541054381e-12
C67_97 V67 V97 2.08176174939981e-19

R67_98 V67 V98 2264.9697677781105
L67_98 V67 V98 1.3794927786446884e-11
C67_98 V67 V98 4.41746442625533e-20

R67_99 V67 V99 767.2122918406934
L67_99 V67 V99 9.509514931023671e-11
C67_99 V67 V99 -8.255183386181186e-20

R67_100 V67 V100 2465.8424901906733
L67_100 V67 V100 -9.345213754543718e-12
C67_100 V67 V100 -1.6139800598714333e-19

R67_101 V67 V101 -1309.6118256888465
L67_101 V67 V101 -2.1063366011269073e-11
C67_101 V67 V101 -1.1583923357777875e-19

R67_102 V67 V102 3272.9532150268396
L67_102 V67 V102 -3.060339545562668e-11
C67_102 V67 V102 -8.167069519945105e-20

R67_103 V67 V103 -19486.86568567739
L67_103 V67 V103 -2.1669645264566094e-12
C67_103 V67 V103 -1.1839217037706858e-19

R67_104 V67 V104 2195.148044908233
L67_104 V67 V104 3.992215376921774e-12
C67_104 V67 V104 4.2978003658585854e-20

R67_105 V67 V105 1321.113973334746
L67_105 V67 V105 -2.5818368184343533e-12
C67_105 V67 V105 -1.2505917470925336e-19

R67_106 V67 V106 -3130.2921111970973
L67_106 V67 V106 2.8721761411802094e-11
C67_106 V67 V106 -8.144057331422521e-21

R67_107 V67 V107 -718.9087448996111
L67_107 V67 V107 2.117500829120397e-12
C67_107 V67 V107 1.5067107132393492e-19

R67_108 V67 V108 -1555.7422050688865
L67_108 V67 V108 -4.7317196416847355e-12
C67_108 V67 V108 -1.8848078585887204e-21

R67_109 V67 V109 1481.7658192931963
L67_109 V67 V109 -1.7825100058271407e-11
C67_109 V67 V109 8.117467728348893e-20

R67_110 V67 V110 -2656.088903879872
L67_110 V67 V110 1.9788003959184372e-10
C67_110 V67 V110 4.99004174800518e-20

R67_111 V67 V111 -2685.400027859898
L67_111 V67 V111 5.5323807113062216e-11
C67_111 V67 V111 1.5382120351945135e-20

R67_112 V67 V112 -3203.5112327594543
L67_112 V67 V112 4.609505811872055e-12
C67_112 V67 V112 7.585443657749716e-20

R67_113 V67 V113 -659.3715392065166
L67_113 V67 V113 2.658252973411532e-12
C67_113 V67 V113 1.397862919394934e-19

R67_114 V67 V114 3752.5166681717055
L67_114 V67 V114 1.3004743044584219e-11
C67_114 V67 V114 2.9985241001266914e-20

R67_115 V67 V115 498.9064149468921
L67_115 V67 V115 -1.486890862232238e-11
C67_115 V67 V115 -8.514441911295222e-20

R67_116 V67 V116 1093.4592250193587
L67_116 V67 V116 -8.047348184724627e-12
C67_116 V67 V116 -4.727330829892847e-20

R67_117 V67 V117 -2332.725432550013
L67_117 V67 V117 -2.4784478531413067e-11
C67_117 V67 V117 6.915355873403737e-21

R67_118 V67 V118 1842.8518469995422
L67_118 V67 V118 -7.671776911600152e-12
C67_118 V67 V118 -1.0956929282026972e-19

R67_119 V67 V119 -963.7066738278461
L67_119 V67 V119 3.388542819285929e-11
C67_119 V67 V119 -3.5719876960733935e-20

R67_120 V67 V120 -4000.4938074260203
L67_120 V67 V120 -6.627549569434063e-12
C67_120 V67 V120 -1.0977774102362578e-19

R67_121 V67 V121 567.0692514457088
L67_121 V67 V121 -2.3501035188552422e-12
C67_121 V67 V121 -1.8040810417594793e-19

R67_122 V67 V122 -3087.741145735593
L67_122 V67 V122 5.840715182186359e-12
C67_122 V67 V122 1.0947125635290213e-19

R67_123 V67 V123 -1850.4456950330798
L67_123 V67 V123 -4.152650562358892e-12
C67_123 V67 V123 -1.0166692597129507e-20

R67_124 V67 V124 -1876.5336309723762
L67_124 V67 V124 1.7115257587390453e-12
C67_124 V67 V124 2.4105922541629646e-19

R67_125 V67 V125 2691.1805878327123
L67_125 V67 V125 -1.0353746043658771e-11
C67_125 V67 V125 -5.125811258195224e-20

R67_126 V67 V126 -961.8356508001175
L67_126 V67 V126 1.544662054737628e-11
C67_126 V67 V126 -1.759419598110159e-20

R67_127 V67 V127 -38180.72871770886
L67_127 V67 V127 1.8209731931021218e-12
C67_127 V67 V127 1.389045903649885e-19

R67_128 V67 V128 20371.267081404792
L67_128 V67 V128 -3.5249957330509905e-12
C67_128 V67 V128 -8.144669572034598e-20

R67_129 V67 V129 -514.2835525225976
L67_129 V67 V129 2.370730941945934e-12
C67_129 V67 V129 2.531332621420287e-19

R67_130 V67 V130 1218.568139932572
L67_130 V67 V130 -4.43853477628081e-12
C67_130 V67 V130 -1.1484018251859338e-19

R67_131 V67 V131 1566.928387746512
L67_131 V67 V131 -6.7335908131127585e-12
C67_131 V67 V131 -8.599688522566612e-20

R67_132 V67 V132 1994.211640921894
L67_132 V67 V132 -7.005986687152539e-12
C67_132 V67 V132 -9.120041493992284e-20

R67_133 V67 V133 197148.271778174
L67_133 V67 V133 -6.319734776519378e-12
C67_133 V67 V133 -8.255544384298181e-20

R67_134 V67 V134 2017.3819814956423
L67_134 V67 V134 4.426933661543547e-12
C67_134 V67 V134 1.9117032405299959e-19

R67_135 V67 V135 759.8062786683735
L67_135 V67 V135 -1.2200283198307004e-12
C67_135 V67 V135 -1.669744300681807e-19

R67_136 V67 V136 2383.856049977114
L67_136 V67 V136 2.505492921947351e-12
C67_136 V67 V136 2.23314647989016e-19

R67_137 V67 V137 533.1384558077735
L67_137 V67 V137 -3.740112428639344e-12
C67_137 V67 V137 -1.246555656610749e-19

R67_138 V67 V138 -1692.3584521869009
L67_138 V67 V138 -1.2973220262085544e-11
C67_138 V67 V138 -7.859256640502151e-20

R67_139 V67 V139 -474.16904346235486
L67_139 V67 V139 1.2021914109716341e-12
C67_139 V67 V139 1.7260413899885562e-19

R67_140 V67 V140 -1156.2592213363262
L67_140 V67 V140 -6.604336173408309e-12
C67_140 V67 V140 -1.8999788731291678e-19

R67_141 V67 V141 3069.0597969593687
L67_141 V67 V141 3.3602639538638333e-12
C67_141 V67 V141 1.5916356330779286e-19

R67_142 V67 V142 -1255.567504010774
L67_142 V67 V142 -1.2789882508600674e-11
C67_142 V67 V142 -8.899751123120482e-20

R67_143 V67 V143 -909.8428064624334
L67_143 V67 V143 1.6536849036692977e-12
C67_143 V67 V143 8.284711982082298e-20

R67_144 V67 V144 -1290.2386961606096
L67_144 V67 V144 -7.096162996783322e-12
C67_144 V67 V144 2.995390725434088e-20

R67_145 V67 V145 -442.7043517711487
L67_145 V67 V145 5.567490670473715e-12
C67_145 V67 V145 9.518978194764092e-20

R67_146 V67 V146 -10694.74860475302
L67_146 V67 V146 8.052464329085835e-12
C67_146 V67 V146 3.527566928656928e-20

R67_147 V67 V147 370.15153055545164
L67_147 V67 V147 -1.2826868245248912e-12
C67_147 V67 V147 -9.218196725746386e-20

R67_148 V67 V148 1127.0430773128514
L67_148 V67 V148 1.542247355130667e-12
C67_148 V67 V148 9.367090586305144e-20

R67_149 V67 V149 -2871.9046788610644
L67_149 V67 V149 -1.2709673260592232e-12
C67_149 V67 V149 -3.7917883305202856e-19

R67_150 V67 V150 525.67318038297
L67_150 V67 V150 -1.3668621189553405e-11
C67_150 V67 V150 2.3951384173030884e-19

R67_151 V67 V151 -1261.1992458644295
L67_151 V67 V151 -1.3940178409796842e-12
C67_151 V67 V151 -4.957804901130584e-20

R67_152 V67 V152 -2161.164883894781
L67_152 V67 V152 -2.933627394378968e-11
C67_152 V67 V152 -1.820557769534055e-20

R67_153 V67 V153 507.38277769195014
L67_153 V67 V153 -2.314642931429952e-11
C67_153 V67 V153 1.7347606140321224e-21

R67_154 V67 V154 7146.713722781865
L67_154 V67 V154 -1.0048650230113791e-11
C67_154 V67 V154 -1.6500616681001084e-19

R67_155 V67 V155 303.2294857463019
L67_155 V67 V155 1.7047785143445185e-12
C67_155 V67 V155 -4.726388255029161e-21

R67_156 V67 V156 1429.3549878738952
L67_156 V67 V156 -5.463595329614792e-12
C67_156 V67 V156 -1.02022514702722e-19

R67_157 V67 V157 510.51912870647374
L67_157 V67 V157 1.6235573757787826e-12
C67_157 V67 V157 4.551456063243379e-19

R67_158 V67 V158 -1017.0398829101372
L67_158 V67 V158 -3.281084628012057e-11
C67_158 V67 V158 -6.086389370282768e-21

R67_159 V67 V159 -371.2633595959704
L67_159 V67 V159 1.5439971446545657e-12
C67_159 V67 V159 -7.512358107356462e-20

R67_160 V67 V160 61580.394387350825
L67_160 V67 V160 -2.4576001678402215e-12
C67_160 V67 V160 3.2607817770607654e-20

R67_161 V67 V161 -512.1238877102732
L67_161 V67 V161 -3.1628411717629254e-10
C67_161 V67 V161 -4.0273781650912796e-20

R67_162 V67 V162 -1104.6295393240719
L67_162 V67 V162 -7.123485189177592e-12
C67_162 V67 V162 -5.1471607247119e-21

R67_163 V67 V163 -424.3279741056223
L67_163 V67 V163 -6.814098997659171e-12
C67_163 V67 V163 1.8112622698946472e-19

R67_164 V67 V164 -661.3252753813845
L67_164 V67 V164 2.4886867988450512e-12
C67_164 V67 V164 -1.861843895300542e-20

R67_165 V67 V165 -806.3870380273144
L67_165 V67 V165 -1.3107740200882074e-12
C67_165 V67 V165 -3.0899542088620705e-19

R67_166 V67 V166 795.0056745110529
L67_166 V67 V166 1.1633119200712566e-11
C67_166 V67 V166 2.0331492628082676e-20

R67_167 V67 V167 395.91716476196035
L67_167 V67 V167 -1.7409721707054912e-12
C67_167 V67 V167 -2.546764926938344e-20

R67_168 V67 V168 -2687.9613209053414
L67_168 V67 V168 1.9177703170981406e-11
C67_168 V67 V168 2.9535289317232084e-20

R67_169 V67 V169 607.3959709679461
L67_169 V67 V169 4.357513971199071e-12
C67_169 V67 V169 1.001503076487143e-19

R67_170 V67 V170 -2759.694812411804
L67_170 V67 V170 -8.176535126051533e-12
C67_170 V67 V170 -1.107044677193745e-19

R67_171 V67 V171 492.78569063036247
L67_171 V67 V171 -5.473987162839313e-12
C67_171 V67 V171 -2.2972483203676123e-19

R67_172 V67 V172 1070.9837889629578
L67_172 V67 V172 -6.041576751682408e-12
C67_172 V67 V172 -9.099084764285743e-20

R67_173 V67 V173 2717.570832403025
L67_173 V67 V173 2.5085514244752632e-12
C67_173 V67 V173 1.5498316161722185e-19

R67_174 V67 V174 -6903.511441341935
L67_174 V67 V174 -7.921288314746326e-12
C67_174 V67 V174 1.3718942483908199e-19

R67_175 V67 V175 -327.4286381055415
L67_175 V67 V175 1.383635405494411e-12
C67_175 V67 V175 9.590805462445956e-20

R67_176 V67 V176 22309.397662182913
L67_176 V67 V176 -8.566053430862426e-12
C67_176 V67 V176 -3.886381629110379e-20

R67_177 V67 V177 -654.2478231155304
L67_177 V67 V177 -2.2008876967825326e-12
C67_177 V67 V177 -9.572619979619974e-20

R67_178 V67 V178 53404.6240903496
L67_178 V67 V178 2.7497229866011037e-12
C67_178 V67 V178 8.057990509341885e-20

R67_179 V67 V179 1320.4299960112203
L67_179 V67 V179 -2.1011309325318787e-11
C67_179 V67 V179 1.4536853965824362e-19

R67_180 V67 V180 -2414.9882316119056
L67_180 V67 V180 3.0497027111852685e-12
C67_180 V67 V180 1.8278325894460638e-19

R67_181 V67 V181 1466.9928037574707
L67_181 V67 V181 -8.821850664852584e-12
C67_181 V67 V181 -5.3721916573968e-20

R67_182 V67 V182 1018.0185396881436
L67_182 V67 V182 -3.206418206025401e-12
C67_182 V67 V182 -1.4155176740733072e-19

R67_183 V67 V183 2094.9464365994845
L67_183 V67 V183 -3.990560440326993e-12
C67_183 V67 V183 5.353301384965562e-20

R67_184 V67 V184 -41400.18200414912
L67_184 V67 V184 4.8047268901695696e-11
C67_184 V67 V184 -4.648952881573613e-20

R67_185 V67 V185 817.1021557084063
L67_185 V67 V185 2.0383167143370892e-12
C67_185 V67 V185 7.472101794489143e-20

R67_186 V67 V186 -5448.749573017818
L67_186 V67 V186 -2.595936576615863e-12
C67_186 V67 V186 -6.260380757591485e-20

R67_187 V67 V187 -2011.5931563719532
L67_187 V67 V187 5.383442500556392e-12
C67_187 V67 V187 -9.35861671465695e-20

R67_188 V67 V188 4765.593154119224
L67_188 V67 V188 -1.4996617211739878e-12
C67_188 V67 V188 -1.405296897948016e-19

R67_189 V67 V189 -968.8911610321138
L67_189 V67 V189 8.84943070590691e-12
C67_189 V67 V189 -5.681455953462948e-20

R67_190 V67 V190 -3273.6062975955583
L67_190 V67 V190 4.405569411617981e-12
C67_190 V67 V190 1.5199791759065682e-19

R67_191 V67 V191 -7049.049500634026
L67_191 V67 V191 -2.1317749426131615e-11
C67_191 V67 V191 -1.8382075007573711e-19

R67_192 V67 V192 6525.733156703297
L67_192 V67 V192 2.136136117946151e-12
C67_192 V67 V192 3.1280933464591747e-20

R67_193 V67 V193 -1590.627904180012
L67_193 V67 V193 -2.4121171993172077e-12
C67_193 V67 V193 8.167815806182184e-20

R67_194 V67 V194 1009.2272459052721
L67_194 V67 V194 2.035541406888404e-12
C67_194 V67 V194 6.039974572116191e-20

R67_195 V67 V195 2702.676035056615
L67_195 V67 V195 3.018205760560104e-12
C67_195 V67 V195 3.0957954385858774e-19

R67_196 V67 V196 -1594.9545293628867
L67_196 V67 V196 8.389457361056328e-10
C67_196 V67 V196 3.3939101496005976e-20

R67_197 V67 V197 1960.397853036495
L67_197 V67 V197 5.921909571995263e-12
C67_197 V67 V197 1.6544116969789054e-21

R67_198 V67 V198 20469.46705063032
L67_198 V67 V198 -2.9538494936014778e-12
C67_198 V67 V198 -2.2675802080912182e-20

R67_199 V67 V199 1470.8415631958426
L67_199 V67 V199 -3.798671074996027e-12
C67_199 V67 V199 1.0119845814499073e-19

R67_200 V67 V200 -2096.079102250632
L67_200 V67 V200 -3.7772518332980494e-12
C67_200 V67 V200 4.1456553635849486e-20

R68_68 V68 0 -2339.4758312118297
L68_68 V68 0 3.210661316616695e-13
C68_68 V68 0 -2.8798761658369746e-19

R68_69 V68 V69 -5020.382267382123
L68_69 V68 V69 3.8253607280974095e-12
C68_69 V68 V69 1.918457695221578e-19

R68_70 V68 V70 6529.097785392049
L68_70 V68 V70 -1.8247062892617726e-11
C68_70 V68 V70 -4.999624007491484e-20

R68_71 V68 V71 8083.306363270861
L68_71 V68 V71 -1.3872625170138327e-11
C68_71 V68 V71 8.530288020473759e-21

R68_72 V68 V72 3665.3904828131376
L68_72 V68 V72 3.832848294586185e-12
C68_72 V68 V72 2.011612832383295e-19

R68_73 V68 V73 4869.7004854770985
L68_73 V68 V73 6.822931195054571e-12
C68_73 V68 V73 1.6934023680367305e-19

R68_74 V68 V74 2894.6307863039033
L68_74 V68 V74 7.024206969951925e-12
C68_74 V68 V74 1.5739199329736793e-19

R68_75 V68 V75 4760.163063991443
L68_75 V68 V75 2.8648547720745108e-12
C68_75 V68 V75 2.2102349848186757e-19

R68_76 V68 V76 803.6260089419364
L68_76 V68 V76 8.996314421212717e-13
C68_76 V68 V76 4.834125640552423e-19

R68_77 V68 V77 1653.8038590238818
L68_77 V68 V77 -1.5085686311551964e-10
C68_77 V68 V77 -3.689452061073865e-20

R68_78 V68 V78 -1424.0419067372284
L68_78 V68 V78 5.2204423132139685e-11
C68_78 V68 V78 -2.674798940559846e-20

R68_79 V68 V79 -5995.316939262768
L68_79 V68 V79 1.820088182139969e-11
C68_79 V68 V79 -3.046954254267139e-20

R68_80 V68 V80 -859.3735131694265
L68_80 V68 V80 -1.789721162945146e-12
C68_80 V68 V80 -2.7372644692285274e-19

R68_81 V68 V81 -1208.0709876365763
L68_81 V68 V81 -2.502566899256587e-12
C68_81 V68 V81 -1.2803969461249363e-19

R68_82 V68 V82 4225.690146910006
L68_82 V68 V82 -7.00616259080674e-12
C68_82 V68 V82 -3.033755242071615e-20

R68_83 V68 V83 -31589.237898881664
L68_83 V68 V83 -6.783395288482318e-12
C68_83 V68 V83 -1.2515582724238033e-19

R68_84 V68 V84 -6658.860524972363
L68_84 V68 V84 -2.4609041217739036e-12
C68_84 V68 V84 -1.223396772794784e-19

R68_85 V68 V85 17051.19137583762
L68_85 V68 V85 1.153837478654028e-11
C68_85 V68 V85 2.945002072629154e-20

R68_86 V68 V86 1339.685467832117
L68_86 V68 V86 7.715722356347228e-11
C68_86 V68 V86 -2.4035104511372848e-21

R68_87 V68 V87 2473.2103576382865
L68_87 V68 V87 8.94794951844915e-12
C68_87 V68 V87 8.0116572074302145e-22

R68_88 V68 V88 982.2460006678562
L68_88 V68 V88 3.0398388117574505e-12
C68_88 V68 V88 1.6652126709829762e-20

R68_89 V68 V89 3005.7936839734166
L68_89 V68 V89 -3.4485565877474567e-12
C68_89 V68 V89 -1.1431998846542595e-19

R68_90 V68 V90 -1668.3269297706881
L68_90 V68 V90 4.398554742569967e-12
C68_90 V68 V90 -1.7323973429603172e-20

R68_91 V68 V91 -1140.8904880517011
L68_91 V68 V91 -2.968135065282579e-11
C68_91 V68 V91 6.439688782787411e-20

R68_92 V68 V92 -602.76631647792
L68_92 V68 V92 -2.819456792931203e-12
C68_92 V68 V92 3.7112846279778146e-20

R68_93 V68 V93 -37881.51719003164
L68_93 V68 V93 1.1364388446651652e-11
C68_93 V68 V93 8.896840411319118e-20

R68_94 V68 V94 -4268.877307245752
L68_94 V68 V94 -3.964943427377059e-11
C68_94 V68 V94 4.888754286258548e-20

R68_95 V68 V95 -15363.578135633235
L68_95 V68 V95 -9.145099299754113e-11
C68_95 V68 V95 4.6312846906982557e-20

R68_96 V68 V96 4539.676991285214
L68_96 V68 V96 2.704719641145846e-12
C68_96 V68 V96 1.0507036352633628e-19

R68_97 V68 V97 3335.0241457894235
L68_97 V68 V97 -5.855736581761383e-11
C68_97 V68 V97 1.8846069350611726e-19

R68_98 V68 V98 3550.4173672743946
L68_98 V68 V98 -4.6931192926874e-12
C68_98 V68 V98 -2.5689636013926328e-20

R68_99 V68 V99 1331.3011198635388
L68_99 V68 V99 5.7835131845810485e-12
C68_99 V68 V99 -1.2535533720946633e-19

R68_100 V68 V100 875.5134043436144
L68_100 V68 V100 6.65513659864503e-12
C68_100 V68 V100 -1.8649670845200995e-20

R68_101 V68 V101 -1003.9838299603229
L68_101 V68 V101 1.2776253336179281e-11
C68_101 V68 V101 -1.6596757347852343e-19

R68_102 V68 V102 2377.4056923787975
L68_102 V68 V102 4.580126678204908e-12
C68_102 V68 V102 9.84945809935499e-21

R68_103 V68 V103 4183.744259305989
L68_103 V68 V103 1.0926110577759416e-11
C68_103 V68 V103 3.1395609194225976e-20

R68_104 V68 V104 4736.94124329621
L68_104 V68 V104 -2.1157778382874574e-12
C68_104 V68 V104 -1.205851477164588e-19

R68_105 V68 V105 1221.468018188017
L68_105 V68 V105 -2.2134127612224926e-12
C68_105 V68 V105 -1.3377479813181835e-19

R68_106 V68 V106 -2518.137545192809
L68_106 V68 V106 9.196835066493734e-12
C68_106 V68 V106 -2.3572836668514327e-20

R68_107 V68 V107 -1002.5086046276055
L68_107 V68 V107 -4.6535377063105165e-11
C68_107 V68 V107 5.523455350629547e-20

R68_108 V68 V108 -600.4975120352589
L68_108 V68 V108 2.6574857506111437e-12
C68_108 V68 V108 -1.4319582817737218e-20

R68_109 V68 V109 957.6579673811988
L68_109 V68 V109 -5.153804500319351e-12
C68_109 V68 V109 3.0091692025507646e-20

R68_110 V68 V110 -2605.85737500104
L68_110 V68 V110 -6.51896853526362e-11
C68_110 V68 V110 3.659938896984143e-20

R68_111 V68 V111 -1861.6987637883128
L68_111 V68 V111 -1.3263496457914783e-11
C68_111 V68 V111 -2.7289565654441796e-20

R68_112 V68 V112 -4275.010821326889
L68_112 V68 V112 -5.5235867431530206e-11
C68_112 V68 V112 8.719338868417343e-20

R68_113 V68 V113 -481.8011048993979
L68_113 V68 V113 2.4900200899258654e-12
C68_113 V68 V113 1.9874941825707485e-19

R68_114 V68 V114 2541.2468340610503
L68_114 V68 V114 -1.1203989314905904e-11
C68_114 V68 V114 2.3903558100287966e-20

R68_115 V68 V115 599.2072817832105
L68_115 V68 V115 -4.127238486437823e-11
C68_115 V68 V115 -3.3448140716999394e-20

R68_116 V68 V116 367.1076470595364
L68_116 V68 V116 6.46503385538456e-12
C68_116 V68 V116 2.8980128194967177e-20

R68_117 V68 V117 -3058.6533070705386
L68_117 V68 V117 6.339278352889439e-12
C68_117 V68 V117 8.915037336034675e-20

R68_118 V68 V118 1625.8879740585119
L68_118 V68 V118 -1.7236502503614147e-11
C68_118 V68 V118 -7.393493327572195e-20

R68_119 V68 V119 -1844.4201072841358
L68_119 V68 V119 1.4127342878932118e-10
C68_119 V68 V119 4.1062025803525274e-21

R68_120 V68 V120 -391.2733541941766
L68_120 V68 V120 5.787013686013046e-12
C68_120 V68 V120 -2.1178260400007193e-20

R68_121 V68 V121 478.65990031432136
L68_121 V68 V121 -1.7986332026125736e-12
C68_121 V68 V121 -3.1090615031044746e-19

R68_122 V68 V122 -1674.1412596034586
L68_122 V68 V122 4.5726832820899756e-12
C68_122 V68 V122 1.0433654551277208e-19

R68_123 V68 V123 -1215.034392313906
L68_123 V68 V123 4.699309271867201e-12
C68_123 V68 V123 1.1540121682180433e-19

R68_124 V68 V124 5929.390933501312
L68_124 V68 V124 -1.5947318726525609e-12
C68_124 V68 V124 -8.876115367681856e-20

R68_125 V68 V125 -9095.385662566836
L68_125 V68 V125 -3.1106084673629485e-12
C68_125 V68 V125 -9.782747162746687e-20

R68_126 V68 V126 -710.4437181697004
L68_126 V68 V126 -5.123387112413479e-12
C68_126 V68 V126 -7.131148646471867e-20

R68_127 V68 V127 7275.283160366381
L68_127 V68 V127 -3.949362810600556e-12
C68_127 V68 V127 -1.0843217935183714e-19

R68_128 V68 V128 1155.4704319699945
L68_128 V68 V128 3.0218961527050447e-12
C68_128 V68 V128 2.0980084798978446e-20

R68_129 V68 V129 -573.7565422904931
L68_129 V68 V129 2.2731323021929343e-12
C68_129 V68 V129 2.482434178830264e-19

R68_130 V68 V130 733.331915911578
L68_130 V68 V130 -1.7380971497049286e-11
C68_130 V68 V130 -3.980996641005224e-20

R68_131 V68 V131 3081.9345927202876
L68_131 V68 V131 1.8676716232345468e-11
C68_131 V68 V131 1.3144050721639848e-20

R68_132 V68 V132 -2981.847909224786
L68_132 V68 V132 5.560662464514643e-12
C68_132 V68 V132 5.604602531157776e-20

R68_133 V68 V133 212039.7462638036
L68_133 V68 V133 1.701029813508339e-11
C68_133 V68 V133 7.871276497512057e-20

R68_134 V68 V134 17579.980926382243
L68_134 V68 V134 3.783576577401429e-12
C68_134 V68 V134 2.2081998999392387e-19

R68_135 V68 V135 2490.9785272747945
L68_135 V68 V135 5.8150478628486675e-12
C68_135 V68 V135 1.4518181243213545e-19

R68_136 V68 V136 653.0049889201458
L68_136 V68 V136 -1.4009214644233848e-12
C68_136 V68 V136 -7.330082031600293e-20

R68_137 V68 V137 512.2965701936943
L68_137 V68 V137 -4.5312599265274784e-12
C68_137 V68 V137 -9.911262048944962e-20

R68_138 V68 V138 -2710.040068947611
L68_138 V68 V138 -3.918850041673881e-12
C68_138 V68 V138 -1.2160059819464154e-19

R68_139 V68 V139 -2156.86805898874
L68_139 V68 V139 -3.6912986760186025e-12
C68_139 V68 V139 -1.992625460705702e-19

R68_140 V68 V140 -398.0752624840982
L68_140 V68 V140 1.2571365134696472e-12
C68_140 V68 V140 1.3582357564393127e-19

R68_141 V68 V141 4320.559929435961
L68_141 V68 V141 -8.281845594861666e-12
C68_141 V68 V141 -5.602245943623979e-20

R68_142 V68 V142 -1838.3874835573004
L68_142 V68 V142 -2.8445556157658514e-11
C68_142 V68 V142 -9.961043314975863e-20

R68_143 V68 V143 -1268.3656323310145
L68_143 V68 V143 8.643744541918307e-12
C68_143 V68 V143 1.1228784864051245e-19

R68_144 V68 V144 -17575.16280368735
L68_144 V68 V144 3.009489400859559e-12
C68_144 V68 V144 -5.350704434238108e-20

R68_145 V68 V145 -435.80871422190785
L68_145 V68 V145 1.0400431859016264e-11
C68_145 V68 V145 7.631089227816461e-20

R68_146 V68 V146 -2756.035913349866
L68_146 V68 V146 3.20764029267617e-12
C68_146 V68 V146 7.485807583527085e-20

R68_147 V68 V147 1118.104758812665
L68_147 V68 V147 1.3359468867993312e-10
C68_147 V68 V147 1.5562808457812844e-20

R68_148 V68 V148 6380.1180317735825
L68_148 V68 V148 -9.459667825469552e-13
C68_148 V68 V148 -1.213048383381399e-19

R68_149 V68 V149 -1919.4583200869336
L68_149 V68 V149 -3.074893891683184e-12
C68_149 V68 V149 -2.8435999746064566e-19

R68_150 V68 V150 567.4630373833907
L68_150 V68 V150 -3.1700242207807055e-12
C68_150 V68 V150 1.184056207886361e-19

R68_151 V68 V151 23537.486021217694
L68_151 V68 V151 2.780431177931553e-11
C68_151 V68 V151 -1.1509328389148435e-19

R68_152 V68 V152 845.1310619881816
L68_152 V68 V152 -5.654202015154954e-12
C68_152 V68 V152 8.049254901612272e-20

R68_153 V68 V153 374.69650679479554
L68_153 V68 V153 5.042307166918271e-12
C68_153 V68 V153 1.4539708958572778e-19

R68_154 V68 V154 904.0704469725069
L68_154 V68 V154 1.1384250816703929e-11
C68_154 V68 V154 -8.752436767404223e-20

R68_155 V68 V155 555.811200823562
L68_155 V68 V155 -9.350310586024218e-12
C68_155 V68 V155 -6.991089673294491e-20

R68_156 V68 V156 -60062.60168216398
L68_156 V68 V156 2.6610631659409908e-12
C68_156 V68 V156 6.019785637996173e-20

R68_157 V68 V157 573.9980649087171
L68_157 V68 V157 2.036370394393874e-11
C68_157 V68 V157 3.289417273923536e-19

R68_158 V68 V158 -627.8599789236578
L68_158 V68 V158 -1.3044189783659221e-11
C68_158 V68 V158 -5.491890087384917e-21

R68_159 V68 V159 -1013.4146127756322
L68_159 V68 V159 -1.609124906796025e-11
C68_159 V68 V159 1.0973105759268463e-19

R68_160 V68 V160 -1193.6235111391948
L68_160 V68 V160 1.293700148179277e-12
C68_160 V68 V160 -7.994115481399593e-20

R68_161 V68 V161 -554.8748490918409
L68_161 V68 V161 9.795236297588766e-12
C68_161 V68 V161 -1.4271602372957436e-19

R68_162 V68 V162 -895.5036800470901
L68_162 V68 V162 1.4660191844926827e-11
C68_162 V68 V162 3.2099896574614363e-20

R68_163 V68 V163 -587.502053830581
L68_163 V68 V163 2.596887007935901e-12
C68_163 V68 V163 8.618277254231016e-20

R68_164 V68 V164 -243.6553448353813
L68_164 V68 V164 -2.225722764115151e-12
C68_164 V68 V164 6.853767149382694e-20

R68_165 V68 V165 -498.17114286945497
L68_165 V68 V165 -9.611855237477749e-13
C68_165 V68 V165 -3.0896085709741973e-19

R68_166 V68 V166 897.6542930273205
L68_166 V68 V166 -6.749018339664126e-12
C68_166 V68 V166 -6.779110842705178e-20

R68_167 V68 V167 -3869.788899081184
L68_167 V68 V167 -4.462577010201982e-11
C68_167 V68 V167 -6.889730007749545e-20

R68_168 V68 V168 238.43904966888928
L68_168 V68 V168 -2.4478851610312572e-12
C68_168 V68 V168 -8.23637857013832e-20

R68_169 V68 V169 487.637128840261
L68_169 V68 V169 2.299052165693676e-12
C68_169 V68 V169 1.620654398864748e-19

R68_170 V68 V170 3175.887445242732
L68_170 V68 V170 -3.529593156242613e-11
C68_170 V68 V170 -8.836529807664764e-20

R68_171 V68 V171 506.5688106527868
L68_171 V68 V171 -2.6400021323792593e-12
C68_171 V68 V171 -1.6969178957577251e-19

R68_172 V68 V172 812.2777536292255
L68_172 V68 V172 -6.305179224656862e-12
C68_172 V68 V172 -7.232613500647461e-20

R68_173 V68 V173 1592.344710873951
L68_173 V68 V173 1.7347632717669273e-12
C68_173 V68 V173 2.1367680365288438e-19

R68_174 V68 V174 -5174.798706928355
L68_174 V68 V174 1.3007584617877477e-11
C68_174 V68 V174 1.947967055255701e-19

R68_175 V68 V175 -1747.930898625232
L68_175 V68 V175 8.941364016901406e-12
C68_175 V68 V175 7.031189651748481e-20

R68_176 V68 V176 -328.6652846731548
L68_176 V68 V176 1.0272682374212853e-12
C68_176 V68 V176 2.1495116816085372e-19

R68_177 V68 V177 -499.9193496027358
L68_177 V68 V177 -1.3867100895584241e-12
C68_177 V68 V177 -1.5608235416745826e-19

R68_178 V68 V178 -1655.280581080951
L68_178 V68 V178 3.688211249762194e-12
C68_178 V68 V178 6.155567340093292e-20

R68_179 V68 V179 -4480.521231880925
L68_179 V68 V179 5.6538333947026504e-12
C68_179 V68 V179 1.6036846438793694e-19

R68_180 V68 V180 -1374.794481943283
L68_180 V68 V180 -4.402996027144705e-12
C68_180 V68 V180 -1.0550597127476068e-20

R68_181 V68 V181 1188.8186110828997
L68_181 V68 V181 -7.612724638455899e-12
C68_181 V68 V181 -1.7380914168005236e-19

R68_182 V68 V182 537.8972300991553
L68_182 V68 V182 -3.2413728271829886e-12
C68_182 V68 V182 -1.549126353636141e-19

R68_183 V68 V183 -2128.5431363606126
L68_183 V68 V183 -9.30867084875763e-12
C68_183 V68 V183 -1.4946875922182867e-20

R68_184 V68 V184 863.799781676404
L68_184 V68 V184 -1.7502531077518368e-12
C68_184 V68 V184 9.685305673643675e-21

R68_185 V68 V185 690.1497969643953
L68_185 V68 V185 1.9274590283443605e-12
C68_185 V68 V185 1.7504852252776975e-19

R68_186 V68 V186 -2938.576122551895
L68_186 V68 V186 -1.341547494237518e-12
C68_186 V68 V186 -9.985217708424558e-20

R68_187 V68 V187 -7284.708774185797
L68_187 V68 V187 -2.17587672221315e-12
C68_187 V68 V187 -1.271026667705734e-19

R68_188 V68 V188 657.8024457408719
L68_188 V68 V188 3.230882778350039e-12
C68_188 V68 V188 -1.468024854686351e-19

R68_189 V68 V189 -947.0850415888511
L68_189 V68 V189 4.437442478827098e-12
C68_189 V68 V189 1.2671781664974426e-22

R68_190 V68 V190 -1188.31870647497
L68_190 V68 V190 2.7619814190834868e-12
C68_190 V68 V190 1.313058110540733e-19

R68_191 V68 V191 938.8159409747844
L68_191 V68 V191 3.059673428705707e-12
C68_191 V68 V191 -3.228756657117578e-20

R68_192 V68 V192 -731.596598392
L68_192 V68 V192 8.576115656772235e-12
C68_192 V68 V192 1.3178646610381182e-20

R68_193 V68 V193 -1721.4255003058379
L68_193 V68 V193 -2.01234899353155e-12
C68_193 V68 V193 8.080545640757281e-20

R68_194 V68 V194 1073.6486506646838
L68_194 V68 V194 1.7462026157037382e-12
C68_194 V68 V194 8.475759593533157e-20

R68_195 V68 V195 -1433.59903605135
L68_195 V68 V195 -1.0952092058018557e-11
C68_195 V68 V195 4.627160529224604e-20

R68_196 V68 V196 -4216.647581802969
L68_196 V68 V196 1.830049909427879e-12
C68_196 V68 V196 2.577706602259403e-19

R68_197 V68 V197 1622.4354518639486
L68_197 V68 V197 2.806600186712542e-11
C68_197 V68 V197 -8.573436531225589e-20

R68_198 V68 V198 7168.126589594527
L68_198 V68 V198 -2.275705446784258e-12
C68_198 V68 V198 -3.6690798552090557e-20

R68_199 V68 V199 -923.2638688494458
L68_199 V68 V199 -4.257314413140239e-12
C68_199 V68 V199 1.3384103874175745e-19

R68_200 V68 V200 739.3920695248935
L68_200 V68 V200 -1.3566911011900104e-12
C68_200 V68 V200 -1.037363103723509e-19

R69_69 V69 0 374.8177622873291
L69_69 V69 0 -8.131013186816878e-13
C69_69 V69 0 -1.4822005577715989e-18

R69_70 V69 V70 2453.726580998882
L69_70 V69 V70 -2.360129058129252e-12
C69_70 V69 V70 -1.9089647866715955e-19

R69_71 V69 V71 1697.8991760131876
L69_71 V69 V71 -1.240748361348505e-11
C69_71 V69 V71 -3.4477250616346065e-20

R69_72 V69 V72 1615.102748010425
L69_72 V69 V72 -3.5441511869295898e-12
C69_72 V69 V72 -1.5758789504913208e-19

R69_73 V69 V73 712.4624019491933
L69_73 V69 V73 2.976423700254358e-12
C69_73 V69 V73 4.376229403144409e-19

R69_74 V69 V74 8458.942690048503
L69_74 V69 V74 -2.0882332901685175e-12
C69_74 V69 V74 -2.4055746789605264e-19

R69_75 V69 V75 18402.48923937858
L69_75 V69 V75 -4.1178378632622555e-12
C69_75 V69 V75 -1.0544323626954274e-19

R69_76 V69 V76 -6154.357352074232
L69_76 V69 V76 -1.6176006746730073e-12
C69_76 V69 V76 -3.5859647329265557e-19

R69_77 V69 V77 768.887575943769
L69_77 V69 V77 9.016658150266796e-13
C69_77 V69 V77 4.156999504747604e-19

R69_78 V69 V78 -997.0295879734216
L69_78 V69 V78 4.115732144330259e-12
C69_78 V69 V78 8.66822916441874e-20

R69_79 V69 V79 -905.488483223179
L69_79 V69 V79 6.322984554275118e-12
C69_79 V69 V79 4.591987913772619e-20

R69_80 V69 V80 -868.0566295736388
L69_80 V69 V80 1.4941221637587447e-12
C69_80 V69 V80 2.921957091947588e-19

R69_81 V69 V81 -272.90188868779563
L69_81 V69 V81 -4.0160793939077555e-12
C69_81 V69 V81 -1.575735928617597e-19

R69_82 V69 V82 1646.2039999350181
L69_82 V69 V82 1.6548314642927988e-12
C69_82 V69 V82 3.906573822262751e-19

R69_83 V69 V83 925.1440063845466
L69_83 V69 V83 4.768043434222738e-12
C69_83 V69 V83 1.1816239588857082e-19

R69_84 V69 V84 1039.6863027079487
L69_84 V69 V84 1.7767303525275619e-12
C69_84 V69 V84 2.6107925636443336e-19

R69_85 V69 V85 1063.7619989267398
L69_85 V69 V85 4.216561192066717e-12
C69_85 V69 V85 2.512562759640411e-19

R69_86 V69 V86 389.7424103409102
L69_86 V69 V86 -6.219054075552022e-12
C69_86 V69 V86 5.601947786161502e-22

R69_87 V69 V87 1290.4434397122297
L69_87 V69 V87 -2.3275945017786378e-12
C69_87 V69 V87 -2.4326589379377337e-19

R69_88 V69 V88 1009.504881647109
L69_88 V69 V88 -1.2330074698781988e-12
C69_88 V69 V88 -4.1256398249962905e-19

R69_89 V69 V89 517.2811048626677
L69_89 V69 V89 -9.331402962332216e-13
C69_89 V69 V89 -5.553173189531443e-19

R69_90 V69 V90 -435.99459877980365
L69_90 V69 V90 -8.741549862759904e-13
C69_90 V69 V90 -6.983277770842595e-19

R69_91 V69 V91 -570.3164997137014
L69_91 V69 V91 2.5415241494877145e-12
C69_91 V69 V91 2.7145702938994075e-19

R69_92 V69 V92 -667.475520052546
L69_92 V69 V92 2.6407515632140085e-12
C69_92 V69 V92 1.723970791547731e-19

R69_93 V69 V93 -281.1078330584684
L69_93 V69 V93 1.521541934288027e-11
C69_93 V69 V93 2.5557339284652083e-20

R69_94 V69 V94 -985.1243582555069
L69_94 V69 V94 1.7191338177977598e-12
C69_94 V69 V94 2.9691784422175995e-19

R69_95 V69 V95 -7670.652054178329
L69_95 V69 V95 3.1179524133453877e-12
C69_95 V69 V95 1.809131203850697e-19

R69_96 V69 V96 -1634.3170428240483
L69_96 V69 V96 2.732374195564085e-12
C69_96 V69 V96 2.524485539060899e-19

R69_97 V69 V97 2188.1336164374775
L69_97 V69 V97 6.589599958462457e-13
C69_97 V69 V97 8.71849308582265e-19

R69_98 V69 V98 366.0036482686589
L69_98 V69 V98 1.7719641477662761e-12
C69_98 V69 V98 4.797406408516265e-19

R69_99 V69 V99 574.223616064559
L69_99 V69 V99 -1.276027655154014e-12
C69_99 V69 V99 -4.980596580897191e-19

R69_100 V69 V100 565.4632633276402
L69_100 V69 V100 -3.3555089650573548e-12
C69_100 V69 V100 -3.516683799908826e-19

R69_101 V69 V101 434.5358115148873
L69_101 V69 V101 -1.0952950170694107e-12
C69_101 V69 V101 -5.883356743363883e-19

R69_102 V69 V102 -7139.428750646192
L69_102 V69 V102 -1.7245971350579909e-12
C69_102 V69 V102 -3.695105854523917e-19

R69_103 V69 V103 17590.894546049487
L69_103 V69 V103 2.1543239799368732e-11
C69_103 V69 V103 3.576354684294859e-20

R69_104 V69 V104 1934.3295776861905
L69_104 V69 V104 1.6027675825145132e-11
C69_104 V69 V104 4.6686596747261704e-20

R69_105 V69 V105 -236.57222938279247
L69_105 V69 V105 -1.5837123851683155e-12
C69_105 V69 V105 -8.097605036357543e-20

R69_106 V69 V106 -1773.2573858993094
L69_106 V69 V106 -3.0217963222193284e-12
C69_106 V69 V106 -3.052065318972071e-19

R69_107 V69 V107 -1886.3347344433546
L69_107 V69 V107 1.9447179376798712e-12
C69_107 V69 V107 3.3753084407715314e-19

R69_108 V69 V108 -1099.959761865374
L69_108 V69 V108 -5.535315255277609e-12
C69_108 V69 V108 3.169147356599658e-20

R69_109 V69 V109 1898.4880544494295
L69_109 V69 V109 1.2953958912741892e-12
C69_109 V69 V109 4.926435212909927e-19

R69_110 V69 V110 8106.3049458981095
L69_110 V69 V110 2.3233360885443287e-12
C69_110 V69 V110 3.267605147558703e-19

R69_111 V69 V111 -9040.045658844208
L69_111 V69 V111 -3.7061952788750183e-10
C69_111 V69 V111 -5.245692787450641e-20

R69_112 V69 V112 -93998.58693958503
L69_112 V69 V112 2.951164050642685e-12
C69_112 V69 V112 1.0732745800186226e-19

R69_113 V69 V113 567.3181766231019
L69_113 V69 V113 5.649973946808798e-10
C69_113 V69 V113 -2.2155517785351867e-19

R69_114 V69 V114 6518.10701737174
L69_114 V69 V114 2.055029715712381e-12
C69_114 V69 V114 2.9812162926903775e-19

R69_115 V69 V115 2919.5805378067357
L69_115 V69 V115 -2.072821229622326e-12
C69_115 V69 V115 -1.7629260399170466e-19

R69_116 V69 V116 1670.66767535195
L69_116 V69 V116 -6.1438984376375765e-12
C69_116 V69 V116 -1.7972040757092568e-20

R69_117 V69 V117 -369.6979999204464
L69_117 V69 V117 1.8762844095938174e-11
C69_117 V69 V117 3.3235345250026283e-20

R69_118 V69 V118 2481.5507461517936
L69_118 V69 V118 -1.3142992257663513e-12
C69_118 V69 V118 -4.633120120122717e-19

R69_119 V69 V119 3817.7782664455403
L69_119 V69 V119 -7.909148185457161e-12
C69_119 V69 V119 -9.720200998960658e-20

R69_120 V69 V120 3488.0182133392714
L69_120 V69 V120 -2.6759139229024165e-12
C69_120 V69 V120 -2.7707431572627314e-19

R69_121 V69 V121 -33942.80145659571
L69_121 V69 V121 -2.18354478779084e-12
C69_121 V69 V121 -6.169458735048635e-20

R69_122 V69 V122 -90244.6503718219
L69_122 V69 V122 4.844562875950935e-12
C69_122 V69 V122 7.85048967391856e-20

R69_123 V69 V123 -4246.215486626044
L69_123 V69 V123 1.8195948456413284e-12
C69_123 V69 V123 1.7991643669171625e-19

R69_124 V69 V124 -2565.1874263103973
L69_124 V69 V124 1.3472079415573775e-12
C69_124 V69 V124 3.570802387966664e-19

R69_125 V69 V125 1045.833025487337
L69_125 V69 V125 -4.030266915748925e-12
C69_125 V69 V125 -9.153422735000126e-20

R69_126 V69 V126 -3035.4882193290036
L69_126 V69 V126 1.9096890262681502e-12
C69_126 V69 V126 2.1614293408462007e-19

R69_127 V69 V127 -3987.1785515116185
L69_127 V69 V127 1.1492469340992725e-11
C69_127 V69 V127 1.166109752499525e-19

R69_128 V69 V128 -2752.748142623096
L69_128 V69 V128 -8.559603628580114e-12
C69_128 V69 V128 5.923355349872404e-20

R69_129 V69 V129 -637.3531305353674
L69_129 V69 V129 1.4827322637946118e-12
C69_129 V69 V129 5.2028221797885245e-19

R69_130 V69 V130 7526.947628140078
L69_130 V69 V130 -1.9999191319006332e-12
C69_130 V69 V130 -1.8830565811460215e-19

R69_131 V69 V131 1764.788191565265
L69_131 V69 V131 -2.518959047221744e-12
C69_131 V69 V131 -1.8753794257485023e-19

R69_132 V69 V132 1082.0361613211082
L69_132 V69 V132 -1.739717554195358e-12
C69_132 V69 V132 -3.285315777684255e-19

R69_133 V69 V133 -25598.66143015219
L69_133 V69 V133 -9.306919424025165e-12
C69_133 V69 V133 -5.18815045193069e-19

R69_134 V69 V134 1536.350280450596
L69_134 V69 V134 2.4483171027812645e-12
C69_134 V69 V134 9.502096694222592e-20

R69_135 V69 V135 -4392106.669402581
L69_135 V69 V135 6.3637012279172515e-12
C69_135 V69 V135 1.258132930833019e-20

R69_136 V69 V136 21293.302769592887
L69_136 V69 V136 2.348666687251219e-12
C69_136 V69 V136 2.702047607148215e-19

R69_137 V69 V137 1192.4061309710387
L69_137 V69 V137 -3.7927819332639784e-12
C69_137 V69 V137 -1.368911914521734e-19

R69_138 V69 V138 -1427.405705129075
L69_138 V69 V138 4.345979379267066e-11
C69_138 V69 V138 -6.74823488596318e-21

R69_139 V69 V139 -3047.188669903437
L69_139 V69 V139 -2.8659270917845415e-12
C69_139 V69 V139 -1.9240290766242758e-19

R69_140 V69 V140 -4187.6735461354265
L69_140 V69 V140 -4.889430676319242e-12
C69_140 V69 V140 -3.5819194333850024e-19

R69_141 V69 V141 3034.447624827594
L69_141 V69 V141 1.6497780322045847e-12
C69_141 V69 V141 6.7705477242030735e-19

R69_142 V69 V142 -2777.0435255961
L69_142 V69 V142 -3.673062919593094e-12
C69_142 V69 V142 -1.2227313622737285e-21

R69_143 V69 V143 7139.671393592862
L69_143 V69 V143 1.883358917696043e-12
C69_143 V69 V143 2.3448126178630187e-19

R69_144 V69 V144 -3930.021665317256
L69_144 V69 V144 1.3675156536024784e-11
C69_144 V69 V144 1.507523700869782e-19

R69_145 V69 V145 -374.2290923668163
L69_145 V69 V145 -3.501752842232646e-10
C69_145 V69 V145 -1.782751639348611e-20

R69_146 V69 V146 2605.6718253480967
L69_146 V69 V146 6.884727496426079e-12
C69_146 V69 V146 -1.9977097951656857e-20

R69_147 V69 V147 -11384.534382969048
L69_147 V69 V147 4.789650212405221e-12
C69_147 V69 V147 2.2257024870120904e-19

R69_148 V69 V148 4138.045646575997
L69_148 V69 V148 1.873153079091667e-12
C69_148 V69 V148 2.681019680306683e-19

R69_149 V69 V149 512.9552357747237
L69_149 V69 V149 -7.293640334696266e-13
C69_149 V69 V149 -7.426298348450356e-19

R69_150 V69 V150 764.031026469404
L69_150 V69 V150 7.585891130807508e-11
C69_150 V69 V150 3.763740081655503e-19

R69_151 V69 V151 -4273.576303039783
L69_151 V69 V151 -2.567810773767107e-12
C69_151 V69 V151 -2.352511176545988e-19

R69_152 V69 V152 22540.454898457203
L69_152 V69 V152 -3.195328131052505e-12
C69_152 V69 V152 -9.747262673415317e-20

R69_153 V69 V153 6048.487362345079
L69_153 V69 V153 9.908788334527355e-12
C69_153 V69 V153 5.1844035773613463e-20

R69_154 V69 V154 -14563.842642118581
L69_154 V69 V154 -1.1717963054466728e-11
C69_154 V69 V154 -2.727908038313911e-19

R69_155 V69 V155 2144.388410596232
L69_155 V69 V155 -1.3616428647690242e-12
C69_155 V69 V155 -1.99495872067485e-19

R69_156 V69 V156 1240.2986888422345
L69_156 V69 V156 -5.873638118959223e-12
C69_156 V69 V156 -2.5698719623308365e-19

R69_157 V69 V157 -906.1502491257664
L69_157 V69 V157 6.657280730478849e-13
C69_157 V69 V157 7.529211617233764e-19

R69_158 V69 V158 -1688.8500448062036
L69_158 V69 V158 -5.46841162075653e-12
C69_158 V69 V158 -8.029872459745781e-20

R69_159 V69 V159 2421.485454756045
L69_159 V69 V159 2.333466006546396e-12
C69_159 V69 V159 7.135589800273102e-20

R69_160 V69 V160 -2774.074520200608
L69_160 V69 V160 6.959380987730427e-12
C69_160 V69 V160 7.044686124038868e-20

R69_161 V69 V161 -990.3025790751302
L69_161 V69 V161 -2.052272307631009e-12
C69_161 V69 V161 -1.1352841778176206e-19

R69_162 V69 V162 -63149.10165355723
L69_162 V69 V162 -3.0221567269371542e-12
C69_162 V69 V162 -3.935852704498714e-20

R69_163 V69 V163 5444.6396555861775
L69_163 V69 V163 1.9032964788446516e-12
C69_163 V69 V163 1.4627447968407643e-19

R69_164 V69 V164 -26968.500695953488
L69_164 V69 V164 3.3432236454180297e-12
C69_164 V69 V164 -4.105348311230493e-20

R69_165 V69 V165 -717.2474910886045
L69_165 V69 V165 -1.7481863545739541e-12
C69_165 V69 V165 -2.8540771156594352e-19

R69_166 V69 V166 550.3506335728435
L69_166 V69 V166 1.1040456501521502e-11
C69_166 V69 V166 1.679292938202537e-19

R69_167 V69 V167 4918.259250062773
L69_167 V69 V167 -2.9519043044888067e-12
C69_167 V69 V167 -5.913686470496362e-20

R69_168 V69 V168 1704.7767486301416
L69_168 V69 V168 -1.956337358779556e-12
C69_168 V69 V168 7.221158267741836e-20

R69_169 V69 V169 1324.4374454655876
L69_169 V69 V169 -6.559008175045637e-11
C69_169 V69 V169 7.208459396172317e-20

R69_170 V69 V170 -689.8290823980738
L69_170 V69 V170 -2.8004690047718752e-12
C69_170 V69 V170 -2.7956107098503853e-19

R69_171 V69 V171 -1301.5708447113248
L69_171 V69 V171 -1.1129492176990401e-12
C69_171 V69 V171 -2.492869159743839e-19

R69_172 V69 V172 -1891.2059879665737
L69_172 V69 V172 -9.808828952799362e-12
C69_172 V69 V172 -1.4800339394197667e-19

R69_173 V69 V173 -3043.250914153936
L69_173 V69 V173 3.435765684324338e-12
C69_173 V69 V173 1.4797446386411648e-19

R69_174 V69 V174 -2333.828415485951
L69_174 V69 V174 1.7780033079445728e-12
C69_174 V69 V174 2.307138724769053e-19

R69_175 V69 V175 2149.466069789246
L69_175 V69 V175 2.8993173807922518e-12
C69_175 V69 V175 -7.86801673684988e-20

R69_176 V69 V176 3720.2043523650145
L69_176 V69 V176 3.845101481537985e-12
C69_176 V69 V176 -1.5703479540480495e-19

R69_177 V69 V177 -1129.435597991888
L69_177 V69 V177 1.4767841925963245e-12
C69_177 V69 V177 2.5737329723690637e-20

R69_178 V69 V178 1343.9895988100316
L69_178 V69 V178 4.9711172661230155e-12
C69_178 V69 V178 1.2867613236682474e-19

R69_179 V69 V179 2610.8542511399028
L69_179 V69 V179 1.8467181092356074e-12
C69_179 V69 V179 3.870436095770522e-19

R69_180 V69 V180 5943.0686581214895
L69_180 V69 V180 2.8954709812820948e-12
C69_180 V69 V180 3.730964811278958e-19

R69_181 V69 V181 820.7351770570978
L69_181 V69 V181 -1.2760182107195848e-12
C69_181 V69 V181 -1.239699171389052e-19

R69_182 V69 V182 9826.006294140743
L69_182 V69 V182 -1.1728938380513505e-12
C69_182 V69 V182 -2.2862181486982413e-19

R69_183 V69 V183 -4254.205024312784
L69_183 V69 V183 2.6320931790871735e-12
C69_183 V69 V183 5.322555246771056e-20

R69_184 V69 V184 -3453.6102308583477
L69_184 V69 V184 8.462817967638656e-12
C69_184 V69 V184 -5.426972343210331e-20

R69_185 V69 V185 -1712.8259498677946
L69_185 V69 V185 -1.5194379765480425e-12
C69_185 V69 V185 2.9415373149425947e-20

R69_186 V69 V186 -7586.479484581101
L69_186 V69 V186 3.37199232795418e-11
C69_186 V69 V186 2.072514827712165e-20

R69_187 V69 V187 -2473.5248015404463
L69_187 V69 V187 -1.5947142360062546e-12
C69_187 V69 V187 -3.302242032358613e-19

R69_188 V69 V188 -2315.217798016941
L69_188 V69 V188 -9.909739402801072e-13
C69_188 V69 V188 -2.5421488177215514e-19

R69_189 V69 V189 1324.465956678282
L69_189 V69 V189 1.2391990080851269e-12
C69_189 V69 V189 -4.6344363798287836e-20

R69_190 V69 V190 5595.440588721204
L69_190 V69 V190 3.0307953861631777e-12
C69_190 V69 V190 2.043883359878969e-19

R69_191 V69 V191 -4465.663621230121
L69_191 V69 V191 -1.08839839702768e-12
C69_191 V69 V191 -9.431453687321348e-20

R69_192 V69 V192 -11699.818175289543
L69_192 V69 V192 4.188952512652724e-11
C69_192 V69 V192 6.105456381868796e-20

R69_193 V69 V193 -27010.997664509858
L69_193 V69 V193 3.1674350098652492e-12
C69_193 V69 V193 7.748952206195721e-20

R69_194 V69 V194 25181.47143605577
L69_194 V69 V194 3.7353965544444164e-12
C69_194 V69 V194 1.41665600104141e-19

R69_195 V69 V195 3775.55377412729
L69_195 V69 V195 9.011326019361002e-13
C69_195 V69 V195 3.3419377712022016e-19

R69_196 V69 V196 4456.254291779253
L69_196 V69 V196 1.2933342815429859e-12
C69_196 V69 V196 8.288180745155808e-20

R69_197 V69 V197 -1161.4650896001149
L69_197 V69 V197 -7.840322599512083e-11
C69_197 V69 V197 8.395719302608782e-20

R69_198 V69 V198 2962.915079973006
L69_198 V69 V198 -7.645915709296268e-12
C69_198 V69 V198 -2.3597353329299528e-20

R69_199 V69 V199 1370.127409112235
L69_199 V69 V199 1.847802911482655e-12
C69_199 V69 V199 9.20505548167087e-20

R69_200 V69 V200 -128885.64679426969
L69_200 V69 V200 5.2164810026040584e-12
C69_200 V69 V200 9.608730051771842e-21

R70_70 V70 0 198.98991449465774
L70_70 V70 0 -1.2165841253456615e-12
C70_70 V70 0 -1.0940449900880029e-18

R70_71 V70 V71 -3951.946867572822
L70_71 V70 V71 4.572781376440267e-12
C70_71 V70 V71 2.0011633956496416e-19

R70_72 V70 V72 -2817.649905467564
L70_72 V70 V72 4.1600932800556485e-12
C70_72 V70 V72 2.576079450891819e-19

R70_73 V70 V73 -1611.0901253575757
L70_73 V70 V73 -5.676117026640492e-12
C70_73 V70 V73 -3.301574579144384e-20

R70_74 V70 V74 29687.42737578466
L70_74 V70 V74 1.7423920527230654e-12
C70_74 V70 V74 4.705402710238734e-19

R70_75 V70 V75 -8599.66688613398
L70_75 V70 V75 -6.783345186669097e-12
C70_75 V70 V75 -7.898917224331967e-20

R70_76 V70 V76 -21761.256884715807
L70_76 V70 V76 -1.9669082215539562e-12
C70_76 V70 V76 -3.7092388983608286e-19

R70_77 V70 V77 -3056.099844954883
L70_77 V70 V77 2.285414956064627e-12
C70_77 V70 V77 2.6806836766758283e-19

R70_78 V70 V78 437.0367802386965
L70_78 V70 V78 2.9530743981219407e-12
C70_78 V70 V78 7.617176956517613e-20

R70_79 V70 V79 1345.4996140684843
L70_79 V70 V79 -2.586456410367651e-11
C70_79 V70 V79 -7.522397182357136e-20

R70_80 V70 V80 1036.341877861742
L70_80 V70 V80 4.107559293370545e-12
C70_80 V70 V80 6.91388943433939e-20

R70_81 V70 V81 812.657839303374
L70_81 V70 V81 4.190600964572674e-11
C70_81 V70 V81 -1.2022352219471666e-20

R70_82 V70 V82 -716.2365174569665
L70_82 V70 V82 6.989779734949582e-11
C70_82 V70 V82 7.758407341870386e-20

R70_83 V70 V83 -1818.1885970334786
L70_83 V70 V83 6.510368681869878e-12
C70_83 V70 V83 1.4922273689098882e-19

R70_84 V70 V84 -1943.7348747973294
L70_84 V70 V84 2.573318070196493e-12
C70_84 V70 V84 2.655585815041581e-19

R70_85 V70 V85 -3403.124170628556
L70_85 V70 V85 -1.1258196508678318e-11
C70_85 V70 V85 -5.417955373309872e-20

R70_86 V70 V86 -333.1682082007151
L70_86 V70 V86 3.603555826722265e-12
C70_86 V70 V86 2.4975130409769776e-19

R70_87 V70 V87 -2484.386318496367
L70_87 V70 V87 -3.490316820477543e-12
C70_87 V70 V87 -1.7517661620450002e-19

R70_88 V70 V88 -1664.9763816488514
L70_88 V70 V88 -1.9261211798545398e-12
C70_88 V70 V88 -3.1152370873576823e-19

R70_89 V70 V89 -1474.8338922500818
L70_89 V70 V89 -2.066978576686222e-12
C70_89 V70 V89 -2.44124667727056e-19

R70_90 V70 V90 280.62110878573634
L70_90 V70 V90 -9.293393119252583e-13
C70_90 V70 V90 -7.921732337850751e-19

R70_91 V70 V91 1030.0698925678932
L70_91 V70 V91 3.020363211291956e-12
C70_91 V70 V91 1.601720128221394e-19

R70_92 V70 V92 1518.0991818072407
L70_92 V70 V92 3.636371179935048e-12
C70_92 V70 V92 1.0634635424323382e-19

R70_93 V70 V93 1147.5687479202631
L70_93 V70 V93 4.94750577688409e-12
C70_93 V70 V93 1.6112996009163766e-19

R70_94 V70 V94 4772.809533176521
L70_94 V70 V94 1.9994421286197818e-12
C70_94 V70 V94 3.834609877324246e-19

R70_95 V70 V95 -44372.67895944192
L70_95 V70 V95 2.929619669171185e-12
C70_95 V70 V95 2.3293618945183147e-19

R70_96 V70 V96 3778.8802910951513
L70_96 V70 V96 2.4367890789408436e-12
C70_96 V70 V96 2.973410859546841e-19

R70_97 V70 V97 3369.4541037165277
L70_97 V70 V97 1.6318652919590729e-12
C70_97 V70 V97 4.105990036405147e-19

R70_98 V70 V98 -427.7928566210115
L70_98 V70 V98 5.093767915142844e-12
C70_98 V70 V98 2.52074345297254e-19

R70_99 V70 V99 -3146.1329385515182
L70_99 V70 V99 -1.4593591118425587e-12
C70_99 V70 V99 -4.0822940200130534e-19

R70_100 V70 V100 -7783.62750444271
L70_100 V70 V100 -2.2320977717030246e-12
C70_100 V70 V100 -3.954272030799807e-19

R70_101 V70 V101 -32290.01112708009
L70_101 V70 V101 -2.3573322305976024e-12
C70_101 V70 V101 -3.2088048244345456e-19

R70_102 V70 V102 593.0619759991688
L70_102 V70 V102 -3.556471985268038e-12
C70_102 V70 V102 -2.6499122927799477e-19

R70_103 V70 V103 -1472.4130598377972
L70_103 V70 V103 1.9577416706225172e-10
C70_103 V70 V103 5.19635683426141e-21

R70_104 V70 V104 -1004.6427712274083
L70_104 V70 V104 8.09862272945551e-11
C70_104 V70 V104 3.8079456847106214e-20

R70_105 V70 V105 -1633.2272565327735
L70_105 V70 V105 -2.287782648973892e-12
C70_105 V70 V105 -1.6118430892995976e-19

R70_106 V70 V106 -352.013570749225
L70_106 V70 V106 -1.2700022382733678e-11
C70_106 V70 V106 4.124294499651442e-20

R70_107 V70 V107 1311.906299743181
L70_107 V70 V107 1.7845795768478932e-12
C70_107 V70 V107 3.0638497120792436e-19

R70_108 V70 V108 1999.6818527706134
L70_108 V70 V108 5.625636255274128e-12
C70_108 V70 V108 1.0126453288997884e-19

R70_109 V70 V109 1604.2282783334517
L70_109 V70 V109 2.6633582601444464e-12
C70_109 V70 V109 2.8662192078434326e-19

R70_110 V70 V110 386.18216936283113
L70_110 V70 V110 -9.473589844811133e-12
C70_110 V70 V110 -2.9879913007815543e-19

R70_111 V70 V111 6549.455749190841
L70_111 V70 V111 -1.077903579056239e-11
C70_111 V70 V111 -1.1232411384175096e-20

R70_112 V70 V112 2168.973610321643
L70_112 V70 V112 2.7867371659490695e-11
C70_112 V70 V112 9.307179816823125e-20

R70_113 V70 V113 642.5777766445659
L70_113 V70 V113 2.7006288914783503e-12
C70_113 V70 V113 1.447438612596615e-19

R70_114 V70 V114 439.61714105807005
L70_114 V70 V114 1.2770653526612673e-12
C70_114 V70 V114 5.140317664335031e-19

R70_115 V70 V115 -1821.048718461777
L70_115 V70 V115 -2.3030123834301168e-12
C70_115 V70 V115 -1.905231563813199e-19

R70_116 V70 V116 -2449.6636655828847
L70_116 V70 V116 -5.27723874862416e-12
C70_116 V70 V116 -2.112978768911015e-20

R70_117 V70 V117 -1387.8571301653064
L70_117 V70 V117 -4.479260821468389e-12
C70_117 V70 V117 -1.4335748283456325e-19

R70_118 V70 V118 -144.8280904822946
L70_118 V70 V118 -1.375797361034585e-12
C70_118 V70 V118 -2.986801427883222e-19

R70_119 V70 V119 -1512.9281305462566
L70_119 V70 V119 5.59033585125303e-12
C70_119 V70 V119 -7.575755800408416e-20

R70_120 V70 V120 -2015.6535334806363
L70_120 V70 V120 8.711733310007461e-12
C70_120 V70 V120 -2.506449480019954e-19

R70_121 V70 V121 -1112.4099230163295
L70_121 V70 V121 -2.9154911620950272e-12
C70_121 V70 V121 -8.242209963551048e-20

R70_122 V70 V122 459.2360340466101
L70_122 V70 V122 -1.228994648542136e-11
C70_122 V70 V122 -1.1643853912714594e-19

R70_123 V70 V123 6719.800541442369
L70_123 V70 V123 6.689657038136537e-12
C70_123 V70 V123 2.0025176879020756e-19

R70_124 V70 V124 4274.616264170709
L70_124 V70 V124 5.715993227621968e-12
C70_124 V70 V124 3.44338882599852e-19

R70_125 V70 V125 4400.01592765472
L70_125 V70 V125 1.2143383535593567e-11
C70_125 V70 V125 -2.469735748473624e-20

R70_126 V70 V126 170.1592919112122
L70_126 V70 V126 1.334069723636896e-12
C70_126 V70 V126 4.1792965694213716e-19

R70_127 V70 V127 503.9362030162714
L70_127 V70 V127 1.4711642049686104e-11
C70_127 V70 V127 6.59228304879678e-20

R70_128 V70 V128 606.6025746538857
L70_128 V70 V128 -9.025457160605552e-12
C70_128 V70 V128 6.793400253408956e-20

R70_129 V70 V129 548.1462069185665
L70_129 V70 V129 1.835033599267789e-12
C70_129 V70 V129 3.5212684483122023e-19

R70_130 V70 V130 -222.76705381769202
L70_130 V70 V130 -1.6835760597590122e-12
C70_130 V70 V130 -3.89365683432939e-19

R70_131 V70 V131 -383.03088634243267
L70_131 V70 V131 -6.065125389145221e-12
C70_131 V70 V131 -1.9103163176613262e-19

R70_132 V70 V132 -306.7691463845816
L70_132 V70 V132 -8.192265508754676e-12
C70_132 V70 V132 -3.7569534373812444e-19

R70_133 V70 V133 -1335.6317582502375
L70_133 V70 V133 -2.4795138785616515e-12
C70_133 V70 V133 -2.565939784052085e-19

R70_134 V70 V134 -551.2005139322599
L70_134 V70 V134 1.991420289500865e-12
C70_134 V70 V134 1.6195875976905163e-19

R70_135 V70 V135 -1154.291689638588
L70_135 V70 V135 -6.6237345510407236e-12
C70_135 V70 V135 3.7628344046508063e-20

R70_136 V70 V136 -618.6558244264112
L70_136 V70 V136 2.0822631994613364e-11
C70_136 V70 V136 2.785230951594936e-19

R70_137 V70 V137 -985.6931636916801
L70_137 V70 V137 -3.370414122968022e-12
C70_137 V70 V137 -1.6899322476133926e-19

R70_138 V70 V138 268.6002212978193
L70_138 V70 V138 -7.086254124880882e-11
C70_138 V70 V138 8.562801891745801e-20

R70_139 V70 V139 304.8013010863283
L70_139 V70 V139 8.524863028583904e-12
C70_139 V70 V139 -9.945626333623964e-20

R70_140 V70 V140 197.5900883675196
L70_140 V70 V140 5.871478444805967e-12
C70_140 V70 V140 -1.770132053707662e-19

R70_141 V70 V141 -942.3580762342067
L70_141 V70 V141 1.696668898242351e-12
C70_141 V70 V141 4.326763475179513e-19

R70_142 V70 V142 847.9884578897406
L70_142 V70 V142 -1.2777887257575945e-12
C70_142 V70 V142 -2.2490233952019197e-19

R70_143 V70 V143 -558.3415416412631
L70_143 V70 V143 3.505087682285493e-12
C70_143 V70 V143 1.6863438186746172e-19

R70_144 V70 V144 -530.4929498081217
L70_144 V70 V144 -2.6102506229471322e-11
C70_144 V70 V144 -3.3762788815221072e-21

R70_145 V70 V145 692.6542389772297
L70_145 V70 V145 5.64598251651933e-12
C70_145 V70 V145 9.206523728819427e-20

R70_146 V70 V146 -225.30095985462816
L70_146 V70 V146 1.5208851695204853e-12
C70_146 V70 V146 6.792791769778393e-20

R70_147 V70 V147 -2031.6883876234674
L70_147 V70 V147 -1.0661404407755985e-11
C70_147 V70 V147 8.382708105019211e-20

R70_148 V70 V148 -930.2561782472552
L70_148 V70 V148 5.952446695901387e-12
C70_148 V70 V148 2.182486766834673e-19

R70_149 V70 V149 1540.1575509449365
L70_149 V70 V149 -8.026427478569654e-13
C70_149 V70 V149 -7.221898940551698e-19

R70_150 V70 V150 -368.65486613435013
L70_150 V70 V150 -8.416116330790409e-11
C70_150 V70 V150 4.333292588729348e-19

R70_151 V70 V151 738.3965127941477
L70_151 V70 V151 -4.861522028202011e-12
C70_151 V70 V151 -1.0991045596465463e-19

R70_152 V70 V152 361.60942745498267
L70_152 V70 V152 -4.730867633894175e-12
C70_152 V70 V152 -1.4583421488658376e-20

R70_153 V70 V153 -2847.4005229182603
L70_153 V70 V153 9.355577821562536e-12
C70_153 V70 V153 6.646977876887752e-20

R70_154 V70 V154 262.02375870339233
L70_154 V70 V154 1.0406878457789237e-11
C70_154 V70 V154 -2.4156590099637946e-19

R70_155 V70 V155 1723.582284147816
L70_155 V70 V155 -5.197683748094081e-12
C70_155 V70 V155 -2.558834651378682e-19

R70_156 V70 V156 -558.4233557710022
L70_156 V70 V156 5.059237196944494e-12
C70_156 V70 V156 -2.1323119514923244e-19

R70_157 V70 V157 -790.2018496422529
L70_157 V70 V157 8.342800692946073e-13
C70_157 V70 V157 7.650269122300899e-19

R70_158 V70 V158 -1455.869726106815
L70_158 V70 V158 -1.2450805497379305e-12
C70_158 V70 V158 -1.1815596558619534e-19

R70_159 V70 V159 -346.11416419971033
L70_159 V70 V159 5.2202431011561704e-12
C70_159 V70 V159 1.3057195659808486e-19

R70_160 V70 V160 -371.4043398309791
L70_160 V70 V160 -1.3951739087675934e-10
C70_160 V70 V160 2.3704679239319257e-20

R70_161 V70 V161 355.24319818416063
L70_161 V70 V161 -9.205546372563008e-12
C70_161 V70 V161 -1.3176753397613603e-19

R70_162 V70 V162 2749.6030978165686
L70_162 V70 V162 1.7433246183696901e-12
C70_162 V70 V162 1.014089320100717e-19

R70_163 V70 V163 398.25944797119325
L70_163 V70 V163 5.119898012493446e-12
C70_163 V70 V163 1.4138023654671377e-19

R70_164 V70 V164 275.03110403612897
L70_164 V70 V164 -1.1778105858203433e-11
C70_164 V70 V164 -7.274861142026963e-21

R70_165 V70 V165 -3168.5438939405376
L70_165 V70 V165 -1.285915517877461e-12
C70_165 V70 V165 -3.309082777212306e-19

R70_166 V70 V166 -1084.1525623823118
L70_166 V70 V166 1.6582704745730884e-11
C70_166 V70 V166 2.5160055358339058e-20

R70_167 V70 V167 2154.532005116498
L70_167 V70 V167 1.6083903086620944e-11
C70_167 V70 V167 -2.711290400999611e-20

R70_168 V70 V168 1281.6404745414725
L70_168 V70 V168 5.953820180050747e-12
C70_168 V70 V168 4.801342275408855e-22

R70_169 V70 V169 -279.67914001452885
L70_169 V70 V169 5.752574593945909e-12
C70_169 V70 V169 2.872679245622737e-19

R70_170 V70 V170 -456.3303462433513
L70_170 V70 V170 -9.436049204211788e-13
C70_170 V70 V170 -1.807994228213314e-19

R70_171 V70 V171 -425.3390806088511
L70_171 V70 V171 -1.3618308315963911e-12
C70_171 V70 V171 -2.6215211751513617e-19

R70_172 V70 V172 -367.7975927833562
L70_172 V70 V172 -4.142504340908324e-12
C70_172 V70 V172 -1.3745052452710896e-19

R70_173 V70 V173 418.1348413022254
L70_173 V70 V173 4.899861715699055e-12
C70_173 V70 V173 2.3601987768724303e-20

R70_174 V70 V174 443.8007542956137
L70_174 V70 V174 7.822637367883777e-13
C70_174 V70 V174 3.4720408941077646e-19

R70_175 V70 V175 12288.100271900916
L70_175 V70 V175 5.655144235338076e-12
C70_175 V70 V175 8.973802820219007e-21

R70_176 V70 V176 1440.1781173924749
L70_176 V70 V176 -1.472730572670063e-11
C70_176 V70 V176 -5.2176740377967487e-20

R70_177 V70 V177 838.501967531958
L70_177 V70 V177 -3.9849584514764996e-12
C70_177 V70 V177 -1.3138915874659606e-19

R70_178 V70 V178 566.0841558339821
L70_178 V70 V178 1.7093316742466646e-11
C70_178 V70 V178 -1.7690657644458797e-20

R70_179 V70 V179 879.777986002384
L70_179 V70 V179 3.123697717499633e-12
C70_179 V70 V179 2.740656806027863e-19

R70_180 V70 V180 948.2142432169886
L70_180 V70 V180 3.498904512015299e-12
C70_180 V70 V180 2.580115652364835e-19

R70_181 V70 V181 -495.96047119743423
L70_181 V70 V181 3.102446818172115e-12
C70_181 V70 V181 6.196332152139291e-20

R70_182 V70 V182 -241.47906340032355
L70_182 V70 V182 -9.433398999315181e-13
C70_182 V70 V182 -1.7683169093807454e-19

R70_183 V70 V183 -2072.0663541710087
L70_183 V70 V183 5.1474271445471454e-12
C70_183 V70 V183 6.250053612938504e-20

R70_184 V70 V184 -2135.231075874725
L70_184 V70 V184 3.164679106748258e-11
C70_184 V70 V184 -8.233021105298343e-20

R70_185 V70 V185 -68647.96098063703
L70_185 V70 V185 -4.0653565187357725e-12
C70_185 V70 V185 3.582494863242303e-20

R70_186 V70 V186 -1582.548700200398
L70_186 V70 V186 1.804572168040145e-12
C70_186 V70 V186 2.5738928631986685e-20

R70_187 V70 V187 2759.2356969077377
L70_187 V70 V187 -4.901748836515122e-12
C70_187 V70 V187 -2.918357283352092e-19

R70_188 V70 V188 1086.598945918441
L70_188 V70 V188 -2.025974846322513e-12
C70_188 V70 V188 -2.0881087766881032e-19

R70_189 V70 V189 1771.144034408135
L70_189 V70 V189 -2.3796744895342373e-12
C70_189 V70 V189 -1.3864429879236995e-19

R70_190 V70 V190 527.8934283438155
L70_190 V70 V190 -2.0282416441874047e-11
C70_190 V70 V190 1.3838818243339679e-19

R70_191 V70 V191 2623.970327984704
L70_191 V70 V191 -1.2546618325623904e-12
C70_191 V70 V191 -1.094475428460004e-19

R70_192 V70 V192 5996.107644270698
L70_192 V70 V192 -4.1617262895196755e-12
C70_192 V70 V192 4.392839012400709e-20

R70_193 V70 V193 1873.4116257749092
L70_193 V70 V193 1.9475444390418915e-12
C70_193 V70 V193 1.4622019632120317e-19

R70_194 V70 V194 -756.1750659622274
L70_194 V70 V194 4.048401514601956e-12
C70_194 V70 V194 2.5738819829709237e-19

R70_195 V70 V195 -1828.1556004312458
L70_195 V70 V195 1.2668872706758892e-12
C70_195 V70 V195 3.2225373085537693e-19

R70_196 V70 V196 -2241.28520676889
L70_196 V70 V196 1.658122173159528e-12
C70_196 V70 V196 1.3697210203199976e-19

R70_197 V70 V197 -2960.20068854633
L70_197 V70 V197 1.3015194134018501e-11
C70_197 V70 V197 -9.118781929876133e-22

R70_198 V70 V198 -629.6884122100817
L70_198 V70 V198 1.3861763504534857e-11
C70_198 V70 V198 -3.4697594970395666e-20

R70_199 V70 V199 -2060.755934219909
L70_199 V70 V199 2.6530209668729284e-12
C70_199 V70 V199 1.2775186668665219e-19

R70_200 V70 V200 1648.70264452064
L70_200 V70 V200 5.18635576057322e-12
C70_200 V70 V200 -7.944602379891698e-20

R71_71 V71 0 420.44563599284925
L71_71 V71 0 3.42710009872664e-13
C71_71 V71 0 1.2612095358396212e-18

R71_72 V71 V72 -2628.1664654518613
L71_72 V71 V72 2.6568716091981137e-11
C71_72 V71 V72 1.2897170267059748e-19

R71_73 V71 V73 -1349.7904167914521
L71_73 V71 V73 1.290585340332248e-11
C71_73 V71 V73 1.129748936123485e-19

R71_74 V71 V74 -4555.326871462738
L71_74 V71 V74 -6.617116432060154e-12
C71_74 V71 V74 -9.904172293193538e-20

R71_75 V71 V75 4219.251171052274
L71_75 V71 V75 7.622517284334157e-13
C71_75 V71 V75 8.689000827215982e-19

R71_76 V71 V76 13165.738558655592
L71_76 V71 V76 6.731257295100404e-12
C71_76 V71 V76 -8.249670470285108e-20

R71_77 V71 V77 -2236.31818435578
L71_77 V71 V77 1.5199647685579315e-11
C71_77 V71 V77 -3.109344737442719e-20

R71_78 V71 V78 1918.3893655097597
L71_78 V71 V78 -8.98842241431017e-12
C71_78 V71 V78 -1.1558256256061361e-19

R71_79 V71 V79 594.7048617560744
L71_79 V71 V79 1.834964638332348e-12
C71_79 V71 V79 3.834735893719452e-19

R71_80 V71 V80 1339.303712844798
L71_80 V71 V80 -4.962835965415783e-12
C71_80 V71 V80 -8.47008150362112e-20

R71_81 V71 V81 712.8181051389923
L71_81 V71 V81 -5.391194414255806e-12
C71_81 V71 V81 -1.2785883775352467e-19

R71_82 V71 V82 -7322.458048559021
L71_82 V71 V82 -7.244800771672075e-11
C71_82 V71 V82 7.798470891289761e-21

R71_83 V71 V83 -1118.2875428259683
L71_83 V71 V83 -9.760414546451202e-13
C71_83 V71 V83 -7.277761277442754e-19

R71_84 V71 V84 -2801.792316101631
L71_84 V71 V84 -1.2732245961724109e-11
C71_84 V71 V84 2.021672309356138e-20

R71_85 V71 V85 -2835.958604025838
L71_85 V71 V85 -4.304810148661423e-12
C71_85 V71 V85 -9.373323299328639e-20

R71_86 V71 V86 -683.4645140479125
L71_86 V71 V86 -4.035593011348087e-12
C71_86 V71 V86 -5.751957635905493e-20

R71_87 V71 V87 -494.5542545780317
L71_87 V71 V87 1.2262339810028317e-12
C71_87 V71 V87 4.676838103238057e-19

R71_88 V71 V88 -1822.2753043674516
L71_88 V71 V88 6.674132101104683e-12
C71_88 V71 V88 4.801074870072207e-20

R71_89 V71 V89 -1147.82753964512
L71_89 V71 V89 3.584614585029821e-12
C71_89 V71 V89 1.3945530316335793e-19

R71_90 V71 V90 1057.9333058528955
L71_90 V71 V90 1.8335148277016445e-12
C71_90 V71 V90 1.8670872282274922e-19

R71_91 V71 V91 342.9565048027725
L71_91 V71 V91 -1.0871975561069374e-12
C71_91 V71 V91 -4.2531408027051807e-19

R71_92 V71 V92 2111.158373271786
L71_92 V71 V92 -2.5580074384649644e-12
C71_92 V71 V92 -1.065234347221326e-19

R71_93 V71 V93 1074.2140732900343
L71_93 V71 V93 6.41226075851737e-12
C71_93 V71 V93 6.892947233163177e-20

R71_94 V71 V94 1143.6119539414467
L71_94 V71 V94 2.0046695358919784e-11
C71_94 V71 V94 -5.3254108292850156e-21

R71_95 V71 V95 669.5252603571791
L71_95 V71 V95 -2.4935222255289704e-12
C71_95 V71 V95 -2.784103643088135e-19

R71_96 V71 V96 1450.9983804838093
L71_96 V71 V96 3.866267641622314e-12
C71_96 V71 V96 1.791037597431601e-20

R71_97 V71 V97 4951.742675226878
L71_97 V71 V97 -3.826957575960553e-12
C71_97 V71 V97 -1.8757401822910502e-19

R71_98 V71 V98 -726.9329667881051
L71_98 V71 V98 -1.9047912931691663e-12
C71_98 V71 V98 -1.9035046746997713e-19

R71_99 V71 V99 -249.2803276532122
L71_99 V71 V99 6.928267892697092e-13
C71_99 V71 V99 7.420096727870768e-19

R71_100 V71 V100 -1813.0369236745885
L71_100 V71 V100 6.936148657147213e-12
C71_100 V71 V100 1.1070589793397321e-19

R71_101 V71 V101 -9188.9919030721
L71_101 V71 V101 1.2821605997144421e-11
C71_101 V71 V101 5.1807013792870865e-20

R71_102 V71 V102 -2599.5876538741727
L71_102 V71 V102 8.223815307818605e-12
C71_102 V71 V102 4.6818472164851104e-20

R71_103 V71 V103 1676.0076006030654
L71_103 V71 V103 -3.601910435495571e-12
C71_103 V71 V103 -1.0035240547813014e-19

R71_104 V71 V104 -1218.7691037382149
L71_104 V71 V104 -2.8214776066836416e-12
C71_104 V71 V104 -1.056057725631132e-19

R71_105 V71 V105 -6954.868750304267
L71_105 V71 V105 1.5033530375471337e-11
C71_105 V71 V105 7.970996622713139e-20

R71_106 V71 V106 2267.060207995015
L71_106 V71 V106 1.844816359670064e-12
C71_106 V71 V106 2.4513455966817e-19

R71_107 V71 V107 446.0414303300043
L71_107 V71 V107 -8.760684290773567e-13
C71_107 V71 V107 -4.853113547332149e-19

R71_108 V71 V108 1721.1014832269443
L71_108 V71 V108 3.3378589294028286e-12
C71_108 V71 V108 5.918322218251357e-20

R71_109 V71 V109 -1848.037509985039
L71_109 V71 V109 -1.5044704854737742e-11
C71_109 V71 V109 -1.399046806061592e-19

R71_110 V71 V110 4436.1433650777335
L71_110 V71 V110 -4.8641735454411115e-12
C71_110 V71 V110 -1.1845405340471955e-19

R71_111 V71 V111 -620.7227120308951
L71_111 V71 V111 2.2869420904987647e-12
C71_111 V71 V111 2.6501828326309458e-20

R71_112 V71 V112 9521.456239680087
L71_112 V71 V112 -1.3581159063442252e-11
C71_112 V71 V112 3.3666116133158934e-20

R71_113 V71 V113 633.9328580666198
L71_113 V71 V113 -5.3527211970927705e-12
C71_113 V71 V113 -2.9039600391067343e-20

R71_114 V71 V114 19518.25303424349
L71_114 V71 V114 -2.3575928902526716e-12
C71_114 V71 V114 -1.9711319348044688e-19

R71_115 V71 V115 -1580.9029758116467
L71_115 V71 V115 1.2363110171615777e-12
C71_115 V71 V115 3.38261647697141e-19

R71_116 V71 V116 -2306.071420053398
L71_116 V71 V116 -3.42752827283426e-11
C71_116 V71 V116 -4.657601166619453e-20

R71_117 V71 V117 1157.714625687353
L71_117 V71 V117 3.727285415959137e-12
C71_117 V71 V117 1.1443158482419392e-19

R71_118 V71 V118 -1424.4774034152376
L71_118 V71 V118 5.306131104162081e-12
C71_118 V71 V118 1.1579442237103457e-19

R71_119 V71 V119 6950.575342461317
L71_119 V71 V119 -1.2157449678882538e-12
C71_119 V71 V119 6.049557693110211e-20

R71_120 V71 V120 8138.769762669271
L71_120 V71 V120 3.5998550574123763e-12
C71_120 V71 V120 1.0052318820396474e-19

R71_121 V71 V121 -532.2791388956223
L71_121 V71 V121 -1.7358668600728946e-11
C71_121 V71 V121 -1.0247738722091593e-19

R71_122 V71 V122 12683.28387537062
L71_122 V71 V122 5.863222037265692e-12
C71_122 V71 V122 4.439220733004027e-20

R71_123 V71 V123 -15944.254762248906
L71_123 V71 V123 -1.1013550693004489e-11
C71_123 V71 V123 -4.484097140495637e-19

R71_124 V71 V124 -34249.405103489284
L71_124 V71 V124 -2.317015280909189e-12
C71_124 V71 V124 -1.057810143023044e-19

R71_125 V71 V125 -1590.0894490978658
L71_125 V71 V125 -5.735723927436086e-12
C71_125 V71 V125 1.62823933966909e-20

R71_126 V71 V126 1366.2416151068862
L71_126 V71 V126 -5.862587568991215e-12
C71_126 V71 V126 -4.1554985337501815e-20

R71_127 V71 V127 610.5099173377963
L71_127 V71 V127 1.58832863553375e-12
C71_127 V71 V127 4.72047198558029e-20

R71_128 V71 V128 18549.60812661669
L71_128 V71 V128 6.22105133328723e-12
C71_128 V71 V128 -2.405966406836351e-20

R71_129 V71 V129 380.3661687077114
L71_129 V71 V129 2.6083196659214977e-11
C71_129 V71 V129 -8.827737170207044e-20

R71_130 V71 V130 -5430.263645260538
L71_130 V71 V130 1.4783537095360944e-11
C71_130 V71 V130 7.208112699798621e-21

R71_131 V71 V131 -483.96634413580523
L71_131 V71 V131 -2.179680485471178e-12
C71_131 V71 V131 2.7091482101127027e-19

R71_132 V71 V132 -1944.5061216506338
L71_132 V71 V132 2.6981045429166323e-11
C71_132 V71 V132 1.8356024413905504e-19

R71_133 V71 V133 268298.91191467724
L71_133 V71 V133 8.695867439380085e-12
C71_133 V71 V133 7.160966679676729e-20

R71_134 V71 V134 -5594.936958454637
L71_134 V71 V134 -6.6240492501047856e-12
C71_134 V71 V134 -3.56810869980495e-20

R71_135 V71 V135 -688.4757053714878
L71_135 V71 V135 5.966470080302899e-12
C71_135 V71 V135 -3.6952856630081905e-19

R71_136 V71 V136 -3604.6718775677236
L71_136 V71 V136 -2.774599314117714e-12
C71_136 V71 V136 -7.184308916018546e-20

R71_137 V71 V137 -538.0368430494996
L71_137 V71 V137 4.446972223491097e-12
C71_137 V71 V137 1.128656772921091e-19

R71_138 V71 V138 2295.3055787012295
L71_138 V71 V138 3.353745859419067e-11
C71_138 V71 V138 -5.2332311918490583e-20

R71_139 V71 V139 323.4363418176855
L71_139 V71 V139 -2.4791025828149496e-11
C71_139 V71 V139 4.0834418750878588e-19

R71_140 V71 V140 769.164087042787
L71_140 V71 V140 1.7743901724197334e-12
C71_140 V71 V140 5.938936631175676e-20

R71_141 V71 V141 -991.5464808177647
L71_141 V71 V141 -2.0085156440906867e-12
C71_141 V71 V141 -2.3800263387429246e-19

R71_142 V71 V142 11989.431581310637
L71_142 V71 V142 3.477028834144665e-12
C71_142 V71 V142 2.17136083463684e-20

R71_143 V71 V143 -3218.4905726632
L71_143 V71 V143 -1.8153362480994185e-12
C71_143 V71 V143 -1.162251548605669e-19

R71_144 V71 V144 -1639.579965267479
L71_144 V71 V144 -4.691771453530015e-12
C71_144 V71 V144 -5.431392066995835e-20

R71_145 V71 V145 376.79799456319523
L71_145 V71 V145 -2.9544422979716754e-12
C71_145 V71 V145 -1.6219705476237645e-19

R71_146 V71 V146 -7461.632363739432
L71_146 V71 V146 -2.4730389512052893e-12
C71_146 V71 V146 9.049560962015964e-20

R71_147 V71 V147 -3755.3760011944087
L71_147 V71 V147 1.3734661869791432e-12
C71_147 V71 V147 -2.834760508940539e-19

R71_148 V71 V148 1788.734641938668
L71_148 V71 V148 -1.8463790553005095e-12
C71_148 V71 V148 -2.6924261525187086e-20

R71_149 V71 V149 3289.735157530222
L71_149 V71 V149 1.0294263386236191e-12
C71_149 V71 V149 4.0374169478113424e-19

R71_150 V71 V150 -824.4727439604391
L71_150 V71 V150 -4.4452758466072095e-12
C71_150 V71 V150 -1.891149281434059e-19

R71_151 V71 V151 -336.41318559247003
L71_151 V71 V151 3.9587839072824675e-12
C71_151 V71 V151 8.757235410323299e-20

R71_152 V71 V152 8331.1316589628
L71_152 V71 V152 3.715366276324153e-12
C71_152 V71 V152 -8.12084756012558e-21

R71_153 V71 V153 -986.7674462919442
L71_153 V71 V153 6.097630627164325e-12
C71_153 V71 V153 6.269018507746505e-20

R71_154 V71 V154 -2552.4215962696962
L71_154 V71 V154 2.7070714914770934e-12
C71_154 V71 V154 6.3472066416147e-20

R71_155 V71 V155 267.86159589477677
L71_155 V71 V155 -2.3772569913289926e-12
C71_155 V71 V155 3.2852462041617073e-19

R71_156 V71 V156 -1262.4933289478165
L71_156 V71 V156 2.5567246938081516e-12
C71_156 V71 V156 5.428543626087201e-20

R71_157 V71 V157 -494.98859183685124
L71_157 V71 V157 -1.305110701677889e-12
C71_157 V71 V157 -2.7708708411336343e-19

R71_158 V71 V158 15437.087854741858
L71_158 V71 V158 9.790355788905368e-12
C71_158 V71 V158 6.949593557787257e-20

R71_159 V71 V159 2656.379083192983
L71_159 V71 V159 -4.260857835712369e-12
C71_159 V71 V159 -1.4097846553786755e-19

R71_160 V71 V160 -1183.3665888952562
L71_160 V71 V160 -4.883018184704531e-12
C71_160 V71 V160 3.2113456359866437e-20

R71_161 V71 V161 536.7937210099755
L71_161 V71 V161 6.951325887834949e-12
C71_161 V71 V161 -6.835518136740553e-20

R71_162 V71 V162 1220.0812549473142
L71_162 V71 V162 5.801570037082108e-12
C71_162 V71 V162 1.2914982377187054e-19

R71_163 V71 V163 636.7144277585601
L71_163 V71 V163 7.561883134127119e-13
C71_163 V71 V163 9.511143230884095e-20

R71_164 V71 V164 623.4798450965598
L71_164 V71 V164 -2.012495313887603e-11
C71_164 V71 V164 3.5276680128063314e-20

R71_165 V71 V165 590.5417621884399
L71_165 V71 V165 4.789325398173676e-12
C71_165 V71 V165 1.0475430411215704e-19

R71_166 V71 V166 -11974.880648736982
L71_166 V71 V166 -1.4065750776755217e-11
C71_166 V71 V166 -1.2857223805359323e-19

R71_167 V71 V167 -262.4450957009789
L71_167 V71 V167 -7.66543518463694e-13
C71_167 V71 V167 -9.214841266483955e-20

R71_168 V71 V168 1216.1968237653984
L71_168 V71 V168 2.396784244056184e-12
C71_168 V71 V168 -7.087588538593085e-20

R71_169 V71 V169 -583.6388364178002
L71_169 V71 V169 -4.775884892787459e-12
C71_169 V71 V169 -3.9159555859878587e-20

R71_170 V71 V170 -1849.3186567772593
L71_170 V71 V170 2.3829154931553955e-11
C71_170 V71 V170 6.237696548000539e-20

R71_171 V71 V171 2474.8805854726143
L71_171 V71 V171 -7.333028015612463e-12
C71_171 V71 V171 4.1608293423386057e-20

R71_172 V71 V172 -944.4757662888437
L71_172 V71 V172 -3.518481607934945e-12
C71_172 V71 V172 -1.6939538670421252e-21

R71_173 V71 V173 -3660.7795447820154
L71_173 V71 V173 5.514087864066612e-12
C71_173 V71 V173 7.42887845605204e-20

R71_174 V71 V174 -7267.12201538906
L71_174 V71 V174 4.668380281905366e-12
C71_174 V71 V174 2.783821907478317e-20

R71_175 V71 V175 410.3856372873233
L71_175 V71 V175 7.0027312680519e-13
C71_175 V71 V175 2.5338278607556136e-19

R71_176 V71 V176 2072.595027836034
L71_176 V71 V176 3.076531430497707e-12
C71_176 V71 V176 1.2960037377004791e-19

R71_177 V71 V177 1246.2340338209967
L71_177 V71 V177 -8.887681561917938e-12
C71_177 V71 V177 -7.471722528641194e-20

R71_178 V71 V178 4216.69436374944
L71_178 V71 V178 -3.009411294911227e-12
C71_178 V71 V178 -7.238424033930957e-20

R71_179 V71 V179 1085.0557161993715
L71_179 V71 V179 -1.3003176960276902e-12
C71_179 V71 V179 -2.4703431773578227e-19

R71_180 V71 V180 -86720.65855207916
L71_180 V71 V180 -2.622465162029022e-12
C71_180 V71 V180 -1.423247167522724e-19

R71_181 V71 V181 -2317.3646709229765
L71_181 V71 V181 3.2280938920789026e-11
C71_181 V71 V181 -7.124789264289125e-20

R71_182 V71 V182 164427.39904897564
L71_182 V71 V182 3.684604843206447e-12
C71_182 V71 V182 8.9013882572312e-20

R71_183 V71 V183 -310.6886582111528
L71_183 V71 V183 -1.8700779787398008e-12
C71_183 V71 V183 1.2896850083952001e-20

R71_184 V71 V184 -2107.310507521202
L71_184 V71 V184 -2.510080506072431e-12
C71_184 V71 V184 -4.657502404122933e-20

R71_185 V71 V185 -2088.150738096988
L71_185 V71 V185 -6.04159958812828e-12
C71_185 V71 V185 1.092334974359799e-19

R71_186 V71 V186 -3371.2833051578527
L71_186 V71 V186 -2.4985309986260643e-11
C71_186 V71 V186 -1.1529686983610612e-19

R71_187 V71 V187 840.5723202206975
L71_187 V71 V187 1.198570631130073e-12
C71_187 V71 V187 1.8368625693878307e-19

R71_188 V71 V188 1040.9260215688305
L71_188 V71 V188 1.3870361316158135e-12
C71_188 V71 V188 1.151765194362991e-19

R71_189 V71 V189 4470.631470999396
L71_189 V71 V189 2.3540323771733713e-11
C71_189 V71 V189 -3.0395713719632095e-20

R71_190 V71 V190 -15055.043060030714
L71_190 V71 V190 -1.0236353043214006e-11
C71_190 V71 V190 -4.906466196174646e-20

R71_191 V71 V191 470.7057407826479
L71_191 V71 V191 8.601548578838221e-12
C71_191 V71 V191 -1.5953926439031105e-19

R71_192 V71 V192 2926.3949563593037
L71_192 V71 V192 -2.4839634917138304e-11
C71_192 V71 V192 -1.466666638012163e-20

R71_193 V71 V193 2358.4323733583756
L71_193 V71 V193 6.4432115351610414e-12
C71_193 V71 V193 4.065348872349655e-23

R71_194 V71 V194 -6528.0300545805285
L71_194 V71 V194 -7.262792823690695e-12
C71_194 V71 V194 -1.5901903905313357e-21

R71_195 V71 V195 -470.82338980059325
L71_195 V71 V195 -4.5396661351740565e-12
C71_195 V71 V195 1.9788265036730743e-19

R71_196 V71 V196 -843.8633270526353
L71_196 V71 V196 -3.0080966592952206e-12
C71_196 V71 V196 -9.301967719000009e-20

R71_197 V71 V197 -1987.0907737034715
L71_197 V71 V197 -3.910277450550279e-12
C71_197 V71 V197 -9.00335623398246e-20

R71_198 V71 V198 -2587.282292257783
L71_198 V71 V198 3.892894217731081e-12
C71_198 V71 V198 1.706862779763196e-20

R71_199 V71 V199 -1037.2891329308745
L71_199 V71 V199 -5.446417522379398e-12
C71_199 V71 V199 4.266623307620397e-20

R71_200 V71 V200 -10816.334059523087
L71_200 V71 V200 1.993904755217699e-11
C71_200 V71 V200 -1.3170462182680628e-21

R72_72 V72 0 139.90582409765815
L72_72 V72 0 2.979308122544291e-13
C72_72 V72 0 1.2340370395318622e-18

R72_73 V72 V73 -1175.8437835333586
L72_73 V72 V73 2.6042142504767698e-11
C72_73 V72 V73 9.903658365749914e-20

R72_74 V72 V74 -3656.9630296411206
L72_74 V72 V74 -3.774183781891915e-12
C72_74 V72 V74 -1.915532196318259e-19

R72_75 V72 V75 -6323.06280651563
L72_75 V72 V75 -4.25261473760506e-12
C72_75 V72 V75 -1.8549512998891332e-19

R72_76 V72 V76 1779.6615439065044
L72_76 V72 V76 6.060626695029698e-13
C72_76 V72 V76 1.0678242908949418e-18

R72_77 V72 V77 -1806.7178603581324
L72_77 V72 V77 1.0964572233728582e-11
C72_77 V72 V77 -3.307039594183065e-20

R72_78 V72 V78 1480.1197108424726
L72_78 V72 V78 -7.306509009719742e-12
C72_78 V72 V78 -1.7015306143207583e-19

R72_79 V72 V79 1311.7065480365754
L72_79 V72 V79 -3.160910145562225e-11
C72_79 V72 V79 -6.599100210155268e-20

R72_80 V72 V80 528.8078508540028
L72_80 V72 V80 2.1823152976317702e-12
C72_80 V72 V80 3.8137560536667096e-19

R72_81 V72 V81 601.3266666534789
L72_81 V72 V81 -1.2647285133753665e-11
C72_81 V72 V81 -3.3769662659201625e-20

R72_82 V72 V82 -3550.8493411740233
L72_82 V72 V82 5.871798974495925e-12
C72_82 V72 V82 1.62709558941922e-19

R72_83 V72 V83 -1734.0956477474544
L72_83 V72 V83 1.806099474807677e-11
C72_83 V72 V83 8.382082284483462e-20

R72_84 V72 V84 -1193.4964910272167
L72_84 V72 V84 -9.406670548480076e-13
C72_84 V72 V84 -8.139475052808525e-19

R72_85 V72 V85 -3098.5659059215254
L72_85 V72 V85 -7.297097067672584e-12
C72_85 V72 V85 -3.9351828228483314e-20

R72_86 V72 V86 -635.8705264017451
L72_86 V72 V86 -4.530719229051029e-12
C72_86 V72 V86 -2.715574717571707e-20

R72_87 V72 V87 -1459.409354383399
L72_87 V72 V87 -4.5374448081782135e-11
C72_87 V72 V87 -9.114330836447712e-21

R72_88 V72 V88 -363.188622284315
L72_88 V72 V88 1.6429825888009356e-12
C72_88 V72 V88 4.2778501570772694e-19

R72_89 V72 V89 -866.5212852609674
L72_89 V72 V89 1.2912697212448821e-11
C72_89 V72 V89 4.895898023819869e-20

R72_90 V72 V90 947.207333124626
L72_90 V72 V90 2.351289084858537e-11
C72_90 V72 V90 -9.715657304796104e-20

R72_91 V72 V91 1159.3093802841447
L72_91 V72 V91 -5.2203833949721215e-12
C72_91 V72 V91 -8.929352304099963e-20

R72_92 V72 V92 260.4457221810075
L72_92 V72 V92 -2.066301222674611e-12
C72_92 V72 V92 -2.267386011404774e-19

R72_93 V72 V93 1135.7444180810812
L72_93 V72 V93 1.2388652783239501e-11
C72_93 V72 V93 3.098965832875268e-20

R72_94 V72 V94 1688.2831580366394
L72_94 V72 V94 4.289475799343417e-12
C72_94 V72 V94 1.1272401765654552e-19

R72_95 V72 V95 1687.2281953920228
L72_95 V72 V95 6.197715919804809e-12
C72_95 V72 V95 5.510451186966476e-20

R72_96 V72 V96 466.41443473138685
L72_96 V72 V96 -4.170336393021019e-12
C72_96 V72 V96 -2.228400176644614e-19

R72_97 V72 V97 2555.822210810602
L72_97 V72 V97 1.3619808984436418e-11
C72_97 V72 V97 -2.2065966905792333e-20

R72_98 V72 V98 -877.7131858230707
L72_98 V72 V98 -4.058448955562038e-12
C72_98 V72 V98 -4.133930608910253e-20

R72_99 V72 V99 -753.0400913861399
L72_99 V72 V99 1.5906350489155499e-10
C72_99 V72 V99 3.2249086749775345e-20

R72_100 V72 V100 -177.63367168697593
L72_100 V72 V100 1.1738816292133133e-12
C72_100 V72 V100 4.735501845749542e-19

R72_101 V72 V101 -6595.732885394215
L72_101 V72 V101 -6.978616568113715e-12
C72_101 V72 V101 -4.200767667718505e-20

R72_102 V72 V102 -3748.0119130469106
L72_102 V72 V102 -8.317428510061804e-12
C72_102 V72 V102 -1.0635798369174192e-19

R72_103 V72 V103 -1883.6282885365513
L72_103 V72 V103 -4.539673820972914e-12
C72_103 V72 V103 -9.925492897658045e-20

R72_104 V72 V104 1986.436790167379
L72_104 V72 V104 -8.585540185745575e-12
C72_104 V72 V104 -5.656580886700541e-20

R72_105 V72 V105 -2334.866153697923
L72_105 V72 V105 -9.743575287084711e-12
C72_105 V72 V105 2.5391749581364305e-20

R72_106 V72 V106 -3408.9086917420095
L72_106 V72 V106 2.7460357913020548e-12
C72_106 V72 V106 1.7975060192553838e-19

R72_107 V72 V107 1034.1871229458616
L72_107 V72 V107 1.140094123594147e-11
C72_107 V72 V107 2.249879739891141e-20

R72_108 V72 V108 260.0525639490323
L72_108 V72 V108 -1.1773443683830844e-12
C72_108 V72 V108 -3.1463862030320587e-19

R72_109 V72 V109 -5304.078652621973
L72_109 V72 V109 1.0232364400026145e-11
C72_109 V72 V109 -4.1831946352983564e-20

R72_110 V72 V110 1010.8457740096883
L72_110 V72 V110 -1.251143451267178e-10
C72_110 V72 V110 -9.778325721488745e-21

R72_111 V72 V111 -5060.372040393668
L72_111 V72 V111 1.700867470255745e-11
C72_111 V72 V111 5.718422277640837e-20

R72_112 V72 V112 -393.99788797372867
L72_112 V72 V112 3.103503174934933e-12
C72_112 V72 V112 -1.0796477660263887e-20

R72_113 V72 V113 504.30066184877484
L72_113 V72 V113 -5.2576541138108377e-11
C72_113 V72 V113 7.78087406016931e-21

R72_114 V72 V114 2985.000438306234
L72_114 V72 V114 -8.186084561623346e-12
C72_114 V72 V114 -7.861140820425262e-20

R72_115 V72 V115 -5746.201277137016
L72_115 V72 V115 -2.233186457576842e-11
C72_115 V72 V115 -5.039844654905518e-20

R72_116 V72 V116 -558.4881619128251
L72_116 V72 V116 1.6023860270578312e-12
C72_116 V72 V116 2.406483620556495e-19

R72_117 V72 V117 2149.388363035017
L72_117 V72 V117 6.053897479300595e-12
C72_117 V72 V117 5.3566418040166375e-20

R72_118 V72 V118 -536.5008008064112
L72_118 V72 V118 -1.0313103647926369e-11
C72_118 V72 V118 -3.7512243812787873e-20

R72_119 V72 V119 11557.940289120097
L72_119 V72 V119 5.168502385688532e-12
C72_119 V72 V119 4.4985250072749384e-20

R72_120 V72 V120 434.19360445123704
L72_120 V72 V120 -1.1625884879740798e-12
C72_120 V72 V120 5.535986777387115e-20

R72_121 V72 V121 -601.6392182899054
L72_121 V72 V121 -3.380585059393751e-12
C72_121 V72 V121 -1.226393825784275e-19

R72_122 V72 V122 1236.3588410854213
L72_122 V72 V122 6.809997213976138e-12
C72_122 V72 V122 8.06220638244061e-20

R72_123 V72 V123 -9406.572513082412
L72_123 V72 V123 -4.571957726507577e-12
C72_123 V72 V123 -6.937390591524573e-21

R72_124 V72 V124 -1090.4458074951676
L72_124 V72 V124 5.147446277085719e-12
C72_124 V72 V124 -3.3025212255747383e-19

R72_125 V72 V125 -6370.761876350596
L72_125 V72 V125 -5.2890165281932924e-12
C72_125 V72 V125 2.0354861824167772e-20

R72_126 V72 V126 683.8388820355906
L72_126 V72 V126 5.471982690915708e-12
C72_126 V72 V126 1.2681903900742932e-19

R72_127 V72 V127 1546.2504792590544
L72_127 V72 V127 9.752719270053708e-11
C72_127 V72 V127 3.3462218328893037e-20

R72_128 V72 V128 2660.6485025415705
L72_128 V72 V128 1.652528365439186e-12
C72_128 V72 V128 5.793216264386719e-21

R72_129 V72 V129 416.1011582644019
L72_129 V72 V129 2.389803151700088e-12
C72_129 V72 V129 7.335847630319409e-20

R72_130 V72 V130 -1065.126051820875
L72_130 V72 V130 -1.0120219690593445e-11
C72_130 V72 V130 -1.252575467657392e-19

R72_131 V72 V131 -1069.46082439795
L72_131 V72 V131 -2.731513726097316e-11
C72_131 V72 V131 -4.644592657614542e-20

R72_132 V72 V132 -799.6643847717137
L72_132 V72 V132 -1.3816056715487425e-12
C72_132 V72 V132 2.660384980695094e-19

R72_133 V72 V133 -5431.050271352728
L72_133 V72 V133 -2.7158623259527358e-11
C72_133 V72 V133 -2.959347260746701e-20

R72_134 V72 V134 5446.210136225906
L72_134 V72 V134 -3.807242859397409e-11
C72_134 V72 V134 1.0046337467244453e-19

R72_135 V72 V135 5014.644059473047
L72_135 V72 V135 -2.917936812129059e-11
C72_135 V72 V135 2.9593843269666985e-20

R72_136 V72 V136 -524.2901490709722
L72_136 V72 V136 1.902671390956154e-11
C72_136 V72 V136 -2.3559984561718157e-19

R72_137 V72 V137 -653.3580267635549
L72_137 V72 V137 2.8790815680802147e-11
C72_137 V72 V137 -2.756777905418043e-20

R72_138 V72 V138 2107.307611378181
L72_138 V72 V138 5.239051955500934e-12
C72_138 V72 V138 -3.828040768027567e-20

R72_139 V72 V139 847.4888167013206
L72_139 V72 V139 2.294595394099917e-12
C72_139 V72 V139 -1.1892686975079517e-21

R72_140 V72 V140 271.48814645646354
L72_140 V72 V140 3.879374384229075e-12
C72_140 V72 V140 2.0611315068839321e-19

R72_141 V72 V141 -1004.5653482894243
L72_141 V72 V141 -5.032403266506574e-12
C72_141 V72 V141 8.109469099189676e-21

R72_142 V72 V142 -4107.26872409699
L72_142 V72 V142 1.0364168529545e-11
C72_142 V72 V142 -4.891543434134763e-20

R72_143 V72 V143 -919.3772419553649
L72_143 V72 V143 -4.41476290015906e-12
C72_143 V72 V143 4.601127848326745e-21

R72_144 V72 V144 1141.952488387623
L72_144 V72 V144 -4.546883585936688e-12
C72_144 V72 V144 3.5013546960630085e-21

R72_145 V72 V145 418.4241146276576
L72_145 V72 V145 -4.511576021267957e-12
C72_145 V72 V145 -3.61910453042954e-20

R72_146 V72 V146 18167.57888656482
L72_146 V72 V146 -2.2453681451380136e-12
C72_146 V72 V146 8.525289615833732e-20

R72_147 V72 V147 2427.2120547409454
L72_147 V72 V147 -4.680315764792844e-12
C72_147 V72 V147 -2.3257367712210608e-20

R72_148 V72 V148 -230.49367087520807
L72_148 V72 V148 5.361756192060218e-12
C72_148 V72 V148 -2.251594287444854e-19

R72_149 V72 V149 1886.356591829305
L72_149 V72 V149 2.3711057282645934e-12
C72_149 V72 V149 -1.9756926180429303e-20

R72_150 V72 V150 -963.5708336206774
L72_150 V72 V150 -8.287116792400475e-12
C72_150 V72 V150 -3.836971393461936e-20

R72_151 V72 V151 18862.998899834925
L72_151 V72 V151 7.786341990344803e-12
C72_151 V72 V151 -3.251743004071855e-20

R72_152 V72 V152 1489.0211638758965
L72_152 V72 V152 1.5753122209182324e-12
C72_152 V72 V152 7.514380594015642e-20

R72_153 V72 V153 -2149.833197783618
L72_153 V72 V153 7.446967697172632e-12
C72_153 V72 V153 8.395706564234726e-20

R72_154 V72 V154 5388.84234166439
L72_154 V72 V154 2.5581253060761855e-12
C72_154 V72 V154 -5.047673901901586e-20

R72_155 V72 V155 5915.372963804393
L72_155 V72 V155 3.860511549950498e-12
C72_155 V72 V155 5.282773781023192e-21

R72_156 V72 V156 -960.1872828528988
L72_156 V72 V156 -7.824031689689715e-13
C72_156 V72 V156 1.3470381033216262e-19

R72_157 V72 V157 -371.6540719627155
L72_157 V72 V157 -2.8542315340832745e-12
C72_157 V72 V157 -5.968962189741244e-20

R72_158 V72 V158 -961.1666821946034
L72_158 V72 V158 -1.0886451048062188e-11
C72_158 V72 V158 2.2318210984253844e-20

R72_159 V72 V159 -529.1857179405685
L72_159 V72 V159 -2.290521296512515e-12
C72_159 V72 V159 2.1116454873878776e-20

R72_160 V72 V160 376.7662706507997
L72_160 V72 V160 -4.626221838230387e-12
C72_160 V72 V160 -5.354983390040303e-20

R72_161 V72 V161 512.0281190076049
L72_161 V72 V161 1.5953809376471163e-11
C72_161 V72 V161 -4.2083434951540415e-20

R72_162 V72 V162 991.401044512341
L72_162 V72 V162 -8.84469421649062e-12
C72_162 V72 V162 4.9286830269831204e-20

R72_163 V72 V163 676.6856233154151
L72_163 V72 V163 -1.891050706944463e-11
C72_163 V72 V163 4.882456748072994e-21

R72_164 V72 V164 17405.31390002562
L72_164 V72 V164 5.986518746481067e-13
C72_164 V72 V164 5.906502027878499e-20

R72_165 V72 V165 811.596857195393
L72_165 V72 V165 -1.8977387661119803e-11
C72_165 V72 V165 -2.437854405657004e-20

R72_166 V72 V166 7639.150879861899
L72_166 V72 V166 5.6518153898151917e-11
C72_166 V72 V166 -1.1385337073229044e-19

R72_167 V72 V167 -1424.2719928090785
L72_167 V72 V167 2.283957103456362e-12
C72_167 V72 V167 -8.608097613242212e-21

R72_168 V72 V168 -1088.0692933698667
L72_168 V72 V168 -7.013123805857461e-13
C72_168 V72 V168 -7.23641059739569e-20

R72_169 V72 V169 -592.473141781326
L72_169 V72 V169 -3.566697971653302e-12
C72_169 V72 V169 -3.986365557542806e-20

R72_170 V72 V170 -705.4203599191268
L72_170 V72 V170 -6.778276476122839e-12
C72_170 V72 V170 -9.203416603437971e-21

R72_171 V72 V171 -1420.240577198507
L72_171 V72 V171 -2.9860644202508266e-12
C72_171 V72 V171 -6.773780310957807e-20

R72_172 V72 V172 -561.197897890725
L72_172 V72 V172 -1.815640953646004e-12
C72_172 V72 V172 2.1659744463447286e-20

R72_173 V72 V173 -3053.557189105706
L72_173 V72 V173 4.783076295202035e-12
C72_173 V72 V173 6.851997484221392e-20

R72_174 V72 V174 3974.6760343287624
L72_174 V72 V174 7.519765694453336e-12
C72_174 V72 V174 9.309606680484317e-20

R72_175 V72 V175 8794.55788484754
L72_175 V72 V175 -1.1018208077724028e-11
C72_175 V72 V175 5.284049766168285e-20

R72_176 V72 V176 401.17376448974596
L72_176 V72 V176 5.661804270125018e-13
C72_176 V72 V176 1.8926416886365158e-19

R72_177 V72 V177 1358.1096537133656
L72_177 V72 V177 1.4028316895861825e-11
C72_177 V72 V177 -7.966223301136976e-20

R72_178 V72 V178 1188.5955049578768
L72_178 V72 V178 4.7086681557024135e-11
C72_178 V72 V178 -1.2220047407992745e-20

R72_179 V72 V179 5825.5633608292355
L72_179 V72 V179 1.0162884697290326e-11
C72_179 V72 V179 1.0381649386788119e-20

R72_180 V72 V180 447.81196524465514
L72_180 V72 V180 -1.3955156574575769e-12
C72_180 V72 V180 -1.691273709893268e-19

R72_181 V72 V181 -2290.5391811660043
L72_181 V72 V181 -6.949314420118946e-12
C72_181 V72 V181 -4.4526836700629435e-21

R72_182 V72 V182 -1442.8024653738676
L72_182 V72 V182 -5.579600499463702e-12
C72_182 V72 V182 -3.0413006830017206e-20

R72_183 V72 V183 -7262.923520275203
L72_183 V72 V183 -5.187339153655236e-12
C72_183 V72 V183 -2.032821157859602e-20

R72_184 V72 V184 -287.09892408258463
L72_184 V72 V184 -2.436364508393706e-12
C72_184 V72 V184 7.389864208426438e-20

R72_185 V72 V185 -1647.3145984332436
L72_185 V72 V185 -4.093655100140821e-12
C72_185 V72 V185 6.018441123215854e-20

R72_186 V72 V186 -1167.1923896855308
L72_186 V72 V186 -2.1962696652495283e-11
C72_186 V72 V186 3.88380166011953e-21

R72_187 V72 V187 2642.901670451687
L72_187 V72 V187 4.365782021776394e-11
C72_187 V72 V187 2.659761747978848e-20

R72_188 V72 V188 729.3928755562554
L72_188 V72 V188 1.413409656230233e-12
C72_188 V72 V188 -7.309076432345142e-21

R72_189 V72 V189 4109.882190676813
L72_189 V72 V189 9.351565491531715e-12
C72_189 V72 V189 -7.278706624434762e-20

R72_190 V72 V190 2772.2397495058303
L72_190 V72 V190 -4.450992778624211e-10
C72_190 V72 V190 -1.2569145453771312e-20

R72_191 V72 V191 3010.5246215166585
L72_191 V72 V191 2.846531268905732e-11
C72_191 V72 V191 -5.2024001025643996e-20

R72_192 V72 V192 415.38979819263454
L72_192 V72 V192 -5.221372598810284e-12
C72_192 V72 V192 -1.1627296741007012e-19

R72_193 V72 V193 1218.400583115343
L72_193 V72 V193 5.800452492246962e-12
C72_193 V72 V193 2.310414344029999e-20

R72_194 V72 V194 -5057.052324895908
L72_194 V72 V194 -8.62061934973321e-12
C72_194 V72 V194 -2.9187233901864185e-20

R72_195 V72 V195 -1584.8338142637308
L72_195 V72 V195 -5.049395317165091e-12
C72_195 V72 V195 -3.313154374422542e-20

R72_196 V72 V196 -383.86959233038453
L72_196 V72 V196 2.970555039425449e-12
C72_196 V72 V196 2.856401210022575e-19

R72_197 V72 V197 -3430.5668866336982
L72_197 V72 V197 -8.601097403563145e-12
C72_197 V72 V197 2.4883344160600446e-20

R72_198 V72 V198 -1054.9134067917878
L72_198 V72 V198 6.480174064442288e-12
C72_198 V72 V198 -6.076316894576462e-20

R72_199 V72 V199 -643.7199787841862
L72_199 V72 V199 5.033917342531114e-12
C72_199 V72 V199 8.224413188735207e-21

R72_200 V72 V200 -2521.1511885209543
L72_200 V72 V200 -3.6811879284362484e-12
C72_200 V72 V200 -2.6852028739886683e-20

R73_73 V73 0 222.56458634595694
L73_73 V73 0 7.427555898826702e-12
C73_73 V73 0 2.962508836351812e-19

R73_74 V73 V74 -3426.0827167218463
L73_74 V73 V74 -9.808249151452725e-12
C73_74 V73 V74 -8.07720628479941e-20

R73_75 V73 V75 14466.888198005816
L73_75 V73 V75 -4.135444823097079e-12
C73_75 V73 V75 -2.010868092863495e-19

R73_76 V73 V76 3527.4102325436
L73_76 V73 V76 -3.557830352939566e-11
C73_76 V73 V76 -6.44602188480078e-20

R73_77 V73 V77 -1009.8633972519948
L73_77 V73 V77 1.8382265977430744e-12
C73_77 V73 V77 1.5411636674055096e-19

R73_78 V73 V78 775.2367731671063
L73_78 V73 V78 -2.051105757545977e-11
C73_78 V73 V78 -1.5557053252715327e-20

R73_79 V73 V79 704.7521023742223
L73_79 V73 V79 9.793761657366692e-12
C73_79 V73 V79 4.4034223799372235e-20

R73_80 V73 V80 642.7548121167423
L73_80 V73 V80 -5.157700502752485e-11
C73_80 V73 V80 -1.0102176233244851e-20

R73_81 V73 V81 284.36966319982696
L73_81 V73 V81 3.867503066352269e-12
C73_81 V73 V81 3.592139694642874e-19

R73_82 V73 V82 -1688.0814253446636
L73_82 V73 V82 6.1299095456733036e-12
C73_82 V73 V82 5.772338210533517e-20

R73_83 V73 V83 -832.227259787153
L73_83 V73 V83 8.87072464222951e-12
C73_83 V73 V83 4.8595921134760315e-20

R73_84 V73 V84 -1144.2574883751158
L73_84 V73 V84 1.20682795393867e-11
C73_84 V73 V84 4.0620579113458433e-20

R73_85 V73 V85 -1564.2314388091158
L73_85 V73 V85 -1.916438938788105e-12
C73_85 V73 V85 -3.9973906362758877e-19

R73_86 V73 V86 -350.0762311316738
L73_86 V73 V86 5.82688153709332e-11
C73_86 V73 V86 -1.7673617381912948e-20

R73_87 V73 V87 -1056.740804212639
L73_87 V73 V87 3.4884810620380145e-11
C73_87 V73 V87 6.417410830143286e-20

R73_88 V73 V88 -831.5659937898943
L73_88 V73 V88 1.4078515736447183e-11
C73_88 V73 V88 1.2927682237372746e-19

R73_89 V73 V89 -341.4058099015006
L73_89 V73 V89 6.6022694319601125e-12
C73_89 V73 V89 3.466449379178999e-19

R73_90 V73 V90 398.76782820979383
L73_90 V73 V90 -4.331265956569517e-12
C73_90 V73 V90 -2.6526373803543844e-21

R73_91 V73 V91 457.77692031932577
L73_91 V73 V91 -4.399838779488499e-12
C73_91 V73 V91 -1.1786209693809416e-19

R73_92 V73 V92 554.6869990592041
L73_92 V73 V92 -3.4949321012654784e-12
C73_92 V73 V92 -1.5128291943668934e-19

R73_93 V73 V93 305.9534274503193
L73_93 V73 V93 2.1230077662706905e-12
C73_93 V73 V93 1.0152502822846817e-19

R73_94 V73 V94 928.1082880406383
L73_94 V73 V94 4.399410976124881e-12
C73_94 V73 V94 7.434950705141746e-20

R73_95 V73 V95 2953.2503078214368
L73_95 V73 V95 1.0806057590001443e-11
C73_95 V73 V95 -5.81351651532967e-20

R73_96 V73 V96 1212.6700713252724
L73_96 V73 V96 5.290211661634275e-12
C73_96 V73 V96 -6.459435651710695e-20

R73_97 V73 V97 -1104.4134383717294
L73_97 V73 V97 -1.3847257977531263e-12
C73_97 V73 V97 -6.650926169453643e-19

R73_98 V73 V98 -358.71599700756576
L73_98 V73 V98 -1.4234005287055267e-11
C73_98 V73 V98 -1.6115377598897963e-19

R73_99 V73 V99 -477.6644992791117
L73_99 V73 V99 5.571611046723793e-12
C73_99 V73 V99 1.822914577574704e-19

R73_100 V73 V100 -567.3903280438695
L73_100 V73 V100 9.494126560148697e-12
C73_100 V73 V100 2.108222137134191e-19

R73_101 V73 V101 -511.8083286278954
L73_101 V73 V101 1.1451832661229859e-11
C73_101 V73 V101 3.4386383072967977e-19

R73_102 V73 V102 5592.160292026309
L73_102 V73 V102 -5.967584422965904e-12
C73_102 V73 V102 -8.280488277483135e-20

R73_103 V73 V103 -16023.976147110669
L73_103 V73 V103 -1.0189625933626121e-11
C73_103 V73 V103 -6.818337355224743e-20

R73_104 V73 V104 -1964.2354732613126
L73_104 V73 V104 -1.9949105158157725e-11
C73_104 V73 V104 -4.2403514099572163e-20

R73_105 V73 V105 292.09984212680604
L73_105 V73 V105 2.5065860678767175e-12
C73_105 V73 V105 8.457395200904538e-20

R73_106 V73 V106 1804.3381446848791
L73_106 V73 V106 4.874395433783805e-12
C73_106 V73 V106 2.9574643079203757e-19

R73_107 V73 V107 957.4494486680342
L73_107 V73 V107 -9.478164202106495e-12
C73_107 V73 V107 -1.0783178295068479e-19

R73_108 V73 V108 903.1715974937576
L73_108 V73 V108 -1.1390957717964666e-11
C73_108 V73 V108 -7.39860721463285e-20

R73_109 V73 V109 -1393.1846206981206
L73_109 V73 V109 -1.984196000138678e-12
C73_109 V73 V109 -2.2597175735265882e-19

R73_110 V73 V110 9866.894998183358
L73_110 V73 V110 2.460971372523192e-11
C73_110 V73 V110 -1.0223768605325147e-19

R73_111 V73 V111 -6682.041921767394
L73_111 V73 V111 -2.5669273883646143e-11
C73_111 V73 V111 9.271824674027696e-20

R73_112 V73 V112 -7830.122920792037
L73_112 V73 V112 -8.56310496165646e-12
C73_112 V73 V112 -2.6924528636609702e-20

R73_113 V73 V113 -637.3072053628733
L73_113 V73 V113 1.9436262311775206e-12
C73_113 V73 V113 3.1491460909573103e-19

R73_114 V73 V114 28789.362243265536
L73_114 V73 V114 -4.928099750352585e-12
C73_114 V73 V114 -1.973240936063427e-19

R73_115 V73 V115 -2027.7497837261396
L73_115 V73 V115 1.277240942814286e-11
C73_115 V73 V115 -4.620286567594174e-20

R73_116 V73 V116 -1345.506361143132
L73_116 V73 V116 4.823773237607173e-12
C73_116 V73 V116 5.0802304361080256e-21

R73_117 V73 V117 457.4639580512661
L73_117 V73 V117 -9.270798730074818e-12
C73_117 V73 V117 -3.6802236499256e-19

R73_118 V73 V118 -1105.8514596622053
L73_118 V73 V118 1.0840655051342978e-11
C73_118 V73 V118 1.2513627698423568e-19

R73_119 V73 V119 -4395.675185359686
L73_119 V73 V119 9.20407764848757e-12
C73_119 V73 V119 5.773152767762885e-20

R73_120 V73 V120 -17382.58117461465
L73_120 V73 V120 6.37389142958122e-11
C73_120 V73 V120 8.750387104243049e-20

R73_121 V73 V121 -4972.5511529210235
L73_121 V73 V121 -3.5665861352127966e-12
C73_121 V73 V121 1.5709037151309427e-19

R73_122 V73 V122 4861.164386068745
L73_122 V73 V122 3.4298513748726953e-11
C73_122 V73 V122 4.8188013632260834e-20

R73_123 V73 V123 3264.357492751419
L73_123 V73 V123 -4.938768829724946e-12
C73_123 V73 V123 -6.853517461588424e-20

R73_124 V73 V124 2025.2650232181275
L73_124 V73 V124 -4.4760722832268e-12
C73_124 V73 V124 -1.4635837336867917e-19

R73_125 V73 V125 -937.8576836633777
L73_125 V73 V125 9.478004955203329e-12
C73_125 V73 V125 1.9155011373860853e-19

R73_126 V73 V126 1120.5247929206485
L73_126 V73 V126 -1.4411385152578652e-11
C73_126 V73 V126 5.2700017466107135e-20

R73_127 V73 V127 1514.0619126640852
L73_127 V73 V127 -2.2368322105862623e-11
C73_127 V73 V127 -1.3767910737979283e-20

R73_128 V73 V128 2539.2470242317067
L73_128 V73 V128 6.352340991350093e-11
C73_128 V73 V128 4.0774886867669994e-20

R73_129 V73 V129 591.5283614783016
L73_129 V73 V129 1.0522161310724841e-11
C73_129 V73 V129 -2.9641822359071623e-19

R73_130 V73 V130 -2027.9783245636017
L73_130 V73 V130 1.3682358197632912e-11
C73_130 V73 V130 -8.007376095714407e-20

R73_131 V73 V131 -855.1344924162928
L73_131 V73 V131 4.7099392376360785e-12
C73_131 V73 V131 7.929902641281466e-20

R73_132 V73 V132 -683.6984219204388
L73_132 V73 V132 2.9959015321822488e-12
C73_132 V73 V132 1.1055338309383044e-19

R73_133 V73 V133 -5089.404171006757
L73_133 V73 V133 -1.249540893229018e-10
C73_133 V73 V133 2.1796078912069054e-19

R73_134 V73 V134 -2176.1391245502164
L73_134 V73 V134 -2.5167151588626427e-11
C73_134 V73 V134 5.543163429496557e-20

R73_135 V73 V135 18236.606411385223
L73_135 V73 V135 -9.466957297426053e-12
C73_135 V73 V135 -6.307274914949792e-20

R73_136 V73 V136 -12759.631411438295
L73_136 V73 V136 -8.101284220952428e-12
C73_136 V73 V136 -2.281300768137003e-19

R73_137 V73 V137 -1250.5767751188744
L73_137 V73 V137 6.246114846698629e-12
C73_137 V73 V137 -3.6253177783156805e-20

R73_138 V73 V138 1268.1693478620914
L73_138 V73 V138 2.7837282366866643e-11
C73_138 V73 V138 -1.597782282219936e-20

R73_139 V73 V139 1681.7223240597416
L73_139 V73 V139 -6.872185764787033e-11
C73_139 V73 V139 9.197835953876492e-20

R73_140 V73 V140 1342.760899127991
L73_140 V73 V140 -1.020038835546681e-11
C73_140 V73 V140 2.284008349187538e-19

R73_141 V73 V141 -3471.5476604979276
L73_141 V73 V141 -3.051347019103388e-12
C73_141 V73 V141 -2.501803605127031e-19

R73_142 V73 V142 4985.918069371078
L73_142 V73 V142 -4.012502724426059e-12
C73_142 V73 V142 -5.60246357369886e-20

R73_143 V73 V143 -2981.4549941377154
L73_143 V73 V143 2.2935113371008683e-11
C73_143 V73 V143 -6.10901334948414e-20

R73_144 V73 V144 8691.891321563528
L73_144 V73 V144 7.60639781136792e-12
C73_144 V73 V144 1.0368760006074891e-21

R73_145 V73 V145 496.3194491512826
L73_145 V73 V145 -8.424960075199685e-12
C73_145 V73 V145 1.879221023709177e-19

R73_146 V73 V146 -1275.7647657730893
L73_146 V73 V146 3.3250589042059874e-12
C73_146 V73 V146 5.217294272816203e-20

R73_147 V73 V147 1543.3279022574193
L73_147 V73 V147 -2.529317750170334e-11
C73_147 V73 V147 -3.2434124453773796e-20

R73_148 V73 V148 -3878.8115570406844
L73_148 V73 V148 -3.590798740047106e-12
C73_148 V73 V148 -1.6397504977261582e-19

R73_149 V73 V149 -626.5187264700583
L73_149 V73 V149 2.8236722602459667e-12
C73_149 V73 V149 8.250629335148425e-20

R73_150 V73 V150 -1352.185193427838
L73_150 V73 V150 -1.4325591297340698e-11
C73_150 V73 V150 -3.4100643506649635e-20

R73_151 V73 V151 -1825.227257184229
L73_151 V73 V151 -7.679655400856776e-12
C73_151 V73 V151 3.52509270699652e-20

R73_152 V73 V152 3227.5727538457386
L73_152 V73 V152 2.4697481017519294e-11
C73_152 V73 V152 6.13102647756029e-20

R73_153 V73 V153 4388.5670212336545
L73_153 V73 V153 -2.243830890221186e-11
C73_153 V73 V153 -9.674346930788001e-20

R73_154 V73 V154 5180.749225420722
L73_154 V73 V154 -5.880461026023272e-11
C73_154 V73 V154 -4.395527080600578e-20

R73_155 V73 V155 3015.7508346253353
L73_155 V73 V155 4.6557489330394896e-12
C73_155 V73 V155 9.159762363335067e-20

R73_156 V73 V156 -612.4032435900257
L73_156 V73 V156 1.2657954676885619e-11
C73_156 V73 V156 5.365595395453584e-20

R73_157 V73 V157 -6753.430848188625
L73_157 V73 V157 -3.577689195620576e-11
C73_157 V73 V157 -1.3459633004428262e-19

R73_158 V73 V158 40121.888558945444
L73_158 V73 V158 -1.0278380723761595e-11
C73_158 V73 V158 3.130954494486938e-20

R73_159 V73 V159 -1647.587702710507
L73_159 V73 V159 -6.205905907045884e-11
C73_159 V73 V159 -1.2312748147386162e-19

R73_160 V73 V160 2025.5926596443426
L73_160 V73 V160 5.590366870783231e-10
C73_160 V73 V160 -9.997224620531465e-20

R73_161 V73 V161 668.5570076207564
L73_161 V73 V161 3.316054549082594e-12
C73_161 V73 V161 1.1818358365066882e-19

R73_162 V73 V162 -6417.845357388448
L73_162 V73 V162 5.02251257065028e-12
C73_162 V73 V162 -8.89843681297926e-21

R73_163 V73 V163 1722.8695909948945
L73_163 V73 V163 -4.271143955820913e-11
C73_163 V73 V163 -1.5415732700225676e-20

R73_164 V73 V164 1074.060471106994
L73_164 V73 V164 -2.0930469829420736e-11
C73_164 V73 V164 7.160108130420787e-20

R73_165 V73 V165 2289.698199525566
L73_165 V73 V165 -1.4064844887014532e-12
C73_165 V73 V165 -9.67483337167406e-20

R73_166 V73 V166 -1021.0389415905922
L73_166 V73 V166 -2.3113781370143625e-12
C73_166 V73 V166 -5.918380020784933e-20

R73_167 V73 V167 -1087.150470345674
L73_167 V73 V167 3.99847917490861e-11
C73_167 V73 V167 7.354894696703531e-20

R73_168 V73 V168 -1408.5728526133341
L73_168 V73 V168 7.519786288144136e-12
C73_168 V73 V168 8.867760471461026e-20

R73_169 V73 V169 -1573.1154313445656
L73_169 V73 V169 3.1312470708593636e-12
C73_169 V73 V169 4.581369795808069e-20

R73_170 V73 V170 1541.8565741575244
L73_170 V73 V170 2.4717703762933747e-12
C73_170 V73 V170 1.082040996737299e-19

R73_171 V73 V171 3858.6332223338554
L73_171 V73 V171 3.905108530896725e-11
C73_171 V73 V171 5.0860963476705414e-20

R73_172 V73 V172 -1558.0698408269334
L73_172 V73 V172 -7.82493434797719e-12
C73_172 V73 V172 -2.5951273108036544e-22

R73_173 V73 V173 3784.53814646406
L73_173 V73 V173 4.495642363113602e-12
C73_173 V73 V173 -1.1265951537271465e-19

R73_174 V73 V174 2712.2970336837047
L73_174 V73 V174 7.531357066422557e-12
C73_174 V73 V174 -1.3008774812837362e-19

R73_175 V73 V175 2892.0033693368655
L73_175 V73 V175 -7.001286155103068e-12
C73_175 V73 V175 -4.288603377524986e-20

R73_176 V73 V176 926.1763900865019
L73_176 V73 V176 8.744607149166049e-12
C73_176 V73 V176 6.352957741289118e-23

R73_177 V73 V177 2330.2897757117016
L73_177 V73 V177 -2.5688252232924893e-12
C73_177 V73 V177 -9.207873522866751e-21

R73_178 V73 V178 -7068.482437758893
L73_178 V73 V178 -2.8248470679447212e-12
C73_178 V73 V178 5.524265322654577e-22

R73_179 V73 V179 -15571.8438743864
L73_179 V73 V179 1.084023141758992e-11
C73_179 V73 V179 -5.1285129020004644e-20

R73_180 V73 V180 7986.785056333837
L73_180 V73 V180 -1.8698910429405617e-11
C73_180 V73 V180 -1.0530397505990672e-19

R73_181 V73 V181 -2429.3223062426
L73_181 V73 V181 1.2888086959863344e-12
C73_181 V73 V181 2.1466004710223579e-19

R73_182 V73 V182 -1799.8886358896755
L73_182 V73 V182 1.8051377154460868e-10
C73_182 V73 V182 2.6849706495850978e-20

R73_183 V73 V183 -1410.0225217781788
L73_183 V73 V183 -2.1326964019861767e-11
C73_183 V73 V183 -1.0187488397016302e-20

R73_184 V73 V184 -945.4408751016812
L73_184 V73 V184 -1.0568719838063383e-11
C73_184 V73 V184 7.630647623004208e-20

R73_185 V73 V185 -3856.2321202271232
L73_185 V73 V185 -2.4286363292334085e-12
C73_185 V73 V185 -1.5868226265566206e-19

R73_186 V73 V186 -1768.8235446070416
L73_186 V73 V186 1.4011583877886075e-11
C73_186 V73 V186 4.376477945982513e-20

R73_187 V73 V187 2662.2553607936984
L73_187 V73 V187 -6.564674971381345e-12
C73_187 V73 V187 8.392330645011223e-20

R73_188 V73 V188 966.999367357676
L73_188 V73 V188 -1.0082213149996981e-10
C73_188 V73 V188 4.504390565758262e-20

R73_189 V73 V189 -7861.337303526974
L73_189 V73 V189 -1.651017016166329e-12
C73_189 V73 V189 -1.0886481530943217e-19

R73_190 V73 V190 3435.6937874325595
L73_190 V73 V190 -1.8872526976433136e-11
C73_190 V73 V190 -4.4792982352147993e-20

R73_191 V73 V191 1016.2147558018627
L73_191 V73 V191 -1.6176170194880384e-11
C73_191 V73 V191 -3.219228345658322e-20

R73_192 V73 V192 1368.0492883887027
L73_192 V73 V192 -7.696047492046374e-12
C73_192 V73 V192 -1.0427425336347161e-19

R73_193 V73 V193 -4051.692192629552
L73_193 V73 V193 1.3139584277742665e-12
C73_193 V73 V193 7.011737227548097e-20

R73_194 V73 V194 1309.0761222498916
L73_194 V73 V194 -1.4031065049260843e-11
C73_194 V73 V194 -1.155672205676888e-19

R73_195 V73 V195 -1588.1769272946192
L73_195 V73 V195 -6.078266784204323e-11
C73_195 V73 V195 -3.530367284048876e-20

R73_196 V73 V196 -1759.0306158028673
L73_196 V73 V196 5.550078554337501e-12
C73_196 V73 V196 7.19068084113495e-20

R73_197 V73 V197 920.8228987129825
L73_197 V73 V197 5.884922971729745e-12
C73_197 V73 V197 1.0972197668281915e-19

R73_198 V73 V198 -1105.6239232548132
L73_198 V73 V198 4.843249816094949e-12
C73_198 V73 V198 -2.896643397950915e-21

R73_199 V73 V199 -677.6462343877214
L73_199 V73 V199 3.649125114490471e-12
C73_199 V73 V199 -2.7964273535217583e-20

R73_200 V73 V200 -1344.931049152957
L73_200 V73 V200 6.633088404094466e-12
C73_200 V73 V200 5.888740341130947e-20

R74_74 V74 0 4239.915231516681
L74_74 V74 0 -8.644896830528172e-13
C74_74 V74 0 -6.022551579561107e-19

R74_75 V74 V75 -13865.404756708
L74_75 V74 V75 -9.988036755839987e-11
C74_75 V74 V75 -2.0041988130186347e-20

R74_76 V74 V76 -3267.984682430031
L74_76 V74 V76 1.970382674258162e-11
C74_76 V74 V76 7.880594689400705e-20

R74_77 V74 V77 -2114.5400062333842
L74_77 V74 V77 3.0977322118822e-12
C74_77 V74 V77 1.094921489628076e-19

R74_78 V74 V78 621.5374414335255
L74_78 V74 V78 1.3287282226558694e-12
C74_78 V74 V78 4.1726502550580422e-19

R74_79 V74 V79 2218.5933509012925
L74_79 V74 V79 1.2796423243095075e-11
C74_79 V74 V79 5.767994264625872e-20

R74_80 V74 V80 1351.6509292458065
L74_80 V74 V80 9.417196370761602e-12
C74_80 V74 V80 7.705602670713616e-20

R74_81 V74 V81 920.1348080160899
L74_81 V74 V81 6.513909351448576e-12
C74_81 V74 V81 9.611298734707682e-20

R74_82 V74 V82 -2983.8523276242104
L74_82 V74 V82 1.23519705930269e-12
C74_82 V74 V82 4.090418455371368e-19

R74_83 V74 V83 -3448.4480212564663
L74_83 V74 V83 -2.0823482337636404e-11
C74_83 V74 V83 -5.737778064765378e-20

R74_84 V74 V84 -65404.74484471501
L74_84 V74 V84 2.5217075654647415e-11
C74_84 V74 V84 6.024462486577544e-22

R74_85 V74 V85 -3913.8593355143325
L74_85 V74 V85 -6.9498076936165395e-12
C74_85 V74 V85 -6.664196170292947e-20

R74_86 V74 V86 -1223.0951671649389
L74_86 V74 V86 -1.0729941665379406e-12
C74_86 V74 V86 -5.573222452021224e-19

R74_87 V74 V87 -1949.0331571741415
L74_87 V74 V87 6.140988436982894e-12
C74_87 V74 V87 1.3400840588731938e-19

R74_88 V74 V88 -1375.5130152020968
L74_88 V74 V88 9.39123364666821e-12
C74_88 V74 V88 1.3126367864619484e-19

R74_89 V74 V89 -1473.7140263637793
L74_89 V74 V89 -2.728909211382556e-10
C74_89 V74 V89 3.711644820854514e-20

R74_90 V74 V90 1398.5732614400736
L74_90 V74 V90 -6.984209699243409e-11
C74_90 V74 V90 1.0545490195209163e-19

R74_91 V74 V91 1065.4035022437688
L74_91 V74 V91 -4.8538493288960065e-12
C74_91 V74 V91 -1.59136766884708e-19

R74_92 V74 V92 1514.630510231918
L74_92 V74 V92 -2.477852772237402e-12
C74_92 V74 V92 -2.184601421057142e-19

R74_93 V74 V93 1911.8247082295445
L74_93 V74 V93 4.182939491480945e-12
C74_93 V74 V93 4.8568917560374444e-20

R74_94 V74 V94 12112.000192251664
L74_94 V74 V94 1.9373358651917062e-12
C74_94 V74 V94 2.142080175871331e-19

R74_95 V74 V95 3201.8128686534224
L74_95 V74 V95 1.6685994523992846e-11
C74_95 V74 V95 -7.077908512454333e-20

R74_96 V74 V96 2225.364715450048
L74_96 V74 V96 4.53739292277758e-12
C74_96 V74 V96 -3.92614718448801e-20

R74_97 V74 V97 -2124.975541593304
L74_97 V74 V97 1.4207150363304606e-11
C74_97 V74 V97 -1.4694499816918632e-19

R74_98 V74 V98 -1908.265354354273
L74_98 V74 V98 -3.0219278847555915e-12
C74_98 V74 V98 -9.600750846779549e-20

R74_99 V74 V99 -861.7296459837646
L74_99 V74 V99 3.945102370612954e-12
C74_99 V74 V99 1.937717584784721e-19

R74_100 V74 V100 -1306.0303798202924
L74_100 V74 V100 2.5638757448066856e-12
C74_100 V74 V100 3.253528944215436e-19

R74_101 V74 V101 1301.725968786928
L74_101 V74 V101 -5.261418807820365e-12
C74_101 V74 V101 2.2708943207656915e-20

R74_102 V74 V102 -1747.5290579812254
L74_102 V74 V102 -3.664847088988414e-12
C74_102 V74 V102 -1.973744156178117e-19

R74_103 V74 V103 -3577.1181931934548
L74_103 V74 V103 -2.343169716474728e-12
C74_103 V74 V103 -2.0181179817006853e-19

R74_104 V74 V104 -2050.8855894088383
L74_104 V74 V104 -2.256395101492999e-12
C74_104 V74 V104 -2.0075076173076037e-19

R74_105 V74 V105 -1798.4182986154185
L74_105 V74 V105 1.666594815485069e-11
C74_105 V74 V105 2.4373033368558004e-20

R74_106 V74 V106 623.2496792661001
L74_106 V74 V106 2.5055074851945823e-12
C74_106 V74 V106 2.0237376317409528e-19

R74_107 V74 V107 840.3071922124404
L74_107 V74 V107 6.7233471623725625e-12
C74_107 V74 V107 1.8572757846462958e-20

R74_108 V74 V108 1080.1633175305192
L74_108 V74 V108 -6.036006612967884e-10
C74_108 V74 V108 -5.242141322099203e-20

R74_109 V74 V109 -985.7749205374623
L74_109 V74 V109 4.424853018529246e-12
C74_109 V74 V109 3.186601731080421e-20

R74_110 V74 V110 -5631.963612296248
L74_110 V74 V110 6.19675952940746e-12
C74_110 V74 V110 2.439053553842119e-19

R74_111 V74 V111 2297.69907631015
L74_111 V74 V111 4.548355066815606e-12
C74_111 V74 V111 7.760116271611641e-20

R74_112 V74 V112 2923.888137500501
L74_112 V74 V112 1.158557837966694e-11
C74_112 V74 V112 -3.6007339778809594e-20

R74_113 V74 V113 519.7197996129012
L74_113 V74 V113 4.779317360909863e-12
C74_113 V74 V113 8.287138444396029e-20

R74_114 V74 V114 -1052.8500220039832
L74_114 V74 V114 -1.7589579334150215e-12
C74_114 V74 V114 -4.2545869869217875e-19

R74_115 V74 V115 -618.6183355259055
L74_115 V74 V115 -5.366616175867887e-12
C74_115 V74 V115 -7.064665121686368e-20

R74_116 V74 V116 -708.6571146469997
L74_116 V74 V116 8.846106129521595e-12
C74_116 V74 V116 4.753486241579908e-20

R74_117 V74 V117 2840.0741662433334
L74_117 V74 V117 -4.6671197111908504e-12
C74_117 V74 V117 -1.8840968533729238e-19

R74_118 V74 V118 -1748.1786031651409
L74_118 V74 V118 9.882013268729774e-12
C74_118 V74 V118 7.867401950153331e-20

R74_119 V74 V119 3816.093960083441
L74_119 V74 V119 -4.229801528804423e-10
C74_119 V74 V119 8.698012576609386e-20

R74_120 V74 V120 1877.5583759591887
L74_120 V74 V120 -9.444162834729749e-12
C74_120 V74 V120 1.1645473033352192e-19

R74_121 V74 V121 -525.758621750712
L74_121 V74 V121 -6.00488221496663e-12
C74_121 V74 V121 -4.1239743997514117e-20

R74_122 V74 V122 832.8576722216362
L74_122 V74 V122 1.8361379748447545e-12
C74_122 V74 V122 3.6280950484730345e-19

R74_123 V74 V123 951.5008173772962
L74_123 V74 V123 -6.556224697498252e-12
C74_123 V74 V123 -2.0860299553110576e-19

R74_124 V74 V124 1119.6011109853591
L74_124 V74 V124 -4.0509717407739056e-12
C74_124 V74 V124 -3.3968482595341555e-19

R74_125 V74 V125 -7331.213624166754
L74_125 V74 V125 4.567216717416634e-12
C74_125 V74 V125 2.188848789402661e-19

R74_126 V74 V126 665.2078070033303
L74_126 V74 V126 -2.779232845866601e-12
C74_126 V74 V126 -2.7535222705783987e-19

R74_127 V74 V127 16831.344046211238
L74_127 V74 V127 5.756939119598015e-12
C74_127 V74 V127 1.118891011323233e-19

R74_128 V74 V128 -5626.501921163262
L74_128 V74 V128 2.724419955447707e-12
C74_128 V74 V128 1.3987223244352687e-19

R74_129 V74 V129 460.1283460029771
L74_129 V74 V129 2.0462186010039817e-12
C74_129 V74 V129 1.0391681370303111e-19

R74_130 V74 V130 -516.8693447362594
L74_130 V74 V130 -2.3775022739518996e-12
C74_130 V74 V130 -8.413381228800554e-20

R74_131 V74 V131 -1115.8306513242471
L74_131 V74 V131 1.1901911262663247e-11
C74_131 V74 V131 1.1704234662817677e-19

R74_132 V74 V132 -949.3502643338455
L74_132 V74 V132 -5.360528213588172e-11
C74_132 V74 V132 1.8579493082665823e-19

R74_133 V74 V133 -1678.2767183109647
L74_133 V74 V133 -1.8625954211193156e-12
C74_133 V74 V133 -3.136221690932102e-19

R74_134 V74 V134 5627.407229985433
L74_134 V74 V134 1.2088759689169906e-12
C74_134 V74 V134 4.524672911881108e-19

R74_135 V74 V135 -10631.561456046547
L74_135 V74 V135 -2.9761778105441863e-12
C74_135 V74 V135 -2.8751898878286196e-19

R74_136 V74 V136 -4129.799168356939
L74_136 V74 V136 -3.2637912194451317e-12
C74_136 V74 V136 -3.5614922020550535e-19

R74_137 V74 V137 -878.4441598052919
L74_137 V74 V137 -3.4505278908237985e-12
C74_137 V74 V137 -1.3656532428178208e-19

R74_138 V74 V138 1166.0469570082525
L74_138 V74 V138 -2.0743926361982967e-12
C74_138 V74 V138 -3.601070706931176e-19

R74_139 V74 V139 1516.6272212082172
L74_139 V74 V139 7.852861562979716e-12
C74_139 V74 V139 2.1065064633748156e-19

R74_140 V74 V140 667.6431850179906
L74_140 V74 V140 1.3122955715675917e-11
C74_140 V74 V140 2.372193511989287e-19

R74_141 V74 V141 -2361.3517404868353
L74_141 V74 V141 1.7128770076005446e-12
C74_141 V74 V141 3.611071738606301e-19

R74_142 V74 V142 -999.9710410107036
L74_142 V74 V142 -2.0848368625508272e-12
C74_142 V74 V142 -9.84938224318144e-21

R74_143 V74 V143 4573.800725215945
L74_143 V74 V143 4.223430608204857e-12
C74_143 V74 V143 7.610050771900071e-20

R74_144 V74 V144 -2036.4368969916138
L74_144 V74 V144 4.900508079903018e-12
C74_144 V74 V144 1.19597391758015e-19

R74_145 V74 V145 624.3286834134083
L74_145 V74 V145 5.888297361574723e-12
C74_145 V74 V145 1.0938006387167774e-19

R74_146 V74 V146 364.03959928409256
L74_146 V74 V146 2.048438770354696e-12
C74_146 V74 V146 8.235678536103134e-20

R74_147 V74 V147 -9365.028930804634
L74_147 V74 V147 -9.565462009354742e-12
C74_147 V74 V147 -1.6864409694889658e-19

R74_148 V74 V148 1039.914555682025
L74_148 V74 V148 -5.538940441385367e-12
C74_148 V74 V148 -2.113147976705532e-19

R74_149 V74 V149 1293.8946041742884
L74_149 V74 V149 -1.561726338051408e-12
C74_149 V74 V149 -3.591179467518974e-19

R74_150 V74 V150 -309.7054003040466
L74_150 V74 V150 2.0141578672400047e-11
C74_150 V74 V150 2.163434009662711e-19

R74_151 V74 V151 -3515.2484115153175
L74_151 V74 V151 -8.49765186512158e-12
C74_151 V74 V151 -2.5929050912733715e-20

R74_152 V74 V152 -982.4209375514607
L74_152 V74 V152 1.9988660353592818e-11
C74_152 V74 V152 4.0507983893551974e-20

R74_153 V74 V153 -670.9793320683449
L74_153 V74 V153 -5.367146392441651e-12
C74_153 V74 V153 -1.2175518845209114e-19

R74_154 V74 V154 -1013.5106850325051
L74_154 V74 V154 -7.570217019555426e-12
C74_154 V74 V154 -3.044777864230945e-19

R74_155 V74 V155 -858.2945541404835
L74_155 V74 V155 -2.5253104203867743e-11
C74_155 V74 V155 1.2039020142138515e-19

R74_156 V74 V156 2158.993222351894
L74_156 V74 V156 -6.4977566744661535e-12
C74_156 V74 V156 7.167998507875694e-20

R74_157 V74 V157 -407.2630433289105
L74_157 V74 V157 1.6747099587138475e-12
C74_157 V74 V157 2.2259611180464163e-19

R74_158 V74 V158 505.4686198365336
L74_158 V74 V158 -8.417377963245564e-12
C74_158 V74 V158 1.691618594172468e-19

R74_159 V74 V159 785.5579587359947
L74_159 V74 V159 -1.9472567052834233e-11
C74_159 V74 V159 -2.14934207992963e-19

R74_160 V74 V160 -10255.862963275826
L74_160 V74 V160 -1.3484134612134787e-11
C74_160 V74 V160 -1.6729334418957973e-19

R74_161 V74 V161 481.89472536464115
L74_161 V74 V161 4.02134326806454e-12
C74_161 V74 V161 2.0651030804658655e-19

R74_162 V74 V162 378.37251070564673
L74_162 V74 V162 -1.8077535898987496e-12
C74_162 V74 V162 -1.2891490973772883e-19

R74_163 V74 V163 742.4196033600316
L74_163 V74 V163 3.476898737986745e-12
C74_163 V74 V163 1.482991840291823e-19

R74_164 V74 V164 430.0528418338398
L74_164 V74 V164 4.673129333732752e-12
C74_164 V74 V164 1.1209312676833557e-19

R74_165 V74 V165 492.0178062599695
L74_165 V74 V165 -2.171479775638193e-12
C74_165 V74 V165 -2.56948906546437e-19

R74_166 V74 V166 -369.578135801979
L74_166 V74 V166 3.3053183763474515e-12
C74_166 V74 V166 -4.5256267307731536e-21

R74_167 V74 V167 14376.24197533728
L74_167 V74 V167 -5.4976862350889434e-12
C74_167 V74 V167 8.548374728305318e-20

R74_168 V74 V168 -2497.1792011136863
L74_168 V74 V168 -1.0072141204068254e-11
C74_168 V74 V168 2.108332757283533e-19

R74_169 V74 V169 -405.0529124567589
L74_169 V74 V169 -3.2188192301406563e-12
C74_169 V74 V169 -2.0011926665731324e-19

R74_170 V74 V170 -596.3573074488953
L74_170 V74 V170 2.1251139173076988e-12
C74_170 V74 V170 -7.075536752125697e-20

R74_171 V74 V171 -593.9165370211722
L74_171 V74 V171 -2.36922123901731e-12
C74_171 V74 V171 -2.253160715315311e-19

R74_172 V74 V172 -707.8913935348661
L74_172 V74 V172 -2.169325670965516e-12
C74_172 V74 V172 -2.0021687962326455e-19

R74_173 V74 V173 2415.976327126994
L74_173 V74 V173 2.5404182270826e-12
C74_173 V74 V173 1.2856245932713664e-19

R74_174 V74 V174 462.0545583038711
L74_174 V74 V174 -8.700136121756847e-13
C74_174 V74 V174 -1.934419715535514e-20

R74_175 V74 V175 3352.673993819381
L74_175 V74 V175 -1.624936187411194e-11
C74_175 V74 V175 -1.0327319328521391e-20

R74_176 V74 V176 1903.8251102272538
L74_176 V74 V176 3.82466248861615e-12
C74_176 V74 V176 1.2335128755015384e-20

R74_177 V74 V177 450.3366640952924
L74_177 V74 V177 2.9425852490285006e-12
C74_177 V74 V177 -8.486825278808423e-21

R74_178 V74 V178 557.2514906011033
L74_178 V74 V178 3.0062869722960217e-12
C74_178 V74 V178 1.4071433201754582e-19

R74_179 V74 V179 1455.8409346475266
L74_179 V74 V179 2.351993342198489e-12
C74_179 V74 V179 1.5713311363591473e-19

R74_180 V74 V180 687.0608617849747
L74_180 V74 V180 3.246123962985222e-12
C74_180 V74 V180 5.712599872801727e-20

R74_181 V74 V181 -700.5298478012395
L74_181 V74 V181 -6.01320861962705e-12
C74_181 V74 V181 1.4107942701353738e-19

R74_182 V74 V182 -264.44749158920933
L74_182 V74 V182 1.4798526777364787e-11
C74_182 V74 V182 -1.2817244794238772e-19

R74_183 V74 V183 3213.0513267831666
L74_183 V74 V183 1.301169175052857e-11
C74_183 V74 V183 1.9829250195128018e-20

R74_184 V74 V184 -2811.585344213491
L74_184 V74 V184 -6.4596232876106045e-12
C74_184 V74 V184 5.825128395382273e-20

R74_185 V74 V185 -674.7454612259884
L74_185 V74 V185 -3.0677548198368886e-12
C74_185 V74 V185 -7.325363674776482e-20

R74_186 V74 V186 -777.8964541027924
L74_186 V74 V186 -1.855781221289535e-12
C74_186 V74 V186 3.523388209395545e-20

R74_187 V74 V187 -3203.066435106149
L74_187 V74 V187 -2.112649434805654e-12
C74_187 V74 V187 -1.5536078618748945e-20

R74_188 V74 V188 -936.1251845606691
L74_188 V74 V188 -9.63569746846076e-12
C74_188 V74 V188 -1.7281070453983213e-20

R74_189 V74 V189 520.3888783864528
L74_189 V74 V189 -8.520693517788369e-12
C74_189 V74 V189 -2.559305641214082e-19

R74_190 V74 V190 318.07077506788727
L74_190 V74 V190 4.795939101265342e-12
C74_190 V74 V190 1.5278863238301097e-19

R74_191 V74 V191 -11482.650186944566
L74_191 V74 V191 -2.761668332253802e-12
C74_191 V74 V191 -2.4866850773734126e-19

R74_192 V74 V192 1231.9579207966926
L74_192 V74 V192 -2.7159830436638745e-12
C74_192 V74 V192 -3.123958640039924e-19

R74_193 V74 V193 2677.677904283077
L74_193 V74 V193 2.353408781382849e-12
C74_193 V74 V193 5.617620846443082e-20

R74_194 V74 V194 -648.6987735871559
L74_194 V74 V194 -2.201386304497816e-12
C74_194 V74 V194 -2.1645592660681012e-19

R74_195 V74 V195 4449.7159988304775
L74_195 V74 V195 1.8873217273494735e-12
C74_195 V74 V195 3.0841676261329667e-19

R74_196 V74 V196 2119.6057829521956
L74_196 V74 V196 1.4646413111093859e-12
C74_196 V74 V196 4.170322411922842e-19

R74_197 V74 V197 -884.2839439676882
L74_197 V74 V197 2.092488044959714e-12
C74_197 V74 V197 3.0502727701859304e-19

R74_198 V74 V198 -357.2075286370849
L74_198 V74 V198 1.896151456154839e-11
C74_198 V74 V198 -6.076832823375591e-20

R74_199 V74 V199 -3739.9765025883153
L74_199 V74 V199 1.7882490612763447e-12
C74_199 V74 V199 1.2675666002977175e-19

R74_200 V74 V200 -3209.1516251899175
L74_200 V74 V200 3.2640806427743935e-12
C74_200 V74 V200 1.504033349826062e-19

R75_75 V75 0 331.70733296412226
L75_75 V75 0 -9.264319954717147e-13
C75_75 V75 0 3.459440039273888e-19

R75_76 V75 V76 -9861.727791556597
L75_76 V75 V76 -1.4772083360570344e-11
C75_76 V75 V76 6.18951863722743e-20

R75_77 V75 V77 -3798.419447059843
L75_77 V75 V77 3.248516585805867e-12
C75_77 V75 V77 1.499842963223606e-19

R75_78 V75 V78 4321.936524724728
L75_78 V75 V78 8.788604476532351e-11
C75_78 V75 V78 5.4193967037515335e-20

R75_79 V75 V79 2031.2189670763755
L75_79 V75 V79 2.22403379264551e-12
C75_79 V75 V79 1.5707517679114712e-19

R75_80 V75 V80 4220.715443847259
L75_80 V75 V80 3.078757914446246e-11
C75_80 V75 V80 1.5076512500004924e-20

R75_81 V75 V81 -11639.155171836745
L75_81 V75 V81 9.312309764160376e-12
C75_81 V75 V81 2.891065162869984e-20

R75_82 V75 V82 -17149.511897049008
L75_82 V75 V82 1.49440162907415e-11
C75_82 V75 V82 -1.5712210853177058e-20

R75_83 V75 V83 3141.660381794631
L75_83 V75 V83 7.634441254873182e-13
C75_83 V75 V83 7.56529077427443e-19

R75_84 V75 V84 6609.144017704326
L75_84 V75 V84 5.742318399662769e-12
C75_84 V75 V84 5.770481820261819e-20

R75_85 V75 V85 6628.134341130663
L75_85 V75 V85 2.958413650220134e-11
C75_85 V75 V85 -1.505459554285978e-20

R75_86 V75 V86 -3508.576356621114
L75_86 V75 V86 5.272134200422667e-12
C75_86 V75 V86 7.103782185556174e-20

R75_87 V75 V87 -2162.765267758497
L75_87 V75 V87 -7.28450440534365e-13
C75_87 V75 V87 -7.126690518608394e-19

R75_88 V75 V88 -1588.738856933418
L75_88 V75 V88 1.3612104978411167e-11
C75_88 V75 V88 1.0773880788182504e-19

R75_89 V75 V89 5616.368947140996
L75_89 V75 V89 1.1913669766827313e-10
C75_89 V75 V89 2.714703657511548e-20

R75_90 V75 V90 4450.511371092401
L75_90 V75 V90 -2.3255960971371867e-12
C75_90 V75 V90 -8.80014892919246e-20

R75_91 V75 V91 983.8374873786298
L75_91 V75 V91 7.487178501446401e-13
C75_91 V75 V91 5.2304143970498e-19

R75_92 V75 V92 1440.9630818253754
L75_92 V75 V92 -4.347886343396163e-12
C75_92 V75 V92 -1.648733020458055e-19

R75_93 V75 V93 -1508.2763280918036
L75_93 V75 V93 -1.8872319151933284e-11
C75_93 V75 V93 -7.17085390800247e-20

R75_94 V75 V94 14883.205444290683
L75_94 V75 V94 -9.496589766091608e-12
C75_94 V75 V94 -1.1805615245919007e-19

R75_95 V75 V95 -2784.727614154737
L75_95 V75 V95 3.5792951642191628e-12
C75_95 V75 V95 2.5995050429100067e-19

R75_96 V75 V96 2060.738854796933
L75_96 V75 V96 9.274050569956575e-11
C75_96 V75 V96 -5.682650636332316e-20

R75_97 V75 V97 3497717.5620614737
L75_97 V75 V97 3.76432982104611e-12
C75_97 V75 V97 1.9136936257693052e-20

R75_98 V75 V98 11097.35349212544
L75_98 V75 V98 2.174152245431867e-12
C75_98 V75 V98 1.423119424707248e-19

R75_99 V75 V99 -1825.9346459469887
L75_99 V75 V99 -5.917729442373481e-13
C75_99 V75 V99 -7.649256375708215e-19

R75_100 V75 V100 -1050.778492237015
L75_100 V75 V100 6.2798577943184585e-12
C75_100 V75 V100 2.2768525107551567e-19

R75_101 V75 V101 919.0824684229855
L75_101 V75 V101 -5.508477679084411e-12
C75_101 V75 V101 -4.081354829897161e-20

R75_102 V75 V102 -4260.267061890466
L75_102 V75 V102 -1.3798210594850797e-10
C75_102 V75 V102 8.567574041384074e-20

R75_103 V75 V103 -5164.009987789875
L75_103 V75 V103 1.209272579908581e-12
C75_103 V75 V103 2.556840462517677e-19

R75_104 V75 V104 -4746.826663918745
L75_104 V75 V104 1.9750501676948245e-11
C75_104 V75 V104 -1.4089374854880502e-20

R75_105 V75 V105 -761.1184336899431
L75_105 V75 V105 6.129209953027021e-12
C75_105 V75 V105 2.1593969489492438e-20

R75_106 V75 V106 -3241.788344423987
L75_106 V75 V106 -1.5166214403297088e-12
C75_106 V75 V106 -2.978011945514925e-19

R75_107 V75 V107 766.1999795947263
L75_107 V75 V107 1.6707257292342023e-12
C75_107 V75 V107 3.205038688651185e-19

R75_108 V75 V108 970.0397418808344
L75_108 V75 V108 -5.338541735719337e-12
C75_108 V75 V108 -1.284876046713402e-19

R75_109 V75 V109 -1560.890006412065
L75_109 V75 V109 5.654437816947453e-12
C75_109 V75 V109 9.18760821177401e-20

R75_110 V75 V110 1151.2948426194364
L75_110 V75 V110 4.176677363455676e-12
C75_110 V75 V110 8.358362164385053e-20

R75_111 V75 V111 2351.1335346066694
L75_111 V75 V111 -2.7884932513314742e-12
C75_111 V75 V111 -2.6818754547272632e-21

R75_112 V75 V112 -6139.385097159343
L75_112 V75 V112 -3.281289568840658e-12
C75_112 V75 V112 -2.0194583979301344e-19

R75_113 V75 V113 544.1285093947159
L75_113 V75 V113 -1.045589043372726e-11
C75_113 V75 V113 -8.674758215767586e-20

R75_114 V75 V114 46888.70035842859
L75_114 V75 V114 1.9579732290832642e-12
C75_114 V75 V114 2.400659186867419e-19

R75_115 V75 V115 -474.75198501575903
L75_115 V75 V115 -1.084365847692674e-12
C75_115 V75 V115 -2.936759184600896e-19

R75_116 V75 V116 -1038.9457702130853
L75_116 V75 V116 2.3447518650213515e-12
C75_116 V75 V116 2.5022038953131125e-19

R75_117 V75 V117 4679.361444778432
L75_117 V75 V117 -6.017049396013608e-12
C75_117 V75 V117 -9.680621313079977e-20

R75_118 V75 V118 -860.1534123379594
L75_118 V75 V118 -4.415370443594139e-12
C75_118 V75 V118 -6.249078426177577e-20

R75_119 V75 V119 541.7294143327057
L75_119 V75 V119 1.2925487469924927e-12
C75_119 V75 V119 1.5460504922358964e-20

R75_120 V75 V120 1868.5838298692847
L75_120 V75 V120 -6.153976069386286e-12
C75_120 V75 V120 4.3094815848505366e-20

R75_121 V75 V121 -541.026297705543
L75_121 V75 V121 3.2485402167420887e-12
C75_121 V75 V121 1.951264489641182e-19

R75_122 V75 V122 2122.224355319842
L75_122 V75 V122 -3.4340811815412673e-12
C75_122 V75 V122 -1.633639597953631e-19

R75_123 V75 V123 -53301.691261985885
L75_123 V75 V123 1.203443284514125e-12
C75_123 V75 V123 6.432925372647909e-19

R75_124 V75 V124 3817.6910351658066
L75_124 V75 V124 -3.1763068544623236e-12
C75_124 V75 V124 -3.771584736248188e-19

R75_125 V75 V125 -2098.0820647184605
L75_125 V75 V125 7.964055571733042e-12
C75_125 V75 V125 1.4256572766390155e-20

R75_126 V75 V126 694.4069475955426
L75_126 V75 V126 3.695031222809886e-12
C75_126 V75 V126 9.414691634968798e-20

R75_127 V75 V127 -1323.619296525171
L75_127 V75 V127 -7.386953731780187e-13
C75_127 V75 V127 -4.358241724281378e-19

R75_128 V75 V128 6252.382202713886
L75_128 V75 V128 3.499290651056384e-12
C75_128 V75 V128 1.987125479650065e-19

R75_129 V75 V129 510.4710288069325
L75_129 V75 V129 -3.776185202893616e-12
C75_129 V75 V129 -1.5066147718683038e-19

R75_130 V75 V130 -1012.5335558707509
L75_130 V75 V130 5.885345104174546e-12
C75_130 V75 V130 1.5285590922324316e-19

R75_131 V75 V131 2067.697151293344
L75_131 V75 V131 2.9461781429785323e-12
C75_131 V75 V131 -1.355914094355057e-19

R75_132 V75 V132 -2082.229611144934
L75_132 V75 V132 -1.5514876762149386e-11
C75_132 V75 V132 -5.2637417211833694e-20

R75_133 V75 V133 2973.9374466148074
L75_133 V75 V133 7.404901224598806e-12
C75_133 V75 V133 9.338395292240177e-20

R75_134 V75 V134 -1683.9295134075949
L75_134 V75 V134 -5.9132094512839314e-12
C75_134 V75 V134 -1.8282465298733577e-19

R75_135 V75 V135 -634.7271686922206
L75_135 V75 V135 9.059143190706422e-13
C75_135 V75 V135 8.641223214472673e-19

R75_136 V75 V136 -1137.5603459490305
L75_136 V75 V136 -6.616742290908752e-12
C75_136 V75 V136 -3.5778695868758803e-19

R75_137 V75 V137 -411.85654032751495
L75_137 V75 V137 5.207249481991881e-12
C75_137 V75 V137 5.53868883794545e-20

R75_138 V75 V138 1961.5865654524714
L75_138 V75 V138 7.124385134882952e-12
C75_138 V75 V138 1.5081296711837598e-19

R75_139 V75 V139 505.33108188860604
L75_139 V75 V139 -7.427376156298742e-13
C75_139 V75 V139 -9.765091933590063e-19

R75_140 V75 V140 852.5883394776151
L75_140 V75 V140 -2.2555616351382205e-11
C75_140 V75 V140 3.8478262970903745e-19

R75_141 V75 V141 -3941.007234869681
L75_141 V75 V141 -1.7381606163094008e-11
C75_141 V75 V141 -6.510643258449166e-20

R75_142 V75 V142 793.6897355822159
L75_142 V75 V142 -6.253117180851452e-12
C75_142 V75 V142 5.736411728352962e-20

R75_143 V75 V143 593.2130892781171
L75_143 V75 V143 4.39746886397461e-12
C75_143 V75 V143 1.0385167672419225e-19

R75_144 V75 V144 641.1568492222747
L75_144 V75 V144 6.569210440051528e-12
C75_144 V75 V144 -3.3373867727709507e-20

R75_145 V75 V145 376.57388258968206
L75_145 V75 V145 -1.1264223310187673e-11
C75_145 V75 V145 1.4320052799744576e-20

R75_146 V75 V146 12968.805926744755
L75_146 V75 V146 1.6475855831534422e-11
C75_146 V75 V146 -9.538046051082874e-20

R75_147 V75 V147 -272.0760472299728
L75_147 V75 V147 7.313439234860648e-12
C75_147 V75 V147 5.106821304000764e-19

R75_148 V75 V148 -465.39237226751266
L75_148 V75 V148 -2.9064779971087202e-12
C75_148 V75 V148 -2.477199951374219e-19

R75_149 V75 V149 2478.451827609495
L75_149 V75 V149 1.1086055633646962e-11
C75_149 V75 V149 5.002251028500966e-20

R75_150 V75 V150 -433.3693166931828
L75_150 V75 V150 4.0501081026785854e-12
C75_150 V75 V150 -1.593475386075104e-19

R75_151 V75 V151 945.1192009524996
L75_151 V75 V151 6.153883764687714e-12
C75_151 V75 V151 -1.3929937619640551e-19

R75_152 V75 V152 1486.7382811203724
L75_152 V75 V152 5.808880641345095e-12
C75_152 V75 V152 1.0659711795146996e-19

R75_153 V75 V153 -387.73391414267064
L75_153 V75 V153 5.925884182718416e-12
C75_153 V75 V153 6.810848167721157e-20

R75_154 V75 V154 -5941.076333198336
L75_154 V75 V154 -1.5499576793595324e-11
C75_154 V75 V154 1.7402733755890109e-19

R75_155 V75 V155 -299.75989274989917
L75_155 V75 V155 -2.1521945921869998e-12
C75_155 V75 V155 -4.384346197827386e-19

R75_156 V75 V156 -958.2456206639308
L75_156 V75 V156 -4.754265955267818e-12
C75_156 V75 V156 1.7712668654999362e-19

R75_157 V75 V157 -504.89972238261714
L75_157 V75 V157 -9.464081165741489e-12
C75_157 V75 V157 -2.555303037278465e-19

R75_158 V75 V158 803.7426933369607
L75_158 V75 V158 -5.278479579946503e-12
C75_158 V75 V158 -8.760253157278607e-20

R75_159 V75 V159 389.7887302432351
L75_159 V75 V159 2.7388151224855025e-12
C75_159 V75 V159 4.2207134799754723e-19

R75_160 V75 V160 1091.8520067411484
L75_160 V75 V160 4.843865075556948e-12
C75_160 V75 V160 -1.18698801958573e-19

R75_161 V75 V161 528.9166466887324
L75_161 V75 V161 -4.359107797801573e-12
C75_161 V75 V161 -3.4561094315695186e-20

R75_162 V75 V162 1117.22031593024
L75_162 V75 V162 -2.6565445996576845e-11
C75_162 V75 V162 -9.051666410237478e-20

R75_163 V75 V163 668.0753777631729
L75_163 V75 V163 -1.023309866920781e-12
C75_163 V75 V163 -3.5132265733342363e-19

R75_164 V75 V164 1238.8301438975482
L75_164 V75 V164 -1.0423079622215711e-11
C75_164 V75 V164 9.635657866318155e-21

R75_165 V75 V165 1200.4223641041083
L75_165 V75 V165 2.251542936733606e-12
C75_165 V75 V165 2.1110999206211353e-19

R75_166 V75 V166 -491.20690839140224
L75_166 V75 V166 -1.0451241426592942e-11
C75_166 V75 V166 1.5351476837131085e-20

R75_167 V75 V167 -750.7465706597054
L75_167 V75 V167 1.070434591675612e-12
C75_167 V75 V167 4.570728131462423e-20

R75_168 V75 V168 2545.8727786847962
L75_168 V75 V168 -2.330494047682426e-12
C75_168 V75 V168 -6.423219442156876e-20

R75_169 V75 V169 -601.9908256154188
L75_169 V75 V169 7.183833377678213e-12
C75_169 V75 V169 3.7667311860424975e-20

R75_170 V75 V170 1378.1305990408102
L75_170 V75 V170 1.6123098452314217e-11
C75_170 V75 V170 7.3755940664928e-20

R75_171 V75 V171 -486.2267586191364
L75_171 V75 V171 2.0596920133292223e-12
C75_171 V75 V171 2.279047167057064e-19

R75_172 V75 V172 -1338.32012220745
L75_172 V75 V172 5.272504594670211e-12
C75_172 V75 V172 1.4612269700160647e-19

R75_173 V75 V173 -3287.1295480405342
L75_173 V75 V173 -1.6407266797071534e-12
C75_173 V75 V173 -2.0009161134676657e-19

R75_174 V75 V174 1063.0860440577708
L75_174 V75 V174 7.877426661441853e-12
C75_174 V75 V174 -8.762009604196512e-20

R75_175 V75 V175 519.4398421575843
L75_175 V75 V175 -5.426150059110239e-13
C75_175 V75 V175 -3.8342651222653084e-19

R75_176 V75 V176 -3839.326018146084
L75_176 V75 V176 7.46425303861107e-12
C75_176 V75 V176 1.0790588214847633e-19

R75_177 V75 V177 695.9518228441567
L75_177 V75 V177 1.858456308875432e-12
C75_177 V75 V177 9.773038930141946e-20

R75_178 V75 V178 -1636.987101444002
L75_178 V75 V178 -1.8701247131271366e-11
C75_178 V75 V178 -3.168535748634513e-20

R75_179 V75 V179 -1434.4325241087824
L75_179 V75 V179 1.8026222206278407e-12
C75_179 V75 V179 1.3157837422607849e-19

R75_180 V75 V180 1484.275338271275
L75_180 V75 V180 -7.00931430467046e-12
C75_180 V75 V180 -1.7229515998818863e-19

R75_181 V75 V181 -1626.13094579019
L75_181 V75 V181 4.599523230193444e-11
C75_181 V75 V181 3.802487631065156e-20

R75_182 V75 V182 -864.5759514668308
L75_182 V75 V182 -1.778276971416431e-11
C75_182 V75 V182 2.1218424419765954e-20

R75_183 V75 V183 1716.682099314387
L75_183 V75 V183 1.1807951120584188e-12
C75_183 V75 V183 -7.05307599804685e-20

R75_184 V75 V184 62758.405532852485
L75_184 V75 V184 4.0031478448235945e-12
C75_184 V75 V184 1.169974554794081e-19

R75_185 V75 V185 -703.3455062743689
L75_185 V75 V185 -1.6471782952314426e-12
C75_185 V75 V185 -9.549186867624218e-20

R75_186 V75 V186 1389.4331354521737
L75_186 V75 V186 2.556480135398296e-12
C75_186 V75 V186 1.5288756847075875e-19

R75_187 V75 V187 -4274.790704713272
L75_187 V75 V187 -8.441915606746992e-13
C75_187 V75 V187 -1.4591717958403058e-19

R75_188 V75 V188 -3246.3100029693237
L75_188 V75 V188 1.2425268003627759e-11
C75_188 V75 V188 1.4348809290162153e-20

R75_189 V75 V189 851.0937284643092
L75_189 V75 V189 4.33828953599839e-12
C75_189 V75 V189 1.4563348077030767e-19

R75_190 V75 V190 4847.386890377808
L75_190 V75 V190 -4.294555792755191e-11
C75_190 V75 V190 -1.1636476098151704e-19

R75_191 V75 V191 -1754.6558145935446
L75_191 V75 V191 -2.1354460368117802e-11
C75_191 V75 V191 4.2922713632309806e-19

R75_192 V75 V192 -3264.654994750656
L75_192 V75 V192 -1.7913638955979855e-12
C75_192 V75 V192 -1.564347282515051e-20

R75_193 V75 V193 1095.4264360431862
L75_193 V75 V193 2.4217957163663343e-12
C75_193 V75 V193 -8.011525464768046e-20

R75_194 V75 V194 -838.4408436210432
L75_194 V75 V194 -4.2341699560060125e-12
C75_194 V75 V194 -1.618175723330557e-20

R75_195 V75 V195 3330.2944992704065
L75_195 V75 V195 -2.531151420872447e-12
C75_195 V75 V195 -7.358281158725351e-19

R75_196 V75 V196 1504.5355619753448
L75_196 V75 V196 1.7526229837227338e-12
C75_196 V75 V196 2.406537793413198e-19

R75_197 V75 V197 -1708.4001532630734
L75_197 V75 V197 -4.627277683061373e-12
C75_197 V75 V197 5.272235381867607e-22

R75_198 V75 V198 -30677.844172760706
L75_198 V75 V198 1.5066250449560442e-11
C75_198 V75 V198 -3.115511413809475e-20

R75_199 V75 V199 -1450.9329235279176
L75_199 V75 V199 2.6031947468105255e-12
C75_199 V75 V199 -1.4514892301152135e-19

R75_200 V75 V200 1061.4552986245542
L75_200 V75 V200 1.2314263558130261e-11
C75_200 V75 V200 -1.3593128174384005e-19

R76_76 V76 0 -207.76749649361423
L76_76 V76 0 -1.4668582358326278e-13
C76_76 V76 0 -2.520535903179891e-18

R76_77 V76 V77 -2322.7297940998474
L76_77 V76 V77 3.64153856897876e-12
C76_77 V76 V77 2.2297825163695264e-19

R76_78 V76 V78 1695.5777172445041
L76_78 V76 V78 -8.31891187313455e-11
C76_78 V76 V78 1.207702077002581e-20

R76_79 V76 V79 -4694.882652188694
L76_79 V76 V79 -4.999096492917317e-12
C76_79 V76 V79 -1.9830693308493418e-20

R76_80 V76 V80 952.4443904430303
L76_80 V76 V80 8.542279656939615e-13
C76_80 V76 V80 3.402300884075797e-19

R76_81 V76 V81 2790.7355410309056
L76_81 V76 V81 2.8108293205532435e-12
C76_81 V76 V81 1.380230867379588e-19

R76_82 V76 V82 -7351.106336210056
L76_82 V76 V82 3.457779883461997e-12
C76_82 V76 V82 1.5904058126529735e-19

R76_83 V76 V83 2887.845930706116
L76_83 V76 V83 7.220755281068489e-12
C76_83 V76 V83 1.0707027291041005e-19

R76_84 V76 V84 1418.7109757858598
L76_84 V76 V84 6.095942006794272e-13
C76_84 V76 V84 9.077404740550548e-19

R76_85 V76 V85 7548.999052758795
L76_85 V76 V85 4.2743844553648555e-12
C76_85 V76 V85 7.477392959152212e-20

R76_86 V76 V86 -6916.8247802851265
L76_86 V76 V86 3.031221726841182e-12
C76_86 V76 V86 1.7521677493579728e-19

R76_87 V76 V87 -2911.7525216727117
L76_87 V76 V87 -4.712743006748405e-12
C76_87 V76 V87 -6.799629986720164e-20

R76_88 V76 V88 -3196.4220536267985
L76_88 V76 V88 -5.031673113984693e-13
C76_88 V76 V88 -9.410371785549996e-19

R76_89 V76 V89 53922.0571256563
L76_89 V76 V89 -1.933273225598287e-12
C76_89 V76 V89 -2.2223937740569257e-19

R76_90 V76 V90 17609.99199456859
L76_90 V76 V90 -7.927406578110987e-13
C76_90 V76 V90 -4.552042405623595e-19

R76_91 V76 V91 1081.7297283912844
L76_91 V76 V91 2.257937955176104e-12
C76_91 V76 V91 1.3912650403056027e-19

R76_92 V76 V92 1158.445024682683
L76_92 V76 V92 5.136016875774918e-13
C76_92 V76 V92 6.200767778432557e-19

R76_93 V76 V93 -2483.1675400108134
L76_93 V76 V93 -9.203002903060135e-12
C76_93 V76 V93 -5.681517760827936e-20

R76_94 V76 V94 -42454.72969187865
L76_94 V76 V94 6.453125605427172e-12
C76_94 V76 V94 8.843691956789411e-20

R76_95 V76 V95 -6568.465756724068
L76_95 V76 V95 7.498200471507131e-11
C76_95 V76 V95 4.032591432954527e-21

R76_96 V76 V96 -570.5093232579036
L76_96 V76 V96 -9.033751753609578e-12
C76_96 V76 V96 3.060702019005918e-19

R76_97 V76 V97 -2695.8268184381527
L76_97 V76 V97 1.1736771695565795e-12
C76_97 V76 V97 4.1967149130883053e-19

R76_98 V76 V98 2205.8740173258475
L76_98 V76 V98 9.38329829011712e-13
C76_98 V76 V98 4.1034461103517174e-19

R76_99 V76 V99 -1525.0757076999855
L76_99 V76 V99 -1.3899832608839986e-12
C76_99 V76 V99 -1.2745567390880489e-19

R76_100 V76 V100 914.542250105163
L76_100 V76 V100 -6.25166761821878e-13
C76_100 V76 V100 -9.542694432021433e-19

R76_101 V76 V101 701.9423018932688
L76_101 V76 V101 -2.337506719638329e-12
C76_101 V76 V101 -1.2449454367539987e-19

R76_102 V76 V102 -2049.479264546108
L76_102 V76 V102 -2.233323440276937e-12
C76_102 V76 V102 -1.5421840224549922e-19

R76_103 V76 V103 8357.315070658378
L76_103 V76 V103 4.293253517727159e-12
C76_103 V76 V103 9.688563867793665e-20

R76_104 V76 V104 -3842.01261222939
L76_104 V76 V104 9.822291325772475e-13
C76_104 V76 V104 3.416706776965556e-19

R76_105 V76 V105 -1076.2171058195966
L76_105 V76 V105 4.3919913155329355e-10
C76_105 V76 V105 -1.0489380232217649e-19

R76_106 V76 V106 2169.621485193074
L76_106 V76 V106 -1.2143014343810327e-12
C76_106 V76 V106 -3.846888921985192e-19

R76_107 V76 V107 1015.5767908383181
L76_107 V76 V107 3.225397239533658e-12
C76_107 V76 V107 9.912372213785845e-20

R76_108 V76 V108 2362.8781553760405
L76_108 V76 V108 4.719784682063348e-12
C76_108 V76 V108 3.09352786055228e-19

R76_109 V76 V109 -727.7882153727129
L76_109 V76 V109 1.9175496399122895e-12
C76_109 V76 V109 3.9268790056012306e-19

R76_110 V76 V110 11712.99190406728
L76_110 V76 V110 3.240985168893488e-12
C76_110 V76 V110 1.0807589482300808e-19

R76_111 V76 V111 1913.1260460503397
L76_111 V76 V111 -1.3612202208493113e-11
C76_111 V76 V111 -1.1002752428370374e-19

R76_112 V76 V112 690.3658263966506
L76_112 V76 V112 2.7835153265419814e-12
C76_112 V76 V112 2.1634378266199488e-19

R76_113 V76 V113 455.1874766486945
L76_113 V76 V113 4.4618115199075426e-11
C76_113 V76 V113 -1.0692610412113974e-19

R76_114 V76 V114 -1895.2518868271713
L76_114 V76 V114 1.2102642982975858e-12
C76_114 V76 V114 3.743230524362405e-19

R76_115 V76 V115 -462.2700002710598
L76_115 V76 V115 -5.81672535914543e-12
C76_115 V76 V115 2.881771041711061e-20

R76_116 V76 V116 -310.7658250885584
L76_116 V76 V116 -7.351712522245436e-13
C76_116 V76 V116 -4.219976754916704e-19

R76_117 V76 V117 -11160.570548128397
L76_117 V76 V117 -1.6956813020660325e-12
C76_117 V76 V117 -2.9202556887471724e-19

R76_118 V76 V118 -16874.460146846148
L76_118 V76 V118 -1.834908343592781e-12
C76_118 V76 V118 -2.942224007923192e-19

R76_119 V76 V119 1294.5660091408347
L76_119 V76 V119 -2.995032789438462e-12
C76_119 V76 V119 -2.257921259311386e-19

R76_120 V76 V120 301.8937986310921
L76_120 V76 V120 2.560265490319761e-12
C76_120 V76 V120 -4.065627477873576e-19

R76_121 V76 V121 -501.31380723715404
L76_121 V76 V121 2.323333102630331e-12
C76_121 V76 V121 3.3629503910544315e-19

R76_122 V76 V122 2295.810002930005
L76_122 V76 V122 -4.815115298879318e-12
C76_122 V76 V122 -1.6100197496800963e-19

R76_123 V76 V123 878.4166487176927
L76_123 V76 V123 3.652241909709958e-12
C76_123 V76 V123 -8.924981029092876e-22

R76_124 V76 V124 -4251.768975899094
L76_124 V76 V124 5.56922625977572e-13
C76_124 V76 V124 1.1984547039956195e-18

R76_125 V76 V125 1351.997090319621
L76_125 V76 V125 1.8453967113416514e-12
C76_125 V76 V125 7.515005166895702e-20

R76_126 V76 V126 700.9765434606605
L76_126 V76 V126 1.287951602584252e-12
C76_126 V76 V126 1.8464127093248166e-19

R76_127 V76 V127 -2673.576134810083
L76_127 V76 V127 1.4557446563687558e-12
C76_127 V76 V127 3.1674173446346305e-19

R76_128 V76 V128 -492.1184243023016
L76_128 V76 V128 -8.24624961337029e-13
C76_128 V76 V128 -1.9838527940138045e-19

R76_129 V76 V129 1322.1661937534934
L76_129 V76 V129 -4.6510761374383534e-12
C76_129 V76 V129 2.6129301034258624e-20

R76_130 V76 V130 -606.8184188698455
L76_130 V76 V130 -2.650880353830391e-12
C76_130 V76 V130 -6.091510083228444e-20

R76_131 V76 V131 -17635.401403724907
L76_131 V76 V131 -1.9457391995254395e-12
C76_131 V76 V131 -2.2639223303304554e-19

R76_132 V76 V132 517.255837412493
L76_132 V76 V132 -3.165899578162203e-12
C76_132 V76 V132 -7.284169909793014e-19

R76_133 V76 V133 27320.309259383383
L76_133 V76 V133 -2.901003766243191e-12
C76_133 V76 V133 -3.385536012453707e-19

R76_134 V76 V134 5090.107875390366
L76_134 V76 V134 -4.987492455033538e-12
C76_134 V76 V134 -3.684916224261182e-19

R76_135 V76 V135 -1650.4457770080337
L76_135 V76 V135 -3.074520261387633e-12
C76_135 V76 V135 -3.1572039138107674e-19

R76_136 V76 V136 -743.157211534827
L76_136 V76 V136 6.944366257257814e-13
C76_136 V76 V136 9.851700983623219e-19

R76_137 V76 V137 -625.2643147097871
L76_137 V76 V137 1.2328356703518577e-10
C76_137 V76 V137 6.623024151351786e-20

R76_138 V76 V138 36864.79546983873
L76_138 V76 V138 2.5030893265019047e-12
C76_138 V76 V138 3.0224612064993765e-19

R76_139 V76 V139 -10563.827552156856
L76_139 V76 V139 4.2530613912299844e-12
C76_139 V76 V139 3.2306260593497974e-19

R76_140 V76 V140 525.2501405981229
L76_140 V76 V140 -7.348380337805827e-13
C76_140 V76 V140 -1.0100716537640964e-18

R76_141 V76 V141 3791.3760329038164
L76_141 V76 V141 1.2184392263318724e-12
C76_141 V76 V141 3.676484231009416e-19

R76_142 V76 V142 1765.697843023126
L76_142 V76 V142 -9.927380215473896e-12
C76_142 V76 V142 1.0701524423434043e-19

R76_143 V76 V143 614.1278658432706
L76_143 V76 V143 2.7477722965322874e-12
C76_143 V76 V143 -3.924858303852016e-21

R76_144 V76 V144 -1293.0657576579647
L76_144 V76 V144 -2.2293108719822278e-11
C76_144 V76 V144 1.1741252357525241e-19

R76_145 V76 V145 623.6452977487603
L76_145 V76 V145 5.852474135942736e-12
C76_145 V76 V145 -1.0996262905094549e-20

R76_146 V76 V146 2327.2628149284046
L76_146 V76 V146 -4.284870680436582e-12
C76_146 V76 V146 -2.195083849131914e-19

R76_147 V76 V147 -708.8281653078373
L76_147 V76 V147 5.954401871107699e-12
C76_147 V76 V147 5.9374478049564e-20

R76_148 V76 V148 441.44433969702976
L76_148 V76 V148 5.892290510157207e-13
C76_148 V76 V148 8.161197544142718e-19

R76_149 V76 V149 3170.4910583456513
L76_149 V76 V149 -9.317782439089575e-13
C76_149 V76 V149 -1.8770055296843812e-19

R76_150 V76 V150 -965.6813886342084
L76_150 V76 V150 2.260377419388762e-12
C76_150 V76 V150 2.2028041429477398e-19

R76_151 V76 V151 -3869.1875471685325
L76_151 V76 V151 -2.969262916728213e-12
C76_151 V76 V151 5.464179572837899e-20

R76_152 V76 V152 -421.1808544021914
L76_152 V76 V152 -8.757276784126464e-13
C76_152 V76 V152 -2.9958337588550995e-19

R76_153 V76 V153 -325.24703423907874
L76_153 V76 V153 -2.1206358970153047e-12
C76_153 V76 V153 -1.5630093806440818e-19

R76_154 V76 V154 -494.4307124887446
L76_154 V76 V154 -1.9923899260600886e-12
C76_154 V76 V154 2.0620742179273806e-21

R76_155 V76 V155 -428.42032955900015
L76_155 V76 V155 -2.032904363073408e-12
C76_155 V76 V155 -2.9855587621712487e-20

R76_156 V76 V156 690.5983798807422
L76_156 V76 V156 1.7865671947632653e-12
C76_156 V76 V156 -5.205184738077281e-19

R76_157 V76 V157 -1728.8883851068058
L76_157 V76 V157 7.052441086023383e-13
C76_157 V76 V157 3.5744400951799563e-19

R76_158 V76 V158 390.27044378701856
L76_158 V76 V158 7.503214668596307e-11
C76_158 V76 V158 -6.270317780819557e-20

R76_159 V76 V159 437.40597861236904
L76_159 V76 V159 3.3227563955509475e-12
C76_159 V76 V159 -1.1252287369464588e-19

R76_160 V76 V160 -1912.6850904334376
L76_160 V76 V160 6.616825024999991e-12
C76_160 V76 V160 3.314446486201147e-19

R76_161 V76 V161 989.6275698628331
L76_161 V76 V161 -1.8239562350699006e-12
C76_161 V76 V161 -2.2120190211825137e-20

R76_162 V76 V162 1116.6403278327375
L76_162 V76 V162 -3.0685717962746737e-12
C76_162 V76 V162 -8.988205192901486e-20

R76_163 V76 V163 648.1153420003008
L76_163 V76 V163 7.314621902046554e-12
C76_163 V76 V163 6.412238565783529e-20

R76_164 V76 V164 181.7826826601053
L76_164 V76 V164 -1.1560597943586025e-12
C76_164 V76 V164 -2.591576576980222e-19

R76_165 V76 V165 449.1780878685805
L76_165 V76 V165 1.7420363074451805e-12
C76_165 V76 V165 1.398436268478423e-19

R76_166 V76 V166 -880.7335915923047
L76_166 V76 V166 2.9007117075799885e-12
C76_166 V76 V166 2.796008047119235e-19

R76_167 V76 V167 1205.569834602124
L76_167 V76 V167 -2.312135943545078e-12
C76_167 V76 V167 -2.1993314761124857e-21

R76_168 V76 V168 -180.74720528111817
L76_168 V76 V168 2.04988192531515e-12
C76_168 V76 V168 1.150135894674819e-19

R76_169 V76 V169 -596.0701265554575
L76_169 V76 V169 1.5058043495550416e-09
C76_169 V76 V169 1.5989650819508244e-19

R76_170 V76 V170 -17222.54931370728
L76_170 V76 V170 -5.041047079165853e-12
C76_170 V76 V170 -5.32937012075424e-20

R76_171 V76 V171 -398.6264812122926
L76_171 V76 V171 -4.105750218139117e-12
C76_171 V76 V171 6.70451101041717e-20

R76_172 V76 V172 -2055.9053054921765
L76_172 V76 V172 8.841999869884015e-13
C76_172 V76 V172 1.3980929713434874e-20

R76_173 V76 V173 -1378.4055486463133
L76_173 V76 V173 -1.5127479573449727e-12
C76_173 V76 V173 -2.662281609030057e-19

R76_174 V76 V174 8452.089220856875
L76_174 V76 V174 2.4484633699954223e-11
C76_174 V76 V174 -6.862409165979361e-20

R76_175 V76 V175 1217.9456972004918
L76_175 V76 V175 3.013491657946727e-12
C76_175 V76 V175 -6.932877181296349e-20

R76_176 V76 V176 407.3585450868929
L76_176 V76 V176 -3.6725829595431473e-13
C76_176 V76 V176 -6.43581816436327e-19

R76_177 V76 V177 459.8264544209256
L76_177 V76 V177 1.3965996727123492e-12
C76_177 V76 V177 1.7308863745746031e-19

R76_178 V76 V178 1550.3578837417854
L76_178 V76 V178 8.82742317440356e-12
C76_178 V76 V178 6.801921221697534e-21

R76_179 V76 V179 2473.7820325597136
L76_179 V76 V179 4.4076080165913105e-12
C76_179 V76 V179 4.538459348036764e-20

R76_180 V76 V180 3631.083418107716
L76_180 V76 V180 9.067705223883092e-13
C76_180 V76 V180 5.288079771999316e-19

R76_181 V76 V181 -1107.3637871130522
L76_181 V76 V181 1.7892418480535713e-11
C76_181 V76 V181 1.456245615237801e-19

R76_182 V76 V182 -445.2843163543317
L76_182 V76 V182 -7.3793922518544e-12
C76_182 V76 V182 3.6671430397591086e-20

R76_183 V76 V183 1447.4870380876775
L76_183 V76 V183 2.1245202282075116e-12
C76_183 V76 V183 1.1068254019335725e-19

R76_184 V76 V184 2768.496507764544
L76_184 V76 V184 8.122511186457531e-13
C76_184 V76 V184 -1.4355765326013707e-19

R76_185 V76 V185 -691.6192388552179
L76_185 V76 V185 -1.9309995673936885e-12
C76_185 V76 V185 -1.9445581681958103e-19

R76_186 V76 V186 983.2929991085408
L76_186 V76 V186 1.1583666683806802e-12
C76_186 V76 V186 5.493021011113935e-20

R76_187 V76 V187 12990.968937556525
L76_187 V76 V187 2.3962185447060937e-11
C76_187 V76 V187 -1.4720949363791823e-19

R76_188 V76 V188 -254.93643543479214
L76_188 V76 V188 -4.199485117555651e-13
C76_188 V76 V188 -1.175628351852861e-19

R76_189 V76 V189 773.3051748426077
L76_189 V76 V189 1.8172347752134207e-11
C76_189 V76 V189 4.4596385964787006e-20

R76_190 V76 V190 888.0270523094224
L76_190 V76 V190 -9.00460257519158e-12
C76_190 V76 V190 4.678300049466548e-20

R76_191 V76 V191 -559.3400687745742
L76_191 V76 V191 -8.223367995421747e-13
C76_191 V76 V191 -4.915672264882517e-20

R76_192 V76 V192 803.5584118990741
L76_192 V76 V192 1.6166904335616898e-12
C76_192 V76 V192 3.1485518966507736e-19

R76_193 V76 V193 3620.820634886262
L76_193 V76 V193 2.05376597184571e-12
C76_193 V76 V193 1.5319193945950157e-20

R76_194 V76 V194 -1084.1319691830993
L76_194 V76 V194 -4.2716293331661086e-11
C76_194 V76 V194 2.141586919758801e-19

R76_195 V76 V195 661.2923893563878
L76_195 V76 V195 7.296752313466429e-13
C76_195 V76 V195 4.3000582513082325e-19

R76_196 V76 V196 614.8220496274797
L76_196 V76 V196 -1.1418171659133524e-12
C76_196 V76 V196 -7.802889475567039e-19

R76_197 V76 V197 -1335.2001853693823
L76_197 V76 V197 -5.0993811826976046e-11
C76_197 V76 V197 -1.0218269488407034e-20

R76_198 V76 V198 5591.682364117237
L76_198 V76 V198 5.6106307340972075e-12
C76_198 V76 V198 1.322481486474846e-19

R76_199 V76 V199 422.2829709010407
L76_199 V76 V199 6.159620580947174e-12
C76_199 V76 V199 -3.671442360245347e-20

R76_200 V76 V200 -434.4424630695969
L76_200 V76 V200 1.229087320971613e-12
C76_200 V76 V200 1.1537937081558619e-19

R77_77 V77 0 -2682.4494410997754
L77_77 V77 0 -6.747528106597111e-13
C77_77 V77 0 4.494128606956321e-19

R77_78 V77 V78 860.5592761793466
L77_78 V77 V78 -3.418818018028496e-12
C77_78 V77 V78 -7.349335788944158e-20

R77_79 V77 V79 1211.784862748676
L77_79 V77 V79 -2.3321259671351964e-12
C77_79 V77 V79 -1.2949668852812074e-19

R77_80 V77 V80 818.5688500830797
L77_80 V77 V80 -1.6859913397319935e-12
C77_80 V77 V80 -2.226828287327215e-19

R77_81 V77 V81 303.23882174787985
L77_81 V77 V81 1.0561012855089862e-12
C77_81 V77 V81 3.5619016395511807e-19

R77_82 V77 V82 -1767.399856151099
L77_82 V77 V82 -1.918612853874357e-12
C77_82 V77 V82 -3.5644533644828194e-19

R77_83 V77 V83 -1447.010667162947
L77_83 V77 V83 -3.371494554182219e-12
C77_83 V77 V83 -1.9389570183753161e-19

R77_84 V77 V84 -2203.011146828953
L77_84 V77 V84 -2.308997223554702e-12
C77_84 V77 V84 -2.403567724874351e-19

R77_85 V77 V85 -1470.2212743823982
L77_85 V77 V85 2.719728590009733e-12
C77_85 V77 V85 3.5615920807349435e-19

R77_86 V77 V86 -510.0305528384533
L77_86 V77 V86 5.025141513928682e-12
C77_86 V77 V86 8.917329523183994e-20

R77_87 V77 V87 -1251.909678008587
L77_87 V77 V87 2.913485798549065e-12
C77_87 V77 V87 2.4212262611215913e-19

R77_88 V77 V88 -846.8967663536775
L77_88 V77 V88 1.781933629377633e-12
C77_88 V77 V88 3.6768492993092806e-19

R77_89 V77 V89 -584.0876537571822
L77_89 V77 V89 7.990938608284778e-13
C77_89 V77 V89 3.3982020768901206e-19

R77_90 V77 V90 531.3250468473175
L77_90 V77 V90 9.66640196700112e-13
C77_90 V77 V90 5.77656148001297e-19

R77_91 V77 V91 489.0409990902976
L77_91 V77 V91 2.7430804178380173e-12
C77_91 V77 V91 4.519709307509775e-20

R77_92 V77 V92 529.4493300597401
L77_92 V77 V92 4.993809134519928e-12
C77_92 V77 V92 6.634121945503975e-21

R77_93 V77 V93 374.7915805203733
L77_93 V77 V93 -1.1468323623095548e-12
C77_93 V77 V93 -5.191206294304956e-19

R77_94 V77 V94 1989.4835985610705
L77_94 V77 V94 -1.6081999332812685e-12
C77_94 V77 V94 -4.1281317708765634e-19

R77_95 V77 V95 -6915049.346697509
L77_95 V77 V95 -1.896662322136373e-12
C77_95 V77 V95 -3.079013224348557e-19

R77_96 V77 V96 3525.5700170904793
L77_96 V77 V96 -1.4605782231968432e-12
C77_96 V77 V96 -3.9095917781716796e-19

R77_97 V77 V97 -1054.2560832675936
L77_97 V77 V97 -1.0639355909259956e-12
C77_97 V77 V97 -5.724540250573362e-19

R77_98 V77 V98 -579.84639835416
L77_98 V77 V98 -4.0707364128486114e-12
C77_98 V77 V98 -2.1073390258663812e-19

R77_99 V77 V99 -499.49280280388183
L77_99 V77 V99 6.622495553422289e-12
C77_99 V77 V99 1.9342413940867986e-19

R77_100 V77 V100 -524.5323630960717
L77_100 V77 V100 1.453048187524629e-10
C77_100 V77 V100 1.8546709290106927e-19

R77_101 V77 V101 -927.0308471668995
L77_101 V77 V101 1.3332662227527238e-12
C77_101 V77 V101 6.546731116197242e-19

R77_102 V77 V102 -13387.593404594809
L77_102 V77 V102 3.2090906979433794e-12
C77_102 V77 V102 2.637692017324765e-19

R77_103 V77 V103 5986.466475866227
L77_103 V77 V103 1.0261297694293345e-11
C77_103 V77 V103 4.044424799433903e-20

R77_104 V77 V104 -8189.052130732819
L77_104 V77 V104 1.0121958319592502e-11
C77_104 V77 V104 3.964201970509543e-20

R77_105 V77 V105 355.24259213666255
L77_105 V77 V105 1.7146989559706221e-12
C77_105 V77 V105 2.2790664314649173e-19

R77_106 V77 V106 2237.3629380098364
L77_106 V77 V106 4.434275443378458e-12
C77_106 V77 V106 1.470549443317273e-19

R77_107 V77 V107 910.0984603330267
L77_107 V77 V107 -8.463163640346821e-12
C77_107 V77 V107 -6.500302184109933e-20

R77_108 V77 V108 766.3364165759214
L77_108 V77 V108 2.7487850330091335e-12
C77_108 V77 V108 1.518173202074627e-19

R77_109 V77 V109 -936.4248072710246
L77_109 V77 V109 1.185151453986189e-11
C77_109 V77 V109 -2.6523707871031266e-19

R77_110 V77 V110 4426.21899356089
L77_110 V77 V110 -4.554335273593787e-12
C77_110 V77 V110 -1.6702013619470944e-19

R77_111 V77 V111 14664.629884523012
L77_111 V77 V111 4.138156427842944e-12
C77_111 V77 V111 4.9742406653567446e-20

R77_112 V77 V112 -7021.357408083123
L77_112 V77 V112 -1.5260261784943016e-11
C77_112 V77 V112 -1.3784511067243064e-19

R77_113 V77 V113 -1929.1877951853307
L77_113 V77 V113 -1.586614562486092e-12
C77_113 V77 V113 -3.458481985068603e-19

R77_114 V77 V114 -3588.8141048202287
L77_114 V77 V114 -4.3044748262092715e-12
C77_114 V77 V114 -2.0435538158113286e-19

R77_115 V77 V115 -824.3199359373752
L77_115 V77 V115 -2.0114330686936315e-11
C77_115 V77 V115 -4.3398183617195975e-20

R77_116 V77 V116 -668.2589135552531
L77_116 V77 V116 -2.5318037555016226e-12
C77_116 V77 V116 -2.078720142413033e-19

R77_117 V77 V117 444.23577582079054
L77_117 V77 V117 -3.4222169163378734e-12
C77_117 V77 V117 4.419718399278033e-21

R77_118 V77 V118 -1566.8340985790883
L77_118 V77 V118 2.1775183921041015e-12
C77_118 V77 V118 3.214732651000786e-19

R77_119 V77 V119 2057.5426721012423
L77_119 V77 V119 4.115700036472493e-11
C77_119 V77 V119 1.4340041034389835e-19

R77_120 V77 V120 967.7850660814978
L77_120 V77 V120 3.199497711073549e-12
C77_120 V77 V120 3.2303174091155305e-19

R77_121 V77 V121 -818.7508698966612
L77_121 V77 V121 1.4957524175525082e-12
C77_121 V77 V121 3.917534288019441e-19

R77_122 V77 V122 3641.969710213935
L77_122 V77 V122 -4.715455526151003e-12
C77_122 V77 V122 -1.0320995104388504e-19

R77_123 V77 V123 2837.811818142783
L77_123 V77 V123 -8.624859659798172e-12
C77_123 V77 V123 -1.3414421392090985e-19

R77_124 V77 V124 9570.032297020884
L77_124 V77 V124 -6.9609149519319055e-12
C77_124 V77 V124 -1.741726504176142e-19

R77_125 V77 V125 -3208.4711801847893
L77_125 V77 V125 1.7331291597375552e-12
C77_125 V77 V125 1.2470165637136183e-19

R77_126 V77 V126 835.775128136964
L77_126 V77 V126 -2.6792772445240388e-11
C77_126 V77 V126 -3.257980274168597e-20

R77_127 V77 V127 7234.915783821377
L77_127 V77 V127 1.1744678331495303e-11
C77_127 V77 V127 -1.3273831331486538e-20

R77_128 V77 V128 -9084.941114643234
L77_128 V77 V128 3.034982302655773e-12
C77_128 V77 V128 1.569511479014348e-20

R77_129 V77 V129 559.9340015924047
L77_129 V77 V129 -1.7252826132128483e-12
C77_129 V77 V129 -3.6039658902110826e-19

R77_130 V77 V130 -1075.7986101077745
L77_130 V77 V130 8.815045118574148e-12
C77_130 V77 V130 8.784922336492696e-20

R77_131 V77 V131 -1945.8438514908175
L77_131 V77 V131 2.0269029266804654e-11
C77_131 V77 V131 5.125027193448901e-20

R77_132 V77 V132 -2109.5147715482162
L77_132 V77 V132 -5.323981104322447e-12
C77_132 V77 V132 2.4010117632136014e-20

R77_133 V77 V133 -2534.1369211735328
L77_133 V77 V133 -5.739199338420539e-11
C77_133 V77 V133 3.30005189242953e-20

R77_134 V77 V134 -1781.7215895396362
L77_134 V77 V134 -2.8470744610936238e-12
C77_134 V77 V134 -1.6349144296049567e-19

R77_135 V77 V135 -1654.1445066859499
L77_135 V77 V135 -9.988972419076149e-12
C77_135 V77 V135 -2.7163314239636654e-20

R77_136 V77 V136 -1167.1242906761292
L77_136 V77 V136 -3.3133952548279088e-12
C77_136 V77 V136 -1.802841481022349e-19

R77_137 V77 V137 -1024.4354638970428
L77_137 V77 V137 -2.6569872922323096e-12
C77_137 V77 V137 -3.7905867674962885e-20

R77_138 V77 V138 1078.5480506335666
L77_138 V77 V138 1.1576927949692283e-11
C77_138 V77 V138 6.798501173946642e-20

R77_139 V77 V139 1035.4684233298944
L77_139 V77 V139 3.859153776154484e-12
C77_139 V77 V139 1.5193195079875498e-19

R77_140 V77 V140 658.4135756191416
L77_140 V77 V140 7.156451869349811e-12
C77_140 V77 V140 1.4346002584134672e-19

R77_141 V77 V141 -2020.5303964973493
L77_141 V77 V141 4.518195770188098e-12
C77_141 V77 V141 2.1663901994526978e-20

R77_142 V77 V142 4205.469013236211
L77_142 V77 V142 2.2343759863353864e-12
C77_142 V77 V142 1.0067141065348069e-19

R77_143 V77 V143 2344.154108623271
L77_143 V77 V143 -2.3405340119268578e-12
C77_143 V77 V143 -2.1208479387812206e-19

R77_144 V77 V144 5165.258213176927
L77_144 V77 V144 3.305781280694174e-11
C77_144 V77 V144 3.7410850058937266e-20

R77_145 V77 V145 370.021674897226
L77_145 V77 V145 1.60833279417883e-12
C77_145 V77 V145 4.2497562823029225e-20

R77_146 V77 V146 6375.2162018658255
L77_146 V77 V146 -2.273612401677572e-12
C77_146 V77 V146 -8.997653714474741e-20

R77_147 V77 V147 -950.7623447645402
L77_147 V77 V147 5.7155531580064944e-12
C77_147 V77 V147 4.704174222096804e-21

R77_148 V77 V148 -3663.493539381292
L77_148 V77 V148 5.899806659940525e-12
C77_148 V77 V148 -4.891760625493666e-21

R77_149 V77 V149 -859.4097927086991
L77_149 V77 V149 3.2871676422126288e-12
C77_149 V77 V149 4.678474589535315e-19

R77_150 V77 V150 -512.8355688093587
L77_150 V77 V150 5.959412384332872e-12
C77_150 V77 V150 -1.7908467545402752e-19

R77_151 V77 V151 3094.946820085592
L77_151 V77 V151 1.6400283375779516e-12
C77_151 V77 V151 2.259190399549656e-19

R77_152 V77 V152 -1301.0093632779697
L77_152 V77 V152 1.37918741603807e-11
C77_152 V77 V152 -5.207226685703351e-20

R77_153 V77 V153 -908.9290566948762
L77_153 V77 V153 -2.4662473040160862e-12
C77_153 V77 V153 -2.6950719418583484e-19

R77_154 V77 V154 -2879.8846424592125
L77_154 V77 V154 -5.973797342326736e-12
C77_154 V77 V154 1.5040804513271596e-19

R77_155 V77 V155 -689.6100748777534
L77_155 V77 V155 2.3117159499193232e-11
C77_155 V77 V155 1.0606011984262986e-19

R77_156 V77 V156 3361.080703672886
L77_156 V77 V156 -5.7741768320279685e-12
C77_156 V77 V156 5.879450245116718e-20

R77_157 V77 V157 -8728.179214045887
L77_157 V77 V157 -1.1359526074570467e-12
C77_157 V77 V157 -6.641235625988893e-19

R77_158 V77 V158 776.1841635544064
L77_158 V77 V158 6.183156555579667e-12
C77_158 V77 V158 9.1309912071891e-21

R77_159 V77 V159 1194.4118371497414
L77_159 V77 V159 -1.7304526331076738e-12
C77_159 V77 V159 -2.0192816115177868e-19

R77_160 V77 V160 2950.1756079627885
L77_160 V77 V160 -2.740628433714821e-12
C77_160 V77 V160 -5.62656898207104e-20

R77_161 V77 V161 513.7943987879513
L77_161 V77 V161 3.661347429178332e-12
C77_161 V77 V161 2.946964659897672e-19

R77_162 V77 V162 1509.2793809231855
L77_162 V77 V162 8.14658100522956e-12
C77_162 V77 V162 -9.260388593952779e-20

R77_163 V77 V163 2158.3805687604095
L77_163 V77 V163 -2.1796783453764866e-12
C77_163 V77 V163 -2.2288224921717104e-19

R77_164 V77 V164 911.2126087941703
L77_164 V77 V164 2.179347909917674e-11
C77_164 V77 V164 4.353905597901656e-21

R77_165 V77 V165 772.2380497716089
L77_165 V77 V165 6.89338873625246e-13
C77_165 V77 V165 5.234440478541251e-19

R77_166 V77 V166 -416.45890409904996
L77_166 V77 V166 2.1600917560879036e-12
C77_166 V77 V166 9.023037886702349e-20

R77_167 V77 V167 -7388.047219342762
L77_167 V77 V167 2.0512504327707734e-12
C77_167 V77 V167 2.067793516763698e-19

R77_168 V77 V168 -896.8949428433756
L77_168 V77 V168 2.3517731031896985e-12
C77_168 V77 V168 1.9827636394635982e-19

R77_169 V77 V169 -557.1570756336295
L77_169 V77 V169 -1.1032657629567628e-12
C77_169 V77 V169 -4.418388065106478e-19

R77_170 V77 V170 929.4175237697087
L77_170 V77 V170 -1.2044664346442481e-11
C77_170 V77 V170 2.249356069619128e-19

R77_171 V77 V171 -1994.7021998428593
L77_171 V77 V171 1.4642596328670762e-12
C77_171 V77 V171 3.1147065805225175e-19

R77_172 V77 V172 11997.881853065037
L77_172 V77 V172 9.687177301352996e-12
C77_172 V77 V172 6.603813500974873e-20

R77_173 V77 V173 1067.1458966664309
L77_173 V77 V173 -1.647380809934218e-12
C77_173 V77 V173 -2.3356365310427985e-19

R77_174 V77 V174 1525.8559727507627
L77_174 V77 V174 -9.944485973874002e-13
C77_174 V77 V174 -4.378646015946638e-19

R77_175 V77 V175 38843.34967013448
L77_175 V77 V175 -1.638923398794462e-12
C77_175 V77 V175 -1.9387367156148803e-19

R77_176 V77 V176 -28024.366665977283
L77_176 V77 V176 -1.2358530591550627e-12
C77_176 V77 V176 -2.3580553320149317e-19

R77_177 V77 V177 902.2892377698417
L77_177 V77 V177 3.035342773701126e-12
C77_177 V77 V177 2.4575978942205477e-19

R77_178 V77 V178 -6927.238269654843
L77_178 V77 V178 3.3838248109921644e-12
C77_178 V77 V178 -9.380250961114058e-20

R77_179 V77 V179 -9832.095731092517
L77_179 V77 V179 -2.9763749558226138e-12
C77_179 V77 V179 -2.848912387726165e-19

R77_180 V77 V180 1935.98203977921
L77_180 V77 V180 -3.6342681488615566e-11
C77_180 V77 V180 -1.4951293908961717e-19

R77_181 V77 V181 -1083.8941882054648
L77_181 V77 V181 5.348411220058608e-12
C77_181 V77 V181 3.572282501717477e-19

R77_182 V77 V182 -767.9987687972956
L77_182 V77 V182 1.2987990897975654e-12
C77_182 V77 V182 2.5389996070401986e-19

R77_183 V77 V183 1608.1129526085515
L77_183 V77 V183 -4.6960850321699975e-12
C77_183 V77 V183 -1.665555286318655e-20

R77_184 V77 V184 3206.1609779192254
L77_184 V77 V184 7.568344092105965e-12
C77_184 V77 V184 9.869622233358193e-20

R77_185 V77 V185 -40836.86163331154
L77_185 V77 V185 1.574124233057044e-12
C77_185 V77 V185 -3.7345957424195217e-19

R77_186 V77 V186 -5649.329911800853
L77_186 V77 V186 4.879247641731667e-12
C77_186 V77 V186 1.949968533294312e-19

R77_187 V77 V187 -7637.298034973273
L77_187 V77 V187 1.7542609194721367e-12
C77_187 V77 V187 2.6394167954669734e-19

R77_188 V77 V188 -836.8523451557892
L77_188 V77 V188 1.4128827993831276e-12
C77_188 V77 V188 2.9411274220388804e-19

R77_189 V77 V189 -2120.65430661353
L77_189 V77 V189 -1.0902213128438754e-12
C77_189 V77 V189 -8.094575533475091e-21

R77_190 V77 V190 1283.9980836048921
L77_190 V77 V190 -3.2673671175663375e-12
C77_190 V77 V190 -2.1385260350522845e-19

R77_191 V77 V191 -3706.186494607141
L77_191 V77 V191 1.561109072566854e-12
C77_191 V77 V191 1.0724664875828394e-19

R77_192 V77 V192 1684.0002557429739
L77_192 V77 V192 -9.47057026553401e-12
C77_192 V77 V192 -1.8762179591633586e-19

R77_193 V77 V193 4432.584883515772
L77_193 V77 V193 -1.3653205356956345e-12
C77_193 V77 V193 -1.430093279269786e-19

R77_194 V77 V194 -2869.874425759632
L77_194 V77 V194 -1.4566059707453633e-12
C77_194 V77 V194 -3.256486331427017e-19

R77_195 V77 V195 2183.632424165286
L77_195 V77 V195 -1.2537137680665237e-12
C77_195 V77 V195 -2.711442655347887e-19

R77_196 V77 V196 1653.355563174299
L77_196 V77 V196 -1.0996748621733241e-12
C77_196 V77 V196 -1.9672661542539989e-19

R77_197 V77 V197 1641.3464766961029
L77_197 V77 V197 2.350739343467882e-12
C77_197 V77 V197 1.9397414196546992e-19

R77_198 V77 V198 -918.4320026167107
L77_198 V77 V198 4.070870432311183e-12
C77_198 V77 V198 8.100855965537381e-20

R77_199 V77 V199 -1347.6960137228484
L77_199 V77 V199 -1.6894907171759281e-12
C77_199 V77 V199 -2.0973918173510568e-19

R77_200 V77 V200 -1621.2449575656171
L77_200 V77 V200 -4.5451312501513495e-11
C77_200 V77 V200 1.3874180772765856e-19

R78_78 V78 0 -150.09674395876115
L78_78 V78 0 9.203682112380786e-13
C78_78 V78 0 5.499687397978716e-19

R78_79 V78 V79 -676.6923687037823
L78_79 V78 V79 2.770602219332384e-11
C78_79 V78 V79 9.17124082205108e-20

R78_80 V78 V80 -452.0064641484376
L78_80 V78 V80 1.510586767469482e-11
C78_80 V78 V80 1.3785085367432882e-19

R78_81 V78 V81 -284.44714094500364
L78_81 V78 V81 1.670713515614054e-11
C78_81 V78 V81 3.99519306500163e-20

R78_82 V78 V82 320.4447274594448
L78_82 V78 V82 1.6498787704189792e-11
C78_82 V78 V82 5.122084608742287e-20

R78_83 V78 V83 797.7929588945241
L78_83 V78 V83 -1.3036895765362208e-11
C78_83 V78 V83 -8.630968333585052e-20

R78_84 V78 V84 1150.8671986389936
L78_84 V78 V84 -5.132184875803064e-12
C78_84 V78 V84 -1.578471377627281e-19

R78_85 V78 V85 1083.175055335217
L78_85 V78 V85 -1.707601542081525e-11
C78_85 V78 V85 -1.3613048203527473e-20

R78_86 V78 V86 159.2350070510169
L78_86 V78 V86 1.0299495310641554e-12
C78_86 V78 V86 5.770627602967063e-19

R78_87 V78 V87 1348.7011990648869
L78_87 V78 V87 -7.746233804958629e-12
C78_87 V78 V87 -1.517841206952551e-19

R78_88 V78 V88 798.0234990175652
L78_88 V78 V88 -1.7431523765464733e-11
C78_88 V78 V88 -1.3333815194969626e-19

R78_89 V78 V89 532.0709637870951
L78_89 V78 V89 4.600979934363952e-12
C78_89 V78 V89 2.800546582956889e-22

R78_90 V78 V90 -131.48465918052747
L78_90 V78 V90 -2.216564867145535e-12
C78_90 V78 V90 -3.7846089541333673e-19

R78_91 V78 V91 -445.1844654321293
L78_91 V78 V91 3.4867919200092916e-12
C78_91 V78 V91 2.981237803407111e-19

R78_92 V78 V92 -807.8536632361164
L78_92 V78 V92 2.4464048205618785e-12
C78_92 V78 V92 3.0902151981983828e-19

R78_93 V78 V93 -388.85771805974827
L78_93 V78 V93 -5.588101594015557e-12
C78_93 V78 V93 -6.002413622618733e-20

R78_94 V78 V94 -14099.166474645634
L78_94 V78 V94 -2.052998133513392e-12
C78_94 V78 V94 -1.6863145889072012e-19

R78_95 V78 V95 3555.5442403393577
L78_95 V78 V95 -8.01713316063215e-12
C78_95 V78 V95 -7.498383048518373e-21

R78_96 V78 V96 -5300.741574063593
L78_96 V78 V96 -3.411431003470084e-12
C78_96 V78 V96 -5.821937157344517e-20

R78_97 V78 V97 2219.4615934452927
L78_97 V78 V97 -6.6538108702398175e-12
C78_97 V78 V97 1.1901323462106915e-19

R78_98 V78 V98 212.4291672862868
L78_98 V78 V98 1.5091692432482749e-12
C78_98 V78 V98 2.982066667117584e-19

R78_99 V78 V99 1023.0212915195493
L78_99 V78 V99 -4.459666413959683e-12
C78_99 V78 V99 -2.5402999397506766e-19

R78_100 V78 V100 -14851.060435302756
L78_100 V78 V100 -4.860570115012013e-12
C78_100 V78 V100 -2.8696144956956034e-19

R78_101 V78 V101 -2032.8249241617425
L78_101 V78 V101 9.756467948340842e-12
C78_101 V78 V101 -3.0634939720077507e-20

R78_102 V78 V102 -374.86402154913594
L78_102 V78 V102 -2.265170737463348e-11
C78_102 V78 V102 1.631275220564203e-20

R78_103 V78 V103 687.5198551750158
L78_103 V78 V103 2.1339486301903126e-12
C78_103 V78 V103 2.6715745091659724e-19

R78_104 V78 V104 449.451132969021
L78_104 V78 V104 2.042709403039613e-12
C78_104 V78 V104 2.507069395607177e-19

R78_105 V78 V105 1553.1312660721812
L78_105 V78 V105 5.1289850947669605e-12
C78_105 V78 V105 2.360510308369619e-20

R78_106 V78 V106 345.6086405899988
L78_106 V78 V106 -3.225770361200805e-12
C78_106 V78 V106 -3.11348073724166e-19

R78_107 V78 V107 -497.22648675042467
L78_107 V78 V107 -3.482135716217769e-12
C78_107 V78 V107 -4.267324662062719e-20

R78_108 V78 V108 -919.1673818316712
L78_108 V78 V108 -4.70351499910934e-12
C78_108 V78 V108 -2.906226410823945e-20

R78_109 V78 V109 11062.549242833637
L78_109 V78 V109 -6.588100198444003e-12
C78_109 V78 V109 5.1353652209790125e-20

R78_110 V78 V110 -277.3297739271671
L78_110 V78 V110 3.3956638116771397e-12
C78_110 V78 V110 1.4389455340574122e-19

R78_111 V78 V111 -807.2334682538487
L78_111 V78 V111 -1.1593784619040332e-11
C78_111 V78 V111 -7.519097589254127e-20

R78_112 V78 V112 -582.2005106465213
L78_112 V78 V112 2.712156543454986e-11
C78_112 V78 V112 5.2033301780853085e-20

R78_113 V78 V113 -246.8223833456464
L78_113 V78 V113 -2.7089693632218536e-12
C78_113 V78 V113 -1.530820278634288e-19

R78_114 V78 V114 -371.5725233675162
L78_114 V78 V114 5.739933608324144e-12
C78_114 V78 V114 2.3921612366315586e-19

R78_115 V78 V115 358.1759647564519
L78_115 V78 V115 5.372266453131558e-12
C78_115 V78 V115 5.506804154546335e-20

R78_116 V78 V116 464.34963621008916
L78_116 V78 V116 -4.81787124820277e-11
C78_116 V78 V116 -4.0816937552618423e-20

R78_117 V78 V117 861.8167008483468
L78_117 V78 V117 4.680605513867875e-12
C78_117 V78 V117 6.531350702614857e-20

R78_118 V78 V118 83.70229690427911
L78_118 V78 V118 1.0333627906602172e-10
C78_118 V78 V118 -2.7060447682371217e-19

R78_119 V78 V119 1009.650439431876
L78_119 V78 V119 -7.112685309229386e-12
C78_119 V78 V119 -1.0550441422740254e-19

R78_120 V78 V120 2486.710139016758
L78_120 V78 V120 -8.109039951592895e-12
C78_120 V78 V120 -1.5819176006163637e-19

R78_121 V78 V121 370.00170998374
L78_121 V78 V121 4.305253952006604e-12
C78_121 V78 V121 1.7956469323628873e-19

R78_122 V78 V122 -195.05705317171444
L78_122 V78 V122 -3.1313852506013483e-12
C78_122 V78 V122 -1.3462543881441295e-19

R78_123 V78 V123 -577.3732552541827
L78_123 V78 V123 3.301185808327761e-12
C78_123 V78 V123 2.3450068392798595e-19

R78_124 V78 V124 -642.6648397193295
L78_124 V78 V124 2.2484829788689215e-12
C78_124 V78 V124 3.8015876261618897e-19

R78_125 V78 V125 -948.1094163253106
L78_125 V78 V125 -9.779488479155731e-12
C78_125 V78 V125 -1.5912417058222632e-19

R78_126 V78 V126 -85.87124412760488
L78_126 V78 V126 5.814540294406459e-12
C78_126 V78 V126 2.684098839078811e-19

R78_127 V78 V127 -328.60773529230624
L78_127 V78 V127 -9.163432966235504e-12
C78_127 V78 V127 -1.272659110658368e-19

R78_128 V78 V128 -435.901469937899
L78_128 V78 V128 -1.0507866214679729e-11
C78_128 V78 V128 -1.3335679191001864e-19

R78_129 V78 V129 -251.28354319953095
L78_129 V78 V129 -1.9151414382167616e-12
C78_129 V78 V129 -1.910545239135922e-19

R78_130 V78 V130 97.33385884952351
L78_130 V78 V130 2.355113732271627e-12
C78_130 V78 V130 3.257650600088727e-20

R78_131 V78 V131 191.82190153808324
L78_131 V78 V131 -8.124969781681741e-12
C78_131 V78 V131 -1.015805207189803e-19

R78_132 V78 V132 152.93933604743697
L78_132 V78 V132 -4.6752195084389476e-12
C78_132 V78 V132 -1.8697805460688742e-19

R78_133 V78 V133 417.80026231724696
L78_133 V78 V133 1.632802347098841e-12
C78_133 V78 V133 3.2753983051858375e-19

R78_134 V78 V134 385.7661541258432
L78_134 V78 V134 -1.3389050102299344e-12
C78_134 V78 V134 -4.966511439028031e-19

R78_135 V78 V135 1157.6989428788202
L78_135 V78 V135 2.397277539742652e-12
C78_135 V78 V135 3.5369286577737815e-19

R78_136 V78 V136 427.04278547209
L78_136 V78 V136 3.003564297611844e-12
C78_136 V78 V136 3.855682173119693e-19

R78_137 V78 V137 917.3908741746219
L78_137 V78 V137 4.365156589042371e-12
C78_137 V78 V137 1.117865621233512e-19

R78_138 V78 V138 -135.71224789816392
L78_138 V78 V138 1.8423384357997928e-12
C78_138 V78 V138 4.612678780931459e-19

R78_139 V78 V139 -185.98389642031327
L78_139 V78 V139 -2.6879892068205247e-12
C78_139 V78 V139 -3.4644817513877068e-19

R78_140 V78 V140 -102.01001930132668
L78_140 V78 V140 -2.9076956925557305e-12
C78_140 V78 V140 -3.97569520484054e-19

R78_141 V78 V141 493.73715615565135
L78_141 V78 V141 -1.7187470147832932e-12
C78_141 V78 V141 -3.4090174815255037e-19

R78_142 V78 V142 -6026.254194627157
L78_142 V78 V142 1.3028980723877908e-12
C78_142 V78 V142 8.989245816557435e-20

R78_143 V78 V143 311.78245658694857
L78_143 V78 V143 -8.053255069443786e-11
C78_143 V78 V143 -4.8672485855795995e-20

R78_144 V78 V144 201.4879561027411
L78_144 V78 V144 2.6223336900326253e-11
C78_144 V78 V144 -1.6200589269806807e-20

R78_145 V78 V145 -494.3130020374383
L78_145 V78 V145 3.651013806084658e-11
C78_145 V78 V145 -3.481386660778799e-20

R78_146 V78 V146 195.49945149267364
L78_146 V78 V146 -8.786313282219306e-13
C78_146 V78 V146 -2.289783935869861e-19

R78_147 V78 V147 1092.9197232195052
L78_147 V78 V147 3.442297239946533e-12
C78_147 V78 V147 3.2326239056142384e-19

R78_148 V78 V148 -2021.5442418660612
L78_148 V78 V148 2.847307857290668e-12
C78_148 V78 V148 2.9635619355507774e-19

R78_149 V78 V149 -426.9370873375632
L78_149 V78 V149 1.6513511301184172e-12
C78_149 V78 V149 3.764285807409681e-19

R78_150 V78 V150 169.39711984262348
L78_150 V78 V150 -2.530874331727114e-11
C78_150 V78 V150 -2.3863329356948173e-19

R78_151 V78 V151 -288.47603942000984
L78_151 V78 V151 -5.142015951335941e-11
C78_151 V78 V151 -3.462410068136467e-20

R78_152 V78 V152 -252.4652530748912
L78_152 V78 V152 -6.095098655979305e-12
C78_152 V78 V152 -1.0596514439362139e-19

R78_153 V78 V153 1574.8628315104609
L78_153 V78 V153 -1.0062315656291269e-11
C78_153 V78 V153 1.8703896643201144e-20

R78_154 V78 V154 -182.5714333959523
L78_154 V78 V154 3.1869237181773497e-12
C78_154 V78 V154 3.6112069820682042e-19

R78_155 V78 V155 446.9948150792641
L78_155 V78 V155 -4.423318464007653e-12
C78_155 V78 V155 -1.2795428201827376e-19

R78_156 V78 V156 433.23823845433844
L78_156 V78 V156 -6.620909100379424e-12
C78_156 V78 V156 -1.2662914670350212e-19

R78_157 V78 V157 227.45532475503626
L78_157 V78 V157 -2.0573492783730074e-12
C78_157 V78 V157 -2.7605326165156187e-19

R78_158 V78 V158 -7484.380277708869
L78_158 V78 V158 4.5600922398959604e-12
C78_158 V78 V158 -1.6507268656984636e-19

R78_159 V78 V159 316.6020299830232
L78_159 V78 V159 4.433580707437431e-12
C78_159 V78 V159 1.8376365540085052e-19

R78_160 V78 V160 165.70600708017952
L78_160 V78 V160 4.5129829150279085e-12
C78_160 V78 V160 1.9284741761511498e-19

R78_161 V78 V161 -157.3256616457634
L78_161 V78 V161 -3.448926959644615e-12
C78_161 V78 V161 -1.6562578002628478e-19

R78_162 V78 V162 -327.8573063493555
L78_162 V78 V162 -4.777477296782923e-12
C78_162 V78 V162 1.9410143041655224e-20

R78_163 V78 V163 -169.03422454456162
L78_163 V78 V163 -3.341175090258726e-12
C78_163 V78 V163 -2.018367527030949e-19

R78_164 V78 V164 -100.64403751828512
L78_164 V78 V164 -1.4604505339190424e-11
C78_164 V78 V164 -1.4531654210362488e-19

R78_165 V78 V165 -555.2882233023494
L78_165 V78 V165 1.935138514114668e-12
C78_165 V78 V165 3.3803498461602425e-19

R78_166 V78 V166 374.83933548423556
L78_166 V78 V166 2.3339617106366162e-11
C78_166 V78 V166 8.617540423664397e-20

R78_167 V78 V167 -742.2023270012589
L78_167 V78 V167 -4.132589687546086e-12
C78_167 V78 V167 -6.868729100204871e-20

R78_168 V78 V168 3104.747717055552
L78_168 V78 V168 -1.943640160244789e-12
C78_168 V78 V168 -1.4008804149982232e-19

R78_169 V78 V169 123.84990870901625
L78_169 V78 V169 6.105799874730429e-12
C78_169 V78 V169 1.0638932580534084e-19

R78_170 V78 V170 163.3266848949189
L78_170 V78 V170 3.12872492652814e-12
C78_170 V78 V170 7.24117245441997e-20

R78_171 V78 V171 158.40114910204665
L78_171 V78 V171 1.5910613623803697e-12
C78_171 V78 V171 3.0770003259702245e-19

R78_172 V78 V172 160.1381524061273
L78_172 V78 V172 1.5214723356323925e-12
C78_172 V78 V172 2.3633578410673016e-19

R78_173 V78 V173 -226.80898084599178
L78_173 V78 V173 -2.8769851183165586e-12
C78_173 V78 V173 -1.7574312227523403e-19

R78_174 V78 V174 -228.2379718692
L78_174 V78 V174 -5.700192192000985e-12
C78_174 V78 V174 -1.2611492402236223e-19

R78_175 V78 V175 -1535.2843675530437
L78_175 V78 V175 -3.1956947562367917e-11
C78_175 V78 V175 -9.73539365180156e-20

R78_176 V78 V176 -417.53870576300915
L78_176 V78 V176 -5.105175202231168e-12
C78_176 V78 V176 -1.3790788887779792e-19

R78_177 V78 V177 -223.01165755253066
L78_177 V78 V177 -6.528821760443613e-12
C78_177 V78 V177 9.852649644071199e-20

R78_178 V78 V178 -156.86062468672216
L78_178 V78 V178 -2.9933237221637226e-12
C78_178 V78 V178 -4.173763975530535e-20

R78_179 V78 V179 -440.57758767054804
L78_179 V78 V179 -2.247693560451156e-12
C78_179 V78 V179 -1.2499387625162861e-19

R78_180 V78 V180 -325.8078224321616
L78_180 V78 V180 -2.2169927313961347e-12
C78_180 V78 V180 -1.6574867643369545e-20

R78_181 V78 V181 191.35699813431106
L78_181 V78 V181 9.766168343525136e-12
C78_181 V78 V181 -9.075341701157891e-20

R78_182 V78 V182 93.35906893502708
L78_182 V78 V182 1.5047550715740735e-12
C78_182 V78 V182 1.1695999115495503e-19

R78_183 V78 V183 7592.84030879616
L78_183 V78 V183 -1.690733991485001e-11
C78_183 V78 V183 -2.2402143306169848e-20

R78_184 V78 V184 839.7487396022535
L78_184 V78 V184 6.773992680141293e-12
C78_184 V78 V184 -1.6912227688629062e-20

R78_185 V78 V185 833.8017608781661
L78_185 V78 V185 4.7657542233951064e-12
C78_185 V78 V185 -2.201302872332005e-20

R78_186 V78 V186 266.16004539078887
L78_186 V78 V186 2.519110868193235e-12
C78_186 V78 V186 -2.774217464892431e-20

R78_187 V78 V187 -12917.82073891338
L78_187 V78 V187 5.157013600212495e-12
C78_187 V78 V187 1.2874090340480024e-20

R78_188 V78 V188 -9453.24217540061
L78_188 V78 V188 5.877644765074295e-11
C78_188 V78 V188 3.50747054269424e-20

R78_189 V78 V189 -300.47105859109223
L78_189 V78 V189 -3.903128638041012e-11
C78_189 V78 V189 2.619928919427182e-19

R78_190 V78 V190 -138.12279126944233
L78_190 V78 V190 -2.2663981803616675e-12
C78_190 V78 V190 -1.2555845415887987e-19

R78_191 V78 V191 -1104.9392601500435
L78_191 V78 V191 3.5120525745535632e-12
C78_191 V78 V191 2.943699865832194e-19

R78_192 V78 V192 -659.2614537953872
L78_192 V78 V192 3.1628081032427395e-12
C78_192 V78 V192 3.0841497695765263e-19

R78_193 V78 V193 -1570.406705301133
L78_193 V78 V193 -3.751584058277913e-12
C78_193 V78 V193 -6.051047668196347e-20

R78_194 V78 V194 277.25188611340064
L78_194 V78 V194 3.6656059106362545e-12
C78_194 V78 V194 1.4353146008851504e-19

R78_195 V78 V195 1414.9237731734786
L78_195 V78 V195 -2.1071189575170327e-12
C78_195 V78 V195 -3.802225183769194e-19

R78_196 V78 V196 -7706.731761828268
L78_196 V78 V196 -1.3151770300639579e-12
C78_196 V78 V196 -5.18775206055885e-19

R78_197 V78 V197 579.6576421166544
L78_197 V78 V197 -3.805996361973618e-12
C78_197 V78 V197 -2.513621887658723e-19

R78_198 V78 V198 170.42139882622135
L78_198 V78 V198 2.844097748181587e-12
C78_198 V78 V198 6.505040477944944e-20

R78_199 V78 V199 1045.894188824131
L78_199 V78 V199 -2.0786858049673616e-12
C78_199 V78 V199 -1.8364865213159315e-19

R78_200 V78 V200 3350.229060080947
L78_200 V78 V200 -3.782881582868177e-12
C78_200 V78 V200 -7.519471238152828e-20

R79_79 V79 0 -150.14188851885825
L79_79 V79 0 -1.0601801160841083e-12
C79_79 V79 0 -6.066663394570023e-19

R79_80 V79 V80 -622.2301685764874
L79_80 V79 V80 6.348887060927028e-12
C79_80 V79 V80 1.0800090073469872e-19

R79_81 V79 V81 -385.42610875035
L79_81 V79 V81 3.682865959377512e-12
C79_81 V79 V81 1.301849310137116e-19

R79_82 V79 V82 1944.8605028193708
L79_82 V79 V82 -1.1542307448485722e-11
C79_82 V79 V82 -6.529775827869332e-20

R79_83 V79 V83 611.1911653821031
L79_83 V79 V83 3.0027987638362814e-12
C79_83 V79 V83 2.572944958417506e-19

R79_84 V79 V84 1396.126488641718
L79_84 V79 V84 -1.2055462438706107e-10
C79_84 V79 V84 -6.638063636840614e-20

R79_85 V79 V85 1865.5182540743629
L79_85 V79 V85 2.7462621754497967e-11
C79_85 V79 V85 6.636313409190652e-20

R79_86 V79 V86 310.42167820626906
L79_86 V79 V86 1.4035161441472543e-11
C79_86 V79 V86 -5.518322481778429e-21

R79_87 V79 V87 231.0776988422317
L79_87 V79 V87 1.4726076943103894e-12
C79_87 V79 V87 2.996006109430359e-19

R79_88 V79 V88 709.566532463676
L79_88 V79 V88 -4.702414282233977e-12
C79_88 V79 V88 -8.698725093082263e-20

R79_89 V79 V89 565.142912234089
L79_89 V79 V89 7.62041836746732e-12
C79_89 V79 V89 -3.4408693863172497e-20

R79_90 V79 V90 -435.5825457202868
L79_90 V79 V90 6.66677085337884e-12
C79_90 V79 V90 8.886675805329959e-20

R79_91 V79 V91 -152.8701195297464
L79_91 V79 V91 -1.2261039546944308e-12
C79_91 V79 V91 -3.7913850999174174e-19

R79_92 V79 V92 -782.7654389717168
L79_92 V79 V92 1.7888629551804793e-12
C79_92 V79 V92 2.2360365405965476e-19

R79_93 V79 V93 -673.3318260469044
L79_93 V79 V93 -9.965543151568321e-12
C79_93 V79 V93 -2.953734432974138e-20

R79_94 V79 V94 -687.9921883091952
L79_94 V79 V94 -1.6075759334968494e-11
C79_94 V79 V94 -1.308400829993047e-20

R79_95 V79 V95 -403.67404222946135
L79_95 V79 V95 1.4503578481469685e-11
C79_95 V79 V95 -1.3895423067458688e-20

R79_96 V79 V96 -650.7580983187264
L79_96 V79 V96 -3.605926829576855e-12
C79_96 V79 V96 -5.57209967475601e-20

R79_97 V79 V97 -1706.0452645837197
L79_97 V79 V97 -5.8787942536374575e-12
C79_97 V79 V97 -3.823394640287718e-20

R79_98 V79 V98 391.5256007490605
L79_98 V79 V98 -4.5211559232759674e-10
C79_98 V79 V98 -2.920959289473847e-20

R79_99 V79 V99 122.51710384662623
L79_99 V79 V99 1.7565168203178769e-12
C79_99 V79 V99 2.9614904485592286e-19

R79_100 V79 V100 673.9008306502212
L79_100 V79 V100 -3.6225330574332466e-12
C79_100 V79 V100 -1.8860256304525453e-19

R79_101 V79 V101 -5001.592971585537
L79_101 V79 V101 8.81410143387576e-12
C79_101 V79 V101 6.089651772290119e-20

R79_102 V79 V102 2881.070603782801
L79_102 V79 V102 7.565893698891931e-10
C79_102 V79 V102 -9.782389816065038e-21

R79_103 V79 V103 -740.9486164286053
L79_103 V79 V103 -1.6016140001723155e-12
C79_103 V79 V103 -2.31116194439334e-19

R79_104 V79 V104 640.7883830591301
L79_104 V79 V104 3.483710068628303e-12
C79_104 V79 V104 6.953852728416761e-20

R79_105 V79 V105 976.1898457707047
L79_105 V79 V105 1.2024021988794898e-11
C79_105 V79 V105 7.529960652449356e-20

R79_106 V79 V106 2849.4854572329004
L79_106 V79 V106 6.460408553069625e-12
C79_106 V79 V106 1.0707600740943927e-19

R79_107 V79 V107 -192.07990710363825
L79_107 V79 V107 1.4398748628496873e-11
C79_107 V79 V107 2.182020590425655e-20

R79_108 V79 V108 -707.9588236570924
L79_108 V79 V108 -1.631011031620225e-11
C79_108 V79 V108 8.695444424759296e-20

R79_109 V79 V109 962.351504694005
L79_109 V79 V109 1.6800915028714506e-11
C79_109 V79 V109 -2.1964799348861436e-20

R79_110 V79 V110 -703.3866007814294
L79_110 V79 V110 -1.1330588700956815e-11
C79_110 V79 V110 -6.976867216869687e-20

R79_111 V79 V111 274.60727467898386
L79_111 V79 V111 5.043073921944984e-12
C79_111 V79 V111 4.0455403308983886e-20

R79_112 V79 V112 9857.095572969763
L79_112 V79 V112 2.616332276721368e-12
C79_112 V79 V112 1.3701905412876476e-19

R79_113 V79 V113 -245.64657798714615
L79_113 V79 V113 -5.030796951715721e-12
C79_113 V79 V113 -1.1180969517942221e-19

R79_114 V79 V114 -1107.5924387855407
L79_114 V79 V114 -7.311597144189683e-12
C79_114 V79 V114 -9.486888166917971e-20

R79_115 V79 V115 459.65177344482726
L79_115 V79 V115 3.794455398288569e-12
C79_115 V79 V115 5.060774398296861e-20

R79_116 V79 V116 1236.619991885826
L79_116 V79 V116 -2.1911309882616826e-12
C79_116 V79 V116 -2.2250248270056914e-19

R79_117 V79 V117 -903.0228507650678
L79_117 V79 V117 -2.2564072074172178e-10
C79_117 V79 V117 5.0256431484295334e-20

R79_118 V79 V118 287.4636138022758
L79_118 V79 V118 3.8532602454947655e-12
C79_118 V79 V118 1.26944903189555e-19

R79_119 V79 V119 -470.87539589734644
L79_119 V79 V119 2.1020506850924732e-11
C79_119 V79 V119 -6.545576957089569e-21

R79_120 V79 V120 -8072.478248194588
L79_120 V79 V120 -4.266754445577821e-11
C79_120 V79 V120 1.1698134975232408e-21

R79_121 V79 V121 252.04190562256844
L79_121 V79 V121 3.54067145247154e-11
C79_121 V79 V121 3.4536447601551686e-20

R79_122 V79 V122 -1318.072492104689
L79_122 V79 V122 -3.8618657440082573e-11
C79_122 V79 V122 1.3710562988713205e-22

R79_123 V79 V123 988.8989811110189
L79_123 V79 V123 -1.2274050704633706e-12
C79_123 V79 V123 -3.5112228351122834e-19

R79_124 V79 V124 23067.778959319214
L79_124 V79 V124 1.5911321907051302e-12
C79_124 V79 V124 2.937515845528158e-19

R79_125 V79 V125 840.9479426386312
L79_125 V79 V125 4.485397871207542e-12
C79_125 V79 V125 2.9360368286602105e-20

R79_126 V79 V126 -304.9765861846251
L79_126 V79 V126 -4.9861538068689255e-12
C79_126 V79 V126 -1.0480407372000141e-19

R79_127 V79 V127 -446.6742221875116
L79_127 V79 V127 1.3054040035027892e-12
C79_127 V79 V127 4.1657125561374224e-19

R79_128 V79 V128 -1545.372921049049
L79_128 V79 V128 -3.2819430136462386e-12
C79_128 V79 V128 -1.638011319349127e-19

R79_129 V79 V129 -184.8075440798644
L79_129 V79 V129 -9.041918839890137e-12
C79_129 V79 V129 -1.5784483494320287e-21

R79_130 V79 V130 574.9696047028505
L79_130 V79 V130 2.7500988884158248e-11
C79_130 V79 V130 -1.5138537362432627e-20

R79_131 V79 V131 337.79278815160245
L79_131 V79 V131 -1.6120968336142195e-11
C79_131 V79 V131 -1.2011927056156638e-19

R79_132 V79 V132 567.5260763477429
L79_132 V79 V132 2.934254246817309e-11
C79_132 V79 V132 -1.0831740021388273e-20

R79_133 V79 V133 -4468.589358022332
L79_133 V79 V133 -1.2305239482123914e-11
C79_133 V79 V133 -6.661585121344884e-20

R79_134 V79 V134 1623.4733341670774
L79_134 V79 V134 1.090305356660508e-11
C79_134 V79 V134 7.991357282701548e-20

R79_135 V79 V135 260.9330057889031
L79_135 V79 V135 -9.86759087149084e-13
C79_135 V79 V135 -5.651970200296249e-19

R79_136 V79 V136 1054.3643984374307
L79_136 V79 V136 2.170305030314167e-12
C79_136 V79 V136 3.1858444677994733e-19

R79_137 V79 V137 235.12903273903666
L79_137 V79 V137 -5.790295877453254e-12
C79_137 V79 V137 -7.736401023486699e-20

R79_138 V79 V138 -640.4380596908034
L79_138 V79 V138 -4.9151678228403e-12
C79_138 V79 V138 -1.113612532674583e-19

R79_139 V79 V139 -134.24905712279363
L79_139 V79 V139 6.797341953090504e-13
C79_139 V79 V139 7.965280790352372e-19

R79_140 V79 V140 -273.5516946943131
L79_140 V79 V140 -1.5665044797376665e-12
C79_140 V79 V140 -4.0665527963637784e-19

R79_141 V79 V141 462.4237597547728
L79_141 V79 V141 4.314111488601e-12
C79_141 V79 V141 1.549810080697656e-19

R79_142 V79 V142 -2258.2497786088848
L79_142 V79 V142 2.2921682712885153e-11
C79_142 V79 V142 1.9797718288133614e-20

R79_143 V79 V143 13714.950026977174
L79_143 V79 V143 -5.74933054755802e-12
C79_143 V79 V143 -1.2760530911906985e-19

R79_144 V79 V144 1152.5887126976836
L79_144 V79 V144 1.2303795525080959e-11
C79_144 V79 V144 1.0974893001820212e-19

R79_145 V79 V145 -179.78106784881336
L79_145 V79 V145 3.4048358033618186e-12
C79_145 V79 V145 6.440030190597383e-20

R79_146 V79 V146 1066.637431946331
L79_146 V79 V146 1.0084192566256767e-11
C79_146 V79 V146 1.3113427458693783e-21

R79_147 V79 V147 286.9767246558976
L79_147 V79 V147 -1.5568969766834085e-12
C79_147 V79 V147 -3.791722281138736e-19

R79_148 V79 V148 3090.4654878839083
L79_148 V79 V148 1.1167452526343422e-12
C79_148 V79 V148 2.6482894691722635e-19

R79_149 V79 V149 -907.2557364333239
L79_149 V79 V149 -2.717197651174872e-12
C79_149 V79 V149 -8.605885311714722e-20

R79_150 V79 V150 341.9792039218574
L79_150 V79 V150 1.599428315347004e-11
C79_150 V79 V150 1.5614092930688737e-19

R79_151 V79 V151 235.90795391017252
L79_151 V79 V151 6.6758943191873015e-12
C79_151 V79 V151 2.5286541818156867e-19

R79_152 V79 V152 -693.2583706541058
L79_152 V79 V152 -2.0379999570064035e-12
C79_152 V79 V152 -1.241305807614697e-19

R79_153 V79 V153 419.43151261219424
L79_153 V79 V153 -2.74435681033105e-12
C79_153 V79 V153 -1.694454600201456e-19

R79_154 V79 V154 -11938.252913533868
L79_154 V79 V154 -3.57832522494667e-12
C79_154 V79 V154 -1.197915481090246e-19

R79_155 V79 V155 -161.5266559978199
L79_155 V79 V155 1.2363304628543761e-12
C79_155 V79 V155 1.155852358076769e-19

R79_156 V79 V156 392.1150325036143
L79_156 V79 V156 -4.414546931588255e-12
C79_156 V79 V156 -2.0194551259470676e-19

R79_157 V79 V157 216.41846107082526
L79_157 V79 V157 2.03702354459164e-12
C79_157 V79 V157 1.4751727844128793e-19

R79_158 V79 V158 24741.20584067331
L79_158 V79 V158 7.148669908168611e-12
C79_158 V79 V158 2.005354945929213e-20

R79_159 V79 V159 -1089.6888579382635
L79_159 V79 V159 -1.4195958944238571e-12
C79_159 V79 V159 -3.1046323053331535e-19

R79_160 V79 V160 615.542902835126
L79_160 V79 V160 5.9533208642999224e-12
C79_160 V79 V160 1.244515730103758e-19

R79_161 V79 V161 -238.6204771802384
L79_161 V79 V161 -1.7390731487854323e-11
C79_161 V79 V161 1.3759969796755366e-19

R79_162 V79 V162 -581.2501625081096
L79_162 V79 V162 -4.209486956657026e-10
C79_162 V79 V162 1.229258865367941e-20

R79_163 V79 V163 -370.6839389396241
L79_163 V79 V163 -2.175205844648587e-12
C79_163 V79 V163 1.3295618866566346e-19

R79_164 V79 V164 -288.08324190221606
L79_164 V79 V164 -2.891758279553122e-11
C79_164 V79 V164 -5.227118198481939e-20

R79_165 V79 V165 -335.49423822970647
L79_165 V79 V165 -1.6206970209411762e-11
C79_165 V79 V165 -5.536812611438707e-20

R79_166 V79 V166 1188.2062763105882
L79_166 V79 V166 9.645133763382933e-12
C79_166 V79 V166 1.0056071745058413e-19

R79_167 V79 V167 171.26147243999674
L79_167 V79 V167 1.3449821741691423e-12
C79_167 V79 V167 1.0402361397664816e-19

R79_168 V79 V168 -524.4755574662335
L79_168 V79 V168 -6.916711510631516e-12
C79_168 V79 V168 1.275685754069097e-19

R79_169 V79 V169 253.2463759814153
L79_169 V79 V169 -2.910793210054251e-12
C79_169 V79 V169 -1.933091555290653e-19

R79_170 V79 V170 739.8883953970858
L79_170 V79 V170 -5.189816529265379e-12
C79_170 V79 V170 -8.352083329669202e-20

R79_171 V79 V171 1633.8238230000188
L79_171 V79 V171 -3.5390727359681513e-12
C79_171 V79 V171 -1.8870946594258996e-19

R79_172 V79 V172 377.4294035610075
L79_172 V79 V172 4.3512756899894145e-12
C79_172 V79 V172 -9.144863288284503e-20

R79_173 V79 V173 3221.0792509896633
L79_173 V79 V173 3.3980337366233497e-12
C79_173 V79 V173 1.0790386309989511e-19

R79_174 V79 V174 -1417.8688919808653
L79_174 V79 V174 -4.9654855511790255e-12
C79_174 V79 V174 -5.230947064157782e-20

R79_175 V79 V175 -253.7032805951893
L79_175 V79 V175 1.0169920225991367e-11
C79_175 V79 V175 2.1263007294415628e-19

R79_176 V79 V176 -1296.9701361394928
L79_176 V79 V176 -1.892770039556765e-12
C79_176 V79 V176 -2.3955869571143825e-19

R79_177 V79 V177 -457.66392840631664
L79_177 V79 V177 -1.1943553555131004e-11
C79_177 V79 V177 5.472842858530173e-20

R79_178 V79 V178 -1542.8991540713437
L79_178 V79 V178 4.282198403926474e-12
C79_178 V79 V178 3.4744610758361293e-20

R79_179 V79 V179 -463.50644882458715
L79_179 V79 V179 3.5654122393146003e-11
C79_179 V79 V179 -1.0698078716345677e-19

R79_180 V79 V180 -2023.2497454826594
L79_180 V79 V180 3.655422265474772e-12
C79_180 V79 V180 1.978076269597943e-19

R79_181 V79 V181 682.4958202814292
L79_181 V79 V181 5.0781071131374294e-11
C79_181 V79 V181 5.468079145135257e-20

R79_182 V79 V182 717.008910789776
L79_182 V79 V182 7.551546466161093e-12
C79_182 V79 V182 4.2222244461983046e-20

R79_183 V79 V183 200.97793071086733
L79_183 V79 V183 -6.9331597708875744e-12
C79_183 V79 V183 1.7497267982695887e-20

R79_184 V79 V184 1121.4376493995087
L79_184 V79 V184 9.371792809840494e-12
C79_184 V79 V184 -7.641675977004677e-20

R79_185 V79 V185 686.9906734654752
L79_185 V79 V185 2.4381281035214742e-12
C79_185 V79 V185 -6.099571837138626e-20

R79_186 V79 V186 3786.345003537016
L79_186 V79 V186 -5.161048547326659e-12
C79_186 V79 V186 -2.8538221230131267e-20

R79_187 V79 V187 -1127.0413381090978
L79_187 V79 V187 1.6974388925147704e-12
C79_187 V79 V187 1.3964012374134625e-19

R79_188 V79 V188 -491.26014690783734
L79_188 V79 V188 -2.2851736428581433e-12
C79_188 V79 V188 1.9880011784518865e-21

R79_189 V79 V189 -746.364884479391
L79_189 V79 V189 -2.301843309608325e-12
C79_189 V79 V189 -9.666043790477425e-20

R79_190 V79 V190 -1933.2918277355682
L79_190 V79 V190 2.703289253218004e-11
C79_190 V79 V190 3.9860904028781464e-20

R79_191 V79 V191 -268.1333561481898
L79_191 V79 V191 -2.4100869039050164e-12
C79_191 V79 V191 -2.0334278956801412e-19

R79_192 V79 V192 -3533.0547017895497
L79_192 V79 V192 2.468276129825985e-12
C79_192 V79 V192 3.679087080117539e-20

R79_193 V79 V193 -948.9492199076328
L79_193 V79 V193 -4.3285023729017475e-12
C79_193 V79 V193 2.770249238373236e-20

R79_194 V79 V194 963.5863750617864
L79_194 V79 V194 -2.5952773509235526e-11
C79_194 V79 V194 -9.430572569811004e-20

R79_195 V79 V195 293.7070142556614
L79_195 V79 V195 1.395775599377963e-12
C79_195 V79 V195 4.378421384056352e-19

R79_196 V79 V196 538.0071624617397
L79_196 V79 V196 -1.6654792464331163e-12
C79_196 V79 V196 -2.7170066110752743e-19

R79_197 V79 V197 793.5074270319803
L79_197 V79 V197 3.1812801864856274e-12
C79_197 V79 V197 8.292281555251904e-20

R79_198 V79 V198 849.9487277781635
L79_198 V79 V198 -2.4443033450180674e-11
C79_198 V79 V198 5.494559527278667e-20

R79_199 V79 V199 427.79863135770785
L79_199 V79 V199 -5.733004037015008e-12
C79_199 V79 V199 -6.411840141702021e-20

R79_200 V79 V200 -2022.6811008282202
L79_200 V79 V200 9.916831366165097e-12
C79_200 V79 V200 1.5385667444343088e-19

R80_80 V80 0 -102.87116184834247
L80_80 V80 0 5.070121176475902e-13
C80_80 V80 0 8.684229603213032e-19

R80_81 V80 V81 -290.5805210612846
L80_81 V80 V81 1.1986076750834356e-11
C80_81 V80 V81 4.950097793841411e-21

R80_82 V80 V82 1094.9483800557293
L80_82 V80 V82 -2.428450158366084e-12
C80_82 V80 V82 -2.8083073146416544e-19

R80_83 V80 V83 976.5732574752774
L80_83 V80 V83 -1.538765034891616e-11
C80_83 V80 V83 -1.0894815927379044e-19

R80_84 V80 V84 769.0955818356834
L80_84 V80 V84 1.6728918196480711e-10
C80_84 V80 V84 1.5803294438245967e-19

R80_85 V80 V85 1817.647516348918
L80_85 V80 V85 -6.881734173803321e-12
C80_85 V80 V85 1.6329983260239596e-20

R80_86 V80 V86 269.06418860049314
L80_86 V80 V86 -2.0051296116314247e-11
C80_86 V80 V86 -5.695592774599924e-20

R80_87 V80 V87 543.3098851799725
L80_87 V80 V87 7.265024669784601e-12
C80_87 V80 V87 2.8758204626854436e-20

R80_88 V80 V88 187.32914297547032
L80_88 V80 V88 7.225209981886001e-13
C80_88 V80 V88 5.330295535744228e-19

R80_89 V80 V89 399.1934306094778
L80_89 V80 V89 1.2998924068474635e-12
C80_89 V80 V89 1.9557332068110111e-19

R80_90 V80 V90 -360.4799130482649
L80_90 V80 V90 9.067863150051402e-13
C80_90 V80 V90 4.685415079980388e-19

R80_91 V80 V91 -376.8393399562141
L80_91 V80 V91 9.525348187653208e-11
C80_91 V80 V91 6.302548399732779e-20

R80_92 V80 V92 -127.98980425754534
L80_92 V80 V92 -5.859026341141734e-13
C80_92 V80 V92 -5.957028353538792e-19

R80_93 V80 V93 -607.4321675583753
L80_93 V80 V93 -1.0406172846121717e-11
C80_93 V80 V93 -5.915754995180086e-20

R80_94 V80 V94 -979.7728209695758
L80_94 V80 V94 -2.9676135353081456e-12
C80_94 V80 V94 -2.210621833748571e-19

R80_95 V80 V95 -873.2883084251245
L80_95 V80 V95 -4.972416263741597e-12
C80_95 V80 V95 -1.0008064342782298e-19

R80_96 V80 V96 -431.6409568056082
L80_96 V80 V96 2.791209684880026e-12
C80_96 V80 V96 -4.7874593808382665e-20

R80_97 V80 V97 -1758.4814958090028
L80_97 V80 V97 -1.1445463631631847e-12
C80_97 V80 V97 -3.798257971509347e-19

R80_98 V80 V98 450.99851754199295
L80_98 V80 V98 -1.6234747398975554e-12
C80_98 V80 V98 -2.51509682009528e-19

R80_99 V80 V99 310.98336362722284
L80_99 V80 V99 2.3691472562561224e-12
C80_99 V80 V99 4.3378840095116104e-20

R80_100 V80 V100 112.4372878103341
L80_100 V80 V100 1.1651970038778734e-12
C80_100 V80 V100 4.8020273981472205e-19

R80_101 V80 V101 -2313.304940282193
L80_101 V80 V101 1.8404749832013627e-12
C80_101 V80 V101 1.9864232679135804e-19

R80_102 V80 V102 3641.3493619102137
L80_102 V80 V102 2.2655172155713138e-12
C80_102 V80 V102 2.0501435826801097e-19

R80_103 V80 V103 1180.9675590564286
L80_103 V80 V103 2.193528464768028e-11
C80_103 V80 V103 3.055980836373982e-20

R80_104 V80 V104 -1835.7835363124168
L80_104 V80 V104 -1.1758849008207258e-12
C80_104 V80 V104 -2.691030544779933e-19

R80_105 V80 V105 703.704230277629
L80_105 V80 V105 2.498123621842719e-12
C80_105 V80 V105 2.201462746359465e-19

R80_106 V80 V106 993.3340786494442
L80_106 V80 V106 2.6348198299941152e-12
C80_106 V80 V106 1.5677995069863995e-19

R80_107 V80 V107 -382.2397565576218
L80_107 V80 V107 -3.4866828178863258e-12
C80_107 V80 V107 -5.156479738968286e-20

R80_108 V80 V108 -142.66357742486366
L80_108 V80 V108 2.9575141227501216e-12
C80_108 V80 V108 4.536806915844522e-20

R80_109 V80 V109 907.0710612832492
L80_109 V80 V109 -3.7264564338093946e-12
C80_109 V80 V109 -2.755127593502519e-19

R80_110 V80 V110 -421.58579747502915
L80_110 V80 V110 -5.6006360505455805e-12
C80_110 V80 V110 -9.130845596340457e-20

R80_111 V80 V111 2527.241826178162
L80_111 V80 V111 6.2752920667302235e-12
C80_111 V80 V111 5.467557166592389e-20

R80_112 V80 V112 293.1546581100187
L80_112 V80 V112 -1.949554460078934e-12
C80_112 V80 V112 -2.014836123235681e-19

R80_113 V80 V113 -189.00026373981964
L80_113 V80 V113 -1.931914213448933e-12
C80_113 V80 V113 -1.7530639786848362e-19

R80_114 V80 V114 -1004.7653112708842
L80_114 V80 V114 -1.5626458334000313e-12
C80_114 V80 V114 -2.56245158616903e-19

R80_115 V80 V115 654.6557650282168
L80_115 V80 V115 1.8023001755662073e-10
C80_115 V80 V115 -5.560582512379252e-20

R80_116 V80 V116 185.07185768219438
L80_116 V80 V116 1.5735897574517337e-12
C80_116 V80 V116 1.301855162801184e-19

R80_117 V80 V117 -2359.6858626827675
L80_117 V80 V117 2.7201526621597765e-12
C80_117 V80 V117 2.390917922603992e-19

R80_118 V80 V118 191.96177164542436
L80_118 V80 V118 1.4772323749549575e-12
C80_118 V80 V118 3.2622067700505794e-19

R80_119 V80 V119 -4039.3332135889955
L80_119 V80 V119 4.573325408999838e-12
C80_119 V80 V119 2.246059452602081e-19

R80_120 V80 V120 -153.29665986184486
L80_120 V80 V120 2.6363230823280823e-12
C80_120 V80 V120 3.642211146707709e-19

R80_121 V80 V121 239.21104082977806
L80_121 V80 V121 5.455201054829306e-12
C80_121 V80 V121 -4.160449323659763e-21

R80_122 V80 V122 -441.97587955246735
L80_122 V80 V122 -4.743585838758589e-11
C80_122 V80 V122 -5.2468436293121476e-21

R80_123 V80 V123 -1767.762127870158
L80_123 V80 V123 -1.1832161904522736e-11
C80_123 V80 V123 -2.9852440955439324e-20

R80_124 V80 V124 476.2562455740846
L80_124 V80 V124 -6.084606148635378e-13
C80_124 V80 V124 -7.788612955553219e-19

R80_125 V80 V125 -12936.526289362118
L80_125 V80 V125 -2.416967198304447e-11
C80_125 V80 V125 -2.4224101133159284e-20

R80_126 V80 V126 -192.9340491790421
L80_126 V80 V126 -1.2546642466063187e-12
C80_126 V80 V126 -2.271124301614979e-19

R80_127 V80 V127 -521.3219480101691
L80_127 V80 V127 -1.5829982296336045e-12
C80_127 V80 V127 -3.4061726934914836e-19

R80_128 V80 V128 1620.1608528604052
L80_128 V80 V128 1.2513948747029099e-12
C80_128 V80 V128 1.9993519733008564e-19

R80_129 V80 V129 -201.74840684689948
L80_129 V80 V129 -2.8665074468125288e-12
C80_129 V80 V129 -2.0236773624773678e-19

R80_130 V80 V130 250.88171123049315
L80_130 V80 V130 1.875043772989792e-12
C80_130 V80 V130 1.5122479985828512e-19

R80_131 V80 V131 346.7567084929257
L80_131 V80 V131 1.7605569927863419e-12
C80_131 V80 V131 2.687328398675836e-19

R80_132 V80 V132 802.2975937338416
L80_132 V80 V132 1.4137873456246268e-12
C80_132 V80 V132 4.0994795619486107e-19

R80_133 V80 V133 11006.892780383925
L80_133 V80 V133 2.7853598132238905e-12
C80_133 V80 V133 2.6793042953150815e-19

R80_134 V80 V134 -5169.504671206851
L80_134 V80 V134 2.5986969902521845e-11
C80_134 V80 V134 1.6112696361393872e-19

R80_135 V80 V135 3578.26365029532
L80_135 V80 V135 2.5310291932103863e-12
C80_135 V80 V135 2.993472707134014e-19

R80_136 V80 V136 216.13519874837755
L80_136 V80 V136 -7.460531350862154e-13
C80_136 V80 V136 -7.644105335830332e-19

R80_137 V80 V137 241.70593988010486
L80_137 V80 V137 -8.936725602688631e-12
C80_137 V80 V137 -6.4551941071147e-20

R80_138 V80 V138 -578.8998263610805
L80_138 V80 V138 -1.9621932324327223e-12
C80_138 V80 V138 -2.4203758749174793e-19

R80_139 V80 V139 -321.70786082571175
L80_139 V80 V139 -1.4242416259761322e-12
C80_139 V80 V139 -4.0783811409729607e-19

R80_140 V80 V140 -108.87987800715683
L80_140 V80 V140 1.0090443745469706e-12
C80_140 V80 V140 7.855708507680315e-19

R80_141 V80 V141 548.9530773457623
L80_141 V80 V141 -1.993551166760584e-12
C80_141 V80 V141 -2.0547629595434884e-19

R80_142 V80 V142 -5037.60736525976
L80_142 V80 V142 2.188220608236595e-11
C80_142 V80 V142 5.098995196945774e-21

R80_143 V80 V143 686.7604792094504
L80_143 V80 V143 -5.227260333801433e-12
C80_143 V80 V143 -1.2517558185686008e-20

R80_144 V80 V144 -12338.031913294568
L80_144 V80 V144 9.493854811280487e-12
C80_144 V80 V144 -1.0543409314265078e-19

R80_145 V80 V145 -185.17407637860188
L80_145 V80 V145 3.450755525421108e-12
C80_145 V80 V145 5.058640332006166e-20

R80_146 V80 V146 1045.4526230585673
L80_146 V80 V146 2.3243299510152855e-12
C80_146 V80 V146 1.0592421164019486e-19

R80_147 V80 V147 23611.072016460937
L80_147 V80 V147 4.383752411666575e-12
C80_147 V80 V147 5.920466891294338e-20

R80_148 V80 V148 171.78558449479254
L80_148 V80 V148 -5.718859002510725e-13
C80_148 V80 V148 -6.115963326216362e-19

R80_149 V80 V149 -673.6127210199938
L80_149 V80 V149 2.0068580423248034e-12
C80_149 V80 V149 2.635226506132555e-19

R80_150 V80 V150 331.16532675430506
L80_150 V80 V150 -6.78113671066677e-12
C80_150 V80 V150 -1.1818831799552224e-19

R80_151 V80 V151 2012.1585250880378
L80_151 V80 V151 4.204171857127954e-12
C80_151 V80 V151 2.3302764092107268e-20

R80_152 V80 V152 10318.825018263893
L80_152 V80 V152 1.274201964514137e-12
C80_152 V80 V152 2.6579915612897845e-19

R80_153 V80 V153 339.9541419185441
L80_153 V80 V153 5.34109863214216e-12
C80_153 V80 V153 -5.161976368250389e-20

R80_154 V80 V154 7017.305849522529
L80_154 V80 V154 2.2102068231540935e-11
C80_154 V80 V154 2.6254705557467478e-20

R80_155 V80 V155 -4950.038653041884
L80_155 V80 V155 1.0906360337747804e-11
C80_155 V80 V155 -5.248889541937647e-20

R80_156 V80 V156 2010.5439419510685
L80_156 V80 V156 1.2070294904645156e-12
C80_156 V80 V156 4.1293146440458554e-19

R80_157 V80 V157 189.6724411715429
L80_157 V80 V157 -1.2174776529929053e-12
C80_157 V80 V157 -3.3713812805547403e-19

R80_158 V80 V158 4396.037523857537
L80_158 V80 V158 1.476271946407517e-11
C80_158 V80 V158 3.456579863091451e-20

R80_159 V80 V159 359.24862853045124
L80_159 V80 V159 4.18806893371799e-12
C80_159 V80 V159 1.3401545344854683e-19

R80_160 V80 V160 -313.73057768798213
L80_160 V80 V160 -1.5213557676578337e-12
C80_160 V80 V160 -3.829202736770409e-19

R80_161 V80 V161 -227.9205678844568
L80_161 V80 V161 2.2790850576480208e-12
C80_161 V80 V161 1.6939065966378202e-19

R80_162 V80 V162 -442.59271008429096
L80_162 V80 V162 2.5075371745445357e-12
C80_162 V80 V162 4.575493902708651e-20

R80_163 V80 V163 -238.7633582174692
L80_163 V80 V163 -2.7124329510332173e-12
C80_163 V80 V163 -1.3623626403277554e-19

R80_164 V80 V164 -238.3951390645241
L80_164 V80 V164 -2.190809405397098e-12
C80_164 V80 V164 2.3671048928200875e-19

R80_165 V80 V165 -275.06853650455724
L80_165 V80 V165 1.2024305349702676e-08
C80_165 V80 V165 6.456396356624707e-20

R80_166 V80 V166 1900.2914147769025
L80_166 V80 V166 -3.4302133458107265e-12
C80_166 V80 V166 -6.153298216910529e-20

R80_167 V80 V167 1035.1737247056994
L80_167 V80 V167 4.649836928506339e-11
C80_167 V80 V167 1.0408478960542992e-19

R80_168 V80 V168 229.68793365019437
L80_168 V80 V168 9.04711524871999e-13
C80_168 V80 V168 -1.1285954472297279e-20

R80_169 V80 V169 207.65568526787814
L80_169 V80 V169 -3.626034261923202e-12
C80_169 V80 V169 -2.847027420565764e-19

R80_170 V80 V170 298.6612879524619
L80_170 V80 V170 3.260039978708937e-12
C80_170 V80 V170 5.758084553706486e-20

R80_171 V80 V171 316.0381916134371
L80_171 V80 V171 1.3370077388126469e-12
C80_171 V80 V171 7.15958934926829e-20

R80_172 V80 V172 278.4271871908515
L80_172 V80 V172 -1.3533964360572977e-12
C80_172 V80 V172 -9.644826077719593e-20

R80_173 V80 V173 1705.2110154448499
L80_173 V80 V173 3.9509810031565995e-12
C80_173 V80 V173 1.2589390949977266e-19

R80_174 V80 V174 -717.4161855949119
L80_174 V80 V174 -2.6160265318881787e-12
C80_174 V80 V174 -1.3084900007234717e-19

R80_175 V80 V175 -875.3244297133382
L80_175 V80 V175 -1.6711054225678421e-12
C80_175 V80 V175 -1.0980931980505752e-19

R80_176 V80 V176 -197.2912781492906
L80_176 V80 V176 1.8259668370686765e-12
C80_176 V80 V176 3.922988104766941e-19

R80_177 V80 V177 -325.9690132344151
L80_177 V80 V177 -3.591916686780062e-12
C80_177 V80 V177 3.9090171934629625e-20

R80_178 V80 V178 -435.6762444079382
L80_178 V80 V178 -1.0261263187937646e-11
C80_178 V80 V178 -2.036431747071996e-20

R80_179 V80 V179 -999.1925914403073
L80_179 V80 V179 -2.9994574308985728e-12
C80_179 V80 V179 -8.73331747383532e-20

R80_180 V80 V180 -226.70171253544353
L80_180 V80 V180 -1.674180988184941e-12
C80_180 V80 V180 -3.585102062085266e-19

R80_181 V80 V181 510.88922174455115
L80_181 V80 V181 1.8918067836134248e-11
C80_181 V80 V181 -2.4624377672637777e-20

R80_182 V80 V182 265.76792819796583
L80_182 V80 V182 2.1730520766925815e-12
C80_182 V80 V182 5.501781152438398e-20

R80_183 V80 V183 2503.4908049039936
L80_183 V80 V183 -3.2434540975236945e-12
C80_183 V80 V183 -1.033524616631934e-19

R80_184 V80 V184 191.04431126797596
L80_184 V80 V184 -3.217824688540402e-12
C80_184 V80 V184 5.997460649281235e-20

R80_185 V80 V185 452.6259918934387
L80_185 V80 V185 1.8568223648784927e-12
C80_185 V80 V185 5.087835178446988e-21

R80_186 V80 V186 1937.9672553627995
L80_186 V80 V186 -2.485474098240251e-12
C80_186 V80 V186 4.494732204814535e-20

R80_187 V80 V187 -763.2333060377728
L80_187 V80 V187 2.3370922305195387e-11
C80_187 V80 V187 1.3770553490513613e-19

R80_188 V80 V188 1076.2236446047261
L80_188 V80 V188 6.039174255438417e-13
C80_188 V80 V188 2.0320035325862333e-19

R80_189 V80 V189 -510.7838260043153
L80_189 V80 V189 -2.2625442085040324e-12
C80_189 V80 V189 -1.4437509610702602e-21

R80_190 V80 V190 -544.483718622771
L80_190 V80 V190 1.77031337269272e-11
C80_190 V80 V190 -5.1728198666134584e-20

R80_191 V80 V191 2023.2221578624244
L80_191 V80 V191 9.899824361338498e-13
C80_191 V80 V191 1.9773632897029628e-19

R80_192 V80 V192 -194.18391102587367
L80_192 V80 V192 -1.1576406398462757e-12
C80_192 V80 V192 -2.2359397877379226e-19

R80_193 V80 V193 -602.5312354037835
L80_193 V80 V193 -2.0645783931244004e-12
C80_193 V80 V193 -9.992829063300404e-20

R80_194 V80 V194 714.0346668371185
L80_194 V80 V194 -2.6380017308264297e-12
C80_194 V80 V194 -2.68383085046726e-19

R80_195 V80 V195 1949.7152203783658
L80_195 V80 V195 -8.042046236590329e-13
C80_195 V80 V195 -4.885599079582937e-19

R80_196 V80 V196 276.0475459490693
L80_196 V80 V196 1.3946659979820386e-12
C80_196 V80 V196 4.693061893557223e-19

R80_197 V80 V197 737.6656866133148
L80_197 V80 V197 4.093970583377088e-12
C80_197 V80 V197 7.42753342651447e-20

R80_198 V80 V198 488.3943608958003
L80_198 V80 V198 5.0005829446338555e-11
C80_198 V80 V198 -7.555490977200828e-21

R80_199 V80 V199 895.8841943916277
L80_199 V80 V199 -8.349144510045714e-12
C80_199 V80 V199 3.6488672011227105e-20

R80_200 V80 V200 542.1477565136396
L80_200 V80 V200 -2.623615538788903e-12
C80_200 V80 V200 -1.826983538565587e-19

R81_81 V81 0 134.77269375403438
L81_81 V81 0 2.3616982528993346e-13
C81_81 V81 0 1.1427402136669286e-18

R81_82 V81 V82 546.6669505155057
L81_82 V81 V82 -4.524541146193708e-12
C81_82 V81 V82 -1.285710609245077e-19

R81_83 V81 V83 338.2450817752871
L81_83 V81 V83 7.636528468191658e-11
C81_83 V81 V83 2.7749044575058483e-20

R81_84 V81 V84 463.8578788309202
L81_84 V81 V84 -7.367004037086131e-12
C81_84 V81 V84 -4.452256614245442e-20

R81_85 V81 V85 473.9997599226878
L81_85 V81 V85 2.0984363067496407e-12
C81_85 V81 V85 2.544786687864454e-19

R81_86 V81 V86 152.00307266445859
L81_86 V81 V86 1.542298232923401e-11
C81_86 V81 V86 1.384933379840545e-20

R81_87 V81 V87 435.1255617740129
L81_87 V81 V87 -1.3191371156414366e-11
C81_87 V81 V87 -1.3520906645734935e-19

R81_88 V81 V88 320.2016051086763
L81_88 V81 V88 5.2388296339793554e-11
C81_88 V81 V88 -6.009935894510185e-20

R81_89 V81 V89 171.86320064459596
L81_89 V81 V89 -1.582812066819065e-12
C81_89 V81 V89 -2.29332710815728e-19

R81_90 V81 V90 -170.46856808126924
L81_90 V81 V90 3.4019144880085475e-11
C81_90 V81 V90 4.374357581693119e-20

R81_91 V81 V91 -179.10091201059657
L81_91 V81 V91 -2.5496679845661996e-12
C81_91 V81 V91 -1.1077469601168873e-19

R81_92 V81 V92 -216.70728395087133
L81_92 V81 V92 -4.072315146140415e-12
C81_92 V81 V92 -6.758261817069692e-20

R81_93 V81 V93 -111.2817169423738
L81_93 V81 V93 5.2073274405735426e-12
C81_93 V81 V93 2.091922724569846e-19

R81_94 V81 V94 -503.79671941533394
L81_94 V81 V94 -1.3275062373313003e-11
C81_94 V81 V94 -3.026491051827154e-20

R81_95 V81 V95 -2141.4695652126816
L81_95 V81 V95 4.489914153460516e-12
C81_95 V81 V95 1.905315940082879e-19

R81_96 V81 V96 -768.000246063349
L81_96 V81 V96 3.855230523709938e-12
C81_96 V81 V96 1.8609160421288978e-19

R81_97 V81 V97 717.8909814006148
L81_97 V81 V97 1.7398904953237619e-12
C81_97 V81 V97 3.4809619042696177e-19

R81_98 V81 V98 157.0911119886474
L81_98 V81 V98 -3.948402484987377e-11
C81_98 V81 V98 -2.1450776509710722e-20

R81_99 V81 V99 156.37149402211455
L81_99 V81 V99 3.360411038003538e-12
C81_99 V81 V99 -1.8580166842257116e-20

R81_100 V81 V100 178.59013175537484
L81_100 V81 V100 3.2327960139959422e-12
C81_100 V81 V100 1.9056949833585388e-20

R81_101 V81 V101 226.23921019236954
L81_101 V81 V101 -1.6584213207657825e-12
C81_101 V81 V101 -5.110500207270919e-19

R81_102 V81 V102 -3983.6478777513216
L81_102 V81 V102 2.9200120120753746e-12
C81_102 V81 V102 1.9888775622731979e-19

R81_103 V81 V103 -1919.8939213754923
L81_103 V81 V103 3.351194447259094e-11
C81_103 V81 V103 7.020290558018887e-20

R81_104 V81 V104 2110.443391763368
L81_104 V81 V104 -2.307334784302266e-11
C81_104 V81 V104 -4.0106001452509705e-20

R81_105 V81 V105 -95.23519270092042
L81_105 V81 V105 -2.8039094945588726e-12
C81_105 V81 V105 6.120659317565516e-21

R81_106 V81 V106 -963.1939722851178
L81_106 V81 V106 -6.507353657334868e-12
C81_106 V81 V106 -2.434183325523432e-19

R81_107 V81 V107 -370.90518978755586
L81_107 V81 V107 -3.899728289861446e-12
C81_107 V81 V107 -1.5007348080489304e-19

R81_108 V81 V108 -353.2887807732081
L81_108 V81 V108 -3.366191191694188e-12
C81_108 V81 V108 -1.2514687386323254e-19

R81_109 V81 V109 406.40434485674905
L81_109 V81 V109 -3.947769900589279e-12
C81_109 V81 V109 3.5291404754121135e-20

R81_110 V81 V110 -6978.2663366833685
L81_110 V81 V110 -6.4790505222757584e-12
C81_110 V81 V110 8.627854468385746e-21

R81_111 V81 V111 1748.170420921899
L81_111 V81 V111 -3.984619049032744e-12
C81_111 V81 V111 -1.1145901601050295e-19

R81_112 V81 V112 1473.2422532737228
L81_112 V81 V112 -9.176995494769157e-12
C81_112 V81 V112 -3.034410447701041e-20

R81_113 V81 V113 390.70125939244616
L81_113 V81 V113 2.993507588968712e-12
C81_113 V81 V113 3.145067562636144e-20

R81_114 V81 V114 2755.1571781242264
L81_114 V81 V114 5.2061488278471594e-12
C81_114 V81 V114 1.6860217108198668e-19

R81_115 V81 V115 466.14254344750833
L81_115 V81 V115 2.6054107817335947e-12
C81_115 V81 V115 2.654572644196492e-19

R81_116 V81 V116 383.08170718679247
L81_116 V81 V116 2.2065377875821453e-12
C81_116 V81 V116 2.485382387529714e-19

R81_117 V81 V117 -164.08107625184763
L81_117 V81 V117 4.294365394145851e-12
C81_117 V81 V117 2.9871792052267987e-19

R81_118 V81 V118 525.3531276229045
L81_118 V81 V118 1.000116399114077e-11
C81_118 V81 V118 -2.199679917752244e-20

R81_119 V81 V119 -6262.14623176143
L81_119 V81 V119 -9.454467773062311e-10
C81_119 V81 V119 -8.39323693670677e-20

R81_120 V81 V120 -1158.4088369791227
L81_120 V81 V120 -2.844872696332797e-11
C81_120 V81 V120 -6.865540103693715e-20

R81_121 V81 V121 830.5008650295379
L81_121 V81 V121 -2.4539895614034768e-11
C81_121 V81 V121 -2.7311226987508233e-19

R81_122 V81 V122 -1800.0935027500527
L81_122 V81 V122 -1.914851216631195e-11
C81_122 V81 V122 -7.995764555394799e-20

R81_123 V81 V123 -1075.1665390164576
L81_123 V81 V123 4.694818154248436e-11
C81_123 V81 V123 6.162752353817527e-20

R81_124 V81 V124 -997.6952256583514
L81_124 V81 V124 -5.376573847044157e-12
C81_124 V81 V124 -1.3302017503238371e-19

R81_125 V81 V125 -1151.9874503959327
L81_125 V81 V125 -9.632295598765903e-13
C81_125 V81 V125 -4.0297274799937224e-19

R81_126 V81 V126 -378.94844516780915
L81_126 V81 V126 -3.1109932871661382e-12
C81_126 V81 V126 -1.6619143251122035e-19

R81_127 V81 V127 -1278.8016728123055
L81_127 V81 V127 -6.026109636325741e-12
C81_127 V81 V127 -1.3160523867664073e-19

R81_128 V81 V128 -5808.283567346315
L81_128 V81 V128 -5.316530599406417e-12
C81_128 V81 V128 -7.421067641172204e-20

R81_129 V81 V129 -330.510258041247
L81_129 V81 V129 3.917177065487563e-12
C81_129 V81 V129 3.128772242961562e-19

R81_130 V81 V130 450.6989542685535
L81_130 V81 V130 2.4268854967709694e-12
C81_130 V81 V130 2.705379537058655e-19

R81_131 V81 V131 503.6306738482742
L81_131 V81 V131 1.3688823726664401e-11
C81_131 V81 V131 8.676904977328463e-20

R81_132 V81 V132 378.33067283735664
L81_132 V81 V132 2.736181078868913e-12
C81_132 V81 V132 2.397700058658004e-19

R81_133 V81 V133 385.3118120307275
L81_133 V81 V133 2.438691747927652e-12
C81_133 V81 V133 7.269569641492205e-20

R81_134 V81 V134 905.8023882389056
L81_134 V81 V134 1.0319011199892377e-11
C81_134 V81 V134 -1.1476302566175598e-19

R81_135 V81 V135 9777.664486002835
L81_135 V81 V135 5.168477259915807e-12
C81_135 V81 V135 1.3120443725720396e-19

R81_136 V81 V136 6503.094760677231
L81_136 V81 V136 1.0702821839811837e-11
C81_136 V81 V136 -3.895082692059113e-20

R81_137 V81 V137 -801.5938283286572
L81_137 V81 V137 3.9242872462956704e-12
C81_137 V81 V137 1.8402460650795738e-19

R81_138 V81 V138 -339.4390430214384
L81_138 V81 V138 -3.0215342458066147e-12
C81_138 V81 V138 -1.8399450370152383e-20

R81_139 V81 V139 -887.792819642913
L81_139 V81 V139 -3.744396330785706e-12
C81_139 V81 V139 -1.9768155985855257e-19

R81_140 V81 V140 -443.457847597444
L81_140 V81 V140 -1.6641425712270894e-11
C81_140 V81 V140 5.506802238046015e-20

R81_141 V81 V141 637.5684726198426
L81_141 V81 V141 -2.056016986066716e-12
C81_141 V81 V141 -3.675370111386769e-19

R81_142 V81 V142 558.7712352196713
L81_142 V81 V142 6.468823419904516e-11
C81_142 V81 V142 2.797592525868112e-20

R81_143 V81 V143 1346.8542574162445
L81_143 V81 V143 4.998465849223311e-12
C81_143 V81 V143 6.303444891731459e-20

R81_144 V81 V144 649.3548420807732
L81_144 V81 V144 -1.0971247510428847e-11
C81_144 V81 V144 -1.1261638942932563e-19

R81_145 V81 V145 -193.4724683999681
L81_145 V81 V145 -1.275584352312388e-12
C81_145 V81 V145 -2.5796012491818246e-19

R81_146 V81 V146 1353.255903335149
L81_146 V81 V146 5.411602191336173e-12
C81_146 V81 V146 6.55208554491501e-20

R81_147 V81 V147 39511.46732315795
L81_147 V81 V147 -4.966832373588242e-12
C81_147 V81 V147 -5.438283835349949e-20

R81_148 V81 V148 -695.3637033009041
L81_148 V81 V148 -3.188674973566928e-12
C81_148 V81 V148 -1.3787340560740795e-19

R81_149 V81 V149 180.343277446136
L81_149 V81 V149 1.7183806393420377e-12
C81_149 V81 V149 2.9057179604262154e-19

R81_150 V81 V150 2730.7618127338733
L81_150 V81 V150 -5.359819303489622e-12
C81_150 V81 V150 -2.1939361714617454e-19

R81_151 V81 V151 -1114.8306833693418
L81_151 V81 V151 -2.8937220795445992e-12
C81_151 V81 V151 -7.313877121827955e-20

R81_152 V81 V152 939.3644226923568
L81_152 V81 V152 8.021491768476213e-12
C81_152 V81 V152 7.233035717856762e-20

R81_153 V81 V153 -358.5986874182088
L81_153 V81 V153 1.4893858513397065e-12
C81_153 V81 V153 3.4608268373550815e-19

R81_154 V81 V154 2559.9206557733846
L81_154 V81 V154 6.997518775512333e-12
C81_154 V81 V154 1.6497001203808388e-19

R81_155 V81 V155 374.7917017714921
L81_155 V81 V155 4.668259303024908e-12
C81_155 V81 V155 -3.366018305876347e-20

R81_156 V81 V156 2009.464837774751
L81_156 V81 V156 5.841887767204083e-12
C81_156 V81 V156 1.4352332489619922e-19

R81_157 V81 V157 -516.3401289155265
L81_157 V81 V157 -2.224698688731827e-12
C81_157 V81 V157 -1.6624034042829184e-19

R81_158 V81 V158 12532.684194971418
L81_158 V81 V158 6.114683962507699e-11
C81_158 V81 V158 -2.8905042041474047e-20

R81_159 V81 V159 -2135.627713521275
L81_159 V81 V159 2.0070234122526936e-12
C81_159 V81 V159 2.4886183358756326e-19

R81_160 V81 V160 1326.2568747941982
L81_160 V81 V160 3.1061890028735414e-12
C81_160 V81 V160 6.920570368667765e-20

R81_161 V81 V161 -260.4608260899886
L81_161 V81 V161 -3.0581134981099664e-12
C81_161 V81 V161 -2.547052285239645e-19

R81_162 V81 V162 -1969.8352639862183
L81_162 V81 V162 7.950212991199928e-12
C81_162 V81 V162 1.6089522688162397e-19

R81_163 V81 V163 -6902.512358116429
L81_163 V81 V163 5.008676830499919e-12
C81_163 V81 V163 6.15407326383197e-20

R81_164 V81 V164 -412.75695690426267
L81_164 V81 V164 -1.0656711980343121e-11
C81_164 V81 V164 1.9217299866965276e-20

R81_165 V81 V165 -308.6679464738138
L81_165 V81 V165 -9.674225060880525e-13
C81_165 V81 V165 -1.950703786172775e-19

R81_166 V81 V166 347.4453504880119
L81_166 V81 V166 -3.6148290654790935e-12
C81_166 V81 V166 -1.6142217503704284e-19

R81_167 V81 V167 1610.6432007550711
L81_167 V81 V167 -1.8141705232621105e-12
C81_167 V81 V167 -2.2385504538660507e-19

R81_168 V81 V168 327.2147106464619
L81_168 V81 V168 -2.4195445787640816e-12
C81_168 V81 V168 -3.3729887171037997e-19

R81_169 V81 V169 459.6528927231614
L81_169 V81 V169 1.058908066447563e-12
C81_169 V81 V169 3.242389173930235e-19

R81_170 V81 V170 -497.8635647469157
L81_170 V81 V170 -3.5739943983887405e-12
C81_170 V81 V170 -6.55342145776418e-20

R81_171 V81 V171 -1455.7592071776971
L81_171 V81 V171 -5.039008836098537e-12
C81_171 V81 V171 -2.616162373140081e-20

R81_172 V81 V172 -9583.598596091353
L81_172 V81 V172 -2.7493529534818548e-11
C81_172 V81 V172 1.1645584465389485e-19

R81_173 V81 V173 -314.0064422959768
L81_173 V81 V173 5.373854569341199e-12
C81_173 V81 V173 1.8080392477346724e-19

R81_174 V81 V174 1302.4022765444813
L81_174 V81 V174 1.170921530144321e-12
C81_174 V81 V174 2.7684383919973707e-19

R81_175 V81 V175 916.6537321922567
L81_175 V81 V175 1.2630492771343889e-12
C81_175 V81 V175 2.4023092774212643e-19

R81_176 V81 V176 -4837.516018266573
L81_176 V81 V176 1.1657186217244076e-12
C81_176 V81 V176 3.611032063206595e-19

R81_177 V81 V177 -1601.5847443334844
L81_177 V81 V177 -7.124572603667898e-12
C81_177 V81 V177 -9.610518826166157e-20

R81_178 V81 V178 -666.166851724957
L81_178 V81 V178 1.0351695845555015e-10
C81_178 V81 V178 -2.2778790437861046e-20

R81_179 V81 V179 -12523.187864429116
L81_179 V81 V179 -3.755120787665471e-12
C81_179 V81 V179 -6.416617660350753e-20

R81_180 V81 V180 -699.1835872462971
L81_180 V81 V180 -3.006378677452443e-12
C81_180 V81 V180 -1.4511646945644986e-19

R81_181 V81 V181 400.8874799484606
L81_181 V81 V181 -1.3036690928509931e-12
C81_181 V81 V181 -6.048780154743223e-19

R81_182 V81 V182 484.30710343926955
L81_182 V81 V182 -2.8168955664584467e-12
C81_182 V81 V182 -5.648973425918879e-20

R81_183 V81 V183 -1890.5910680190714
L81_183 V81 V183 -6.502015805284347e-12
C81_183 V81 V183 -3.624259925632167e-20

R81_184 V81 V184 2629.524451759738
L81_184 V81 V184 -2.5749295858186875e-12
C81_184 V81 V184 -7.068714853513559e-20

R81_185 V81 V185 -300.40976682662114
L81_185 V81 V185 -8.473802394928285e-12
C81_185 V81 V185 3.9339106748539263e-19

R81_186 V81 V186 320.6441805941348
L81_186 V81 V186 -2.3108177595966837e-12
C81_186 V81 V186 -1.8791051627099766e-19

R81_187 V81 V187 2519.678344556551
L81_187 V81 V187 -1.0233808086324917e-11
C81_187 V81 V187 -1.4457800447977452e-20

R81_188 V81 V188 1000.3041670932165
L81_188 V81 V188 -1.874582477005421e-11
C81_188 V81 V188 -8.732225660001746e-20

R81_189 V81 V189 265.7653222692283
L81_189 V81 V189 7.689298503852419e-13
C81_189 V81 V189 2.640049779879223e-19

R81_190 V81 V190 -400.4055929698569
L81_190 V81 V190 3.5103739190064944e-12
C81_190 V81 V190 -1.9500994982028147e-21

R81_191 V81 V191 -470.07790991898656
L81_191 V81 V191 7.15173397094862e-12
C81_191 V81 V191 1.0238740969664677e-19

R81_192 V81 V192 -390.7188694661546
L81_192 V81 V192 2.3268494442656823e-12
C81_192 V81 V192 2.622692989360266e-19

R81_193 V81 V193 1587.3034937942211
L81_193 V81 V193 -2.628983223168934e-12
C81_193 V81 V193 -1.8475690792295675e-20

R81_194 V81 V194 -627.3477187732414
L81_194 V81 V194 1.1929394268793328e-12
C81_194 V81 V194 2.617541644465608e-19

R81_195 V81 V195 6135.479411436586
L81_195 V81 V195 -1.1142548030590902e-11
C81_195 V81 V195 -1.7060556537078343e-19

R81_196 V81 V196 -4006.9155590467008
L81_196 V81 V196 4.370482675757761e-12
C81_196 V81 V196 9.254957375372032e-21

R81_197 V81 V197 -293.3342573486776
L81_197 V81 V197 -2.0134596843490275e-12
C81_197 V81 V197 -2.543323677040695e-19

R81_198 V81 V198 262.4062929095285
L81_198 V81 V198 -2.827422587614735e-12
C81_198 V81 V198 -3.4837609758253946e-20

R81_199 V81 V199 247.49506754667075
L81_199 V81 V199 -7.328349439361516e-12
C81_199 V81 V199 7.71660160282941e-20

R81_200 V81 V200 284.66451585252804
L81_200 V81 V200 -1.8678511416397742e-12
C81_200 V81 V200 -1.7007896924233166e-19

R82_82 V82 0 270.24940777690574
L82_82 V82 0 4.686145924019353e-13
C82_82 V82 0 1.8239592624725553e-18

R82_83 V82 V83 -1403.7564053072197
L82_83 V82 V83 -3.6612346639404145e-11
C82_83 V82 V83 2.5403047837650028e-20

R82_84 V82 V84 -1467.7551567631936
L82_84 V82 V84 -3.700314602461857e-12
C82_84 V82 V84 -1.0340140429230059e-19

R82_85 V82 V85 -1908.447483263024
L82_85 V82 V85 3.988170372007555e-12
C82_85 V82 V85 1.8420640939948333e-19

R82_86 V82 V86 -314.8395206536781
L82_86 V82 V86 1.1661398824348195e-11
C82_86 V82 V86 1.3658726834482387e-19

R82_87 V82 V87 32447.81654755441
L82_87 V82 V87 5.535576140332844e-12
C82_87 V82 V87 1.4672777768747793e-19

R82_88 V82 V88 -2962.8040890495877
L82_88 V82 V88 2.7965987698825576e-12
C82_88 V82 V88 2.8539914409863917e-19

R82_89 V82 V89 -1291.1559239383785
L82_89 V82 V89 2.839180640021944e-12
C82_89 V82 V89 2.5101629179669807e-19

R82_90 V82 V90 207.19043889953696
L82_90 V82 V90 7.854346417389327e-13
C82_90 V82 V90 8.940151979291635e-19

R82_91 V82 V91 1276.663247079182
L82_91 V82 V91 -3.0433985406886864e-12
C82_91 V82 V91 -2.640969365134271e-19

R82_92 V82 V92 1827.0396974694686
L82_92 V82 V92 -7.783779923833282e-12
C82_92 V82 V92 -1.2110446549109269e-19

R82_93 V82 V93 611.4294351277643
L82_93 V82 V93 -3.5370579664402097e-12
C82_93 V82 V93 -2.223138794723113e-19

R82_94 V82 V94 -1130.2805635750672
L82_94 V82 V94 -1.6872358013296799e-12
C82_94 V82 V94 -5.503001868620753e-19

R82_95 V82 V95 -1529.895137840243
L82_95 V82 V95 -8.368280400164609e-12
C82_95 V82 V95 -1.2781092428057802e-19

R82_96 V82 V96 -2662.982608744123
L82_96 V82 V96 -6.235793332361845e-12
C82_96 V82 V96 -2.0184009926391276e-19

R82_97 V82 V97 -4380.423243360482
L82_97 V82 V97 -2.1760274933695974e-12
C82_97 V82 V97 -4.553833690256788e-19

R82_98 V82 V98 -393.9781150223703
L82_98 V82 V98 -1.7362355795052666e-12
C82_98 V82 V98 -4.257464370351291e-19

R82_99 V82 V99 5044.803575621007
L82_99 V82 V99 1.819088023468831e-12
C82_99 V82 V99 4.1421111969432285e-19

R82_100 V82 V100 3469.6233826716416
L82_100 V82 V100 8.152238236211733e-12
C82_100 V82 V100 2.3753928688335407e-19

R82_101 V82 V101 -2823.123948885112
L82_101 V82 V101 2.0389690230352425e-12
C82_101 V82 V101 3.894378786500942e-19

R82_102 V82 V102 326.7428269919711
L82_102 V82 V102 1.2219356114181207e-12
C82_102 V82 V102 5.979431831668371e-19

R82_103 V82 V103 -2291.2167660780765
L82_103 V82 V103 -1.4057520871999254e-11
C82_103 V82 V103 -1.833210789813445e-21

R82_104 V82 V104 -1586.8654619828674
L82_104 V82 V104 -1.3353526529965541e-11
C82_104 V82 V104 -2.4507060213047375e-20

R82_105 V82 V105 1864.0152253787587
L82_105 V82 V105 5.803034090061255e-12
C82_105 V82 V105 2.0351055149629494e-19

R82_106 V82 V106 -257.65034840305765
L82_106 V82 V106 2.353624188922913e-11
C82_106 V82 V106 4.7949382932610745e-20

R82_107 V82 V107 4421.70578640397
L82_107 V82 V107 -2.97037069816925e-12
C82_107 V82 V107 -2.951922518825697e-19

R82_108 V82 V108 -52919.53675388536
L82_108 V82 V108 4.9788948831537305e-12
C82_108 V82 V108 5.065170434997247e-20

R82_109 V82 V109 1271.5510675498772
L82_109 V82 V109 -2.7979735349368056e-12
C82_109 V82 V109 -4.1637575103853986e-19

R82_110 V82 V110 435.6280513964978
L82_110 V82 V110 -1.6490640207883866e-12
C82_110 V82 V110 -4.414021547663759e-19

R82_111 V82 V111 3882.4569181453326
L82_111 V82 V111 -6.865094229286561e-11
C82_111 V82 V111 2.131878106246126e-21

R82_112 V82 V112 2394.843163268854
L82_112 V82 V112 -6.9677001867562875e-12
C82_112 V82 V112 -1.1737711694825001e-19

R82_113 V82 V113 1077.4118003724982
L82_113 V82 V113 -6.407960072434053e-12
C82_113 V82 V113 -1.9981530729317966e-19

R82_114 V82 V114 323.6433624059741
L82_114 V82 V114 6.785848823381978e-12
C82_114 V82 V114 4.723366918197508e-21

R82_115 V82 V115 -2613.1640877317363
L82_115 V82 V115 2.434344892167857e-12
C82_115 V82 V115 2.4020913560876526e-19

R82_116 V82 V116 -5393.360112791548
L82_116 V82 V116 4.5669583429754256e-11
C82_116 V82 V116 -2.6574440517478006e-20

R82_117 V82 V117 -675.7828576714046
L82_117 V82 V117 4.58562832527124e-12
C82_117 V82 V117 2.9532926047178715e-19

R82_118 V82 V118 -127.64417503870746
L82_118 V82 V118 1.898073474035169e-12
C82_118 V82 V118 5.309235262600335e-19

R82_119 V82 V119 -1270.4346048637783
L82_119 V82 V119 2.1123685668638574e-11
C82_119 V82 V119 6.868765784732571e-20

R82_120 V82 V120 -3024.4888055741158
L82_120 V82 V120 3.1509166691958935e-12
C82_120 V82 V120 2.867855530296732e-19

R82_121 V82 V121 2058.5203125416174
L82_121 V82 V121 4.050478569494928e-12
C82_121 V82 V121 1.0184148083149027e-19

R82_122 V82 V122 389.366420157335
L82_122 V82 V122 -3.0712489160692016e-12
C82_122 V82 V122 -4.030961751140622e-19

R82_123 V82 V123 6813.233609314386
L82_123 V82 V123 -3.3821805855860006e-12
C82_123 V82 V123 -1.7485664531388694e-19

R82_124 V82 V124 -70953.43940049381
L82_124 V82 V124 -2.722902753633413e-12
C82_124 V82 V124 -2.9172094488434093e-19

R82_125 V82 V125 633.319328005829
L82_125 V82 V125 -6.296901039714214e-12
C82_125 V82 V125 -1.1731810654373537e-19

R82_126 V82 V126 143.79396284234906
L82_126 V82 V126 -2.9056488794958813e-12
C82_126 V82 V126 -1.8855553947558988e-19

R82_127 V82 V127 483.2622760783721
L82_127 V82 V127 -1.723338833517711e-11
C82_127 V82 V127 -7.508415368685316e-20

R82_128 V82 V128 613.2097276323108
L82_128 V82 V128 -1.5215741808014018e-11
C82_128 V82 V128 -8.51133223356964e-20

R82_129 V82 V129 -2364.4886888835995
L82_129 V82 V129 -2.5847682402723935e-12
C82_129 V82 V129 -3.6400006953307334e-19

R82_130 V82 V130 -169.27816987209647
L82_130 V82 V130 1.6065173085431112e-12
C82_130 V82 V130 4.443934825695849e-19

R82_131 V82 V131 -357.04821177752217
L82_131 V82 V131 6.075479662081016e-12
C82_131 V82 V131 1.3783812260646185e-19

R82_132 V82 V132 -288.7105634790771
L82_132 V82 V132 2.7108225228309016e-12
C82_132 V82 V132 2.902317138673273e-19

R82_133 V82 V133 -783.3330597191479
L82_133 V82 V133 2.6521908713832262e-12
C82_133 V82 V133 3.5197771842774736e-19

R82_134 V82 V134 -686.9788068865469
L82_134 V82 V134 -2.053846650831716e-12
C82_134 V82 V134 -3.857228230100407e-19

R82_135 V82 V135 -2296.268008504969
L82_135 V82 V135 1.5102469856194724e-11
C82_135 V82 V135 -2.3138997887961908e-20

R82_136 V82 V136 -652.9800115974055
L82_136 V82 V136 -1.0786473923874328e-11
C82_136 V82 V136 -2.341397607376592e-19

R82_137 V82 V137 563.0425253873291
L82_137 V82 V137 3.1527047789379246e-12
C82_137 V82 V137 2.309315696996347e-19

R82_138 V82 V138 210.0261530501151
L82_138 V82 V138 -2.7652326798058467e-11
C82_138 V82 V138 8.611431794237761e-20

R82_139 V82 V139 305.34617124650185
L82_139 V82 V139 4.245401347695166e-12
C82_139 V82 V139 1.886578067603307e-19

R82_140 V82 V140 163.38248293103334
L82_140 V82 V140 7.1714496593160484e-12
C82_140 V82 V140 2.842954332574499e-19

R82_141 V82 V141 -698.336793552598
L82_141 V82 V141 -1.6132858999557912e-12
C82_141 V82 V141 -5.864675644515595e-19

R82_142 V82 V142 -2253.4332682832696
L82_142 V82 V142 6.326367533319613e-12
C82_142 V82 V142 8.671367198462077e-20

R82_143 V82 V143 -364.6333530346664
L82_143 V82 V143 -2.010639372600761e-12
C82_143 V82 V143 -2.6316945237665487e-19

R82_144 V82 V144 -273.12433174127085
L82_144 V82 V144 -4.501073632902086e-12
C82_144 V82 V144 -1.3786313005057197e-19

R82_145 V82 V145 -687.2296637453477
L82_145 V82 V145 -2.285335391478065e-12
C82_145 V82 V145 -2.2619732287404973e-19

R82_146 V82 V146 -163.4328297991341
L82_146 V82 V146 2.0466997020678387e-11
C82_146 V82 V146 5.202708239730322e-20

R82_147 V82 V147 -931.672457439988
L82_147 V82 V147 -8.891797306131735e-12
C82_147 V82 V147 -1.5613936155387773e-19

R82_148 V82 V148 -2590.3944258919314
L82_148 V82 V148 -2.9916726652961268e-12
C82_148 V82 V148 -1.9327760695066364e-19

R82_149 V82 V149 824.6820914601132
L82_149 V82 V149 7.271710495613861e-13
C82_149 V82 V149 9.573365618649148e-19

R82_150 V82 V150 3501.8478167588773
L82_150 V82 V150 1.2281629401185218e-11
C82_150 V82 V150 -5.02736922806552e-19

R82_151 V82 V151 309.4536511056064
L82_151 V82 V151 3.1312952174165163e-12
C82_151 V82 V151 2.2199301768699335e-19

R82_152 V82 V152 348.50408721984536
L82_152 V82 V152 4.446593131756448e-12
C82_152 V82 V152 5.108120919023155e-20

R82_153 V82 V153 388.40533233800005
L82_153 V82 V153 3.936548406693324e-12
C82_153 V82 V153 4.752025935487827e-20

R82_154 V82 V154 166.11243083392716
L82_154 V82 V154 -5.160028980853309e-12
C82_154 V82 V154 3.252487470164288e-19

R82_155 V82 V155 -820.1071055563515
L82_155 V82 V155 1.922063724267933e-12
C82_155 V82 V155 2.1617943858343163e-19

R82_156 V82 V156 -2981.204537429141
L82_156 V82 V156 4.754376345510474e-12
C82_156 V82 V156 2.1196087161653741e-19

R82_157 V82 V157 -1942.4667692066323
L82_157 V82 V157 -7.150708163602636e-13
C82_157 V82 V157 -9.320619071958766e-19

R82_158 V82 V158 -230.86058161565586
L82_158 V82 V158 -1.6992965789950922e-11
C82_158 V82 V158 6.384397008427504e-21

R82_159 V82 V159 -424.5048312202171
L82_159 V82 V159 -3.0686067105109007e-12
C82_159 V82 V159 -4.6462304989547735e-20

R82_160 V82 V160 -257.07258707907107
L82_160 V82 V160 -1.3061188418482227e-11
C82_160 V82 V160 2.0823647945763938e-20

R82_161 V82 V161 626.1985566654628
L82_161 V82 V161 5.261462237094784e-11
C82_161 V82 V161 4.3459099840965795e-20

R82_162 V82 V162 -698.452097002453
L82_162 V82 V162 1.18521008606624e-12
C82_162 V82 V162 1.132307990363217e-19

R82_163 V82 V163 428.66142877899097
L82_163 V82 V163 -2.8736605271118175e-12
C82_163 V82 V163 -1.7621926297415176e-19

R82_164 V82 V164 237.9334842463681
L82_164 V82 V164 -3.4620902484837076e-12
C82_164 V82 V164 1.3312108446133239e-20

R82_165 V82 V165 -1387.673540329754
L82_165 V82 V165 1.4036626114051229e-12
C82_165 V82 V165 4.436461239227078e-19

R82_166 V82 V166 223.42170783290626
L82_166 V82 V166 -4.608500912596891e-12
C82_166 V82 V166 -1.2977392597064821e-19

R82_167 V82 V167 6109.159303796905
L82_167 V82 V167 4.9154000029993705e-12
C82_167 V82 V167 3.733751349121671e-21

R82_168 V82 V168 -685.7540143342358
L82_168 V82 V168 3.0835239905188947e-12
C82_168 V82 V168 -1.3637549837123206e-19

R82_169 V82 V169 -411.83960200064496
L82_169 V82 V169 -8.713977639973324e-11
C82_169 V82 V169 -1.3294252704102676e-19

R82_170 V82 V170 -272.0274783179902
L82_170 V82 V170 -2.0888292170131342e-12
C82_170 V82 V170 2.612522967919635e-19

R82_171 V82 V171 -416.25925928210313
L82_171 V82 V171 2.0439643951224982e-12
C82_171 V82 V171 3.4294144708314435e-19

R82_172 V82 V172 -482.2058523341271
L82_172 V82 V172 1.7245770625578728e-11
C82_172 V82 V172 2.0338379802536361e-19

R82_173 V82 V173 375.4276294708416
L82_173 V82 V173 -1.926635905246226e-12
C82_173 V82 V173 -1.232858517125169e-19

R82_174 V82 V174 -369.79076896557433
L82_174 V82 V174 1.9247654923325373e-12
C82_174 V82 V174 -2.502330361038779e-19

R82_175 V82 V175 1447.3139815019194
L82_175 V82 V175 -1.4178181510252027e-10
C82_175 V82 V175 7.550410427036832e-20

R82_176 V82 V176 485.72768541251247
L82_176 V82 V176 -8.450344423344193e-12
C82_176 V82 V176 1.2047646655945805e-19

R82_177 V82 V177 1030.9925508233916
L82_177 V82 V177 -3.028278258966783e-11
C82_177 V82 V177 1.1113425038614904e-19

R82_178 V82 V178 212.70232996936926
L82_178 V82 V178 6.251149445221846e-11
C82_178 V82 V178 -1.8808215406442596e-19

R82_179 V82 V179 2904.5238507101217
L82_179 V82 V179 -1.6349779813813052e-12
C82_179 V82 V179 -4.420671105199719e-19

R82_180 V82 V180 2628.301157183792
L82_180 V82 V180 -2.3820157824496427e-12
C82_180 V82 V180 -3.561217257576108e-19

R82_181 V82 V181 -432.1949759472853
L82_181 V82 V181 -4.089804254032312e-11
C82_181 V82 V181 -1.0205117355448878e-19

R82_182 V82 V182 -350.11653855699996
L82_182 V82 V182 5.662279461683607e-12
C82_182 V82 V182 2.8831180376551727e-19

R82_183 V82 V183 -232771.08695799866
L82_183 V82 V183 -2.7465618419015494e-12
C82_183 V82 V183 -7.192391360256344e-20

R82_184 V82 V184 -1612.5240810607377
L82_184 V82 V184 -6.801027389899698e-12
C82_184 V82 V184 3.1774730199260426e-20

R82_185 V82 V185 1162.6983782558823
L82_185 V82 V185 5.0330124789919276e-12
C82_185 V82 V185 -4.4950791971724467e-23

R82_186 V82 V186 -375.55800738165095
L82_186 V82 V186 3.4708996310911463e-11
C82_186 V82 V186 2.064784611291194e-20

R82_187 V82 V187 14076.04906196547
L82_187 V82 V187 1.4412850730244392e-12
C82_187 V82 V187 3.5649374402813763e-19

R82_188 V82 V188 1710.7749306831374
L82_188 V82 V188 1.3581725633535362e-12
C82_188 V82 V188 2.685004049612257e-19

R82_189 V82 V189 1787.5601536462325
L82_189 V82 V189 3.6530431112025496e-12
C82_189 V82 V189 2.2607873781359533e-19

R82_190 V82 V190 630.1515460634785
L82_190 V82 V190 8.537960871765188e-12
C82_190 V82 V190 -2.9036195569206675e-19

R82_191 V82 V191 1594.4491173918811
L82_191 V82 V191 1.5698565929746274e-12
C82_191 V82 V191 1.889837438127363e-19

R82_192 V82 V192 1159.2768396272356
L82_192 V82 V192 7.400785418348327e-12
C82_192 V82 V192 6.415952366003759e-20

R82_193 V82 V193 -3058.178518206732
L82_193 V82 V193 -1.930984007519228e-12
C82_193 V82 V193 -1.795184128451238e-19

R82_194 V82 V194 -1309.7268981785953
L82_194 V82 V194 -2.0873189356716644e-11
C82_194 V82 V194 -1.1750977473363719e-19

R82_195 V82 V195 -3131.6612208075326
L82_195 V82 V195 -1.0621283301531067e-12
C82_195 V82 V195 -4.334508732036681e-19

R82_196 V82 V196 -11419.61164578982
L82_196 V82 V196 -1.3972061257991086e-12
C82_196 V82 V196 -2.7278368003787203e-19

R82_197 V82 V197 5923.910555287273
L82_197 V82 V197 -2.8664481032463425e-12
C82_197 V82 V197 -1.288209324044045e-19

R82_198 V82 V198 -932.6056465688713
L82_198 V82 V198 -4.0949777012938396e-12
C82_198 V82 V198 4.91110638631676e-20

R82_199 V82 V199 -1695.004762074211
L82_199 V82 V199 -2.035124090071489e-12
C82_199 V82 V199 -1.6836573502013345e-19

R82_200 V82 V200 -1933.6771836749945
L82_200 V82 V200 -3.6070014122760577e-12
C82_200 V82 V200 -3.4290352526785064e-20

R83_83 V83 0 -8384.444441763504
L83_83 V83 0 -6.561103909802085e-12
C83_83 V83 0 1.2884723411162958e-19

R83_84 V83 V84 -1068.9810278085408
L83_84 V83 V84 -3.38571208382203e-12
C83_84 V83 V84 -1.215720911341962e-19

R83_85 V83 V85 -1448.2925467068603
L83_85 V83 V85 2.406954795130448e-11
C83_85 V83 V85 1.506056755843996e-20

R83_86 V83 V86 -403.68748609213645
L83_86 V83 V86 -6.8534883790983915e-12
C83_86 V83 V86 -6.210676874669725e-20

R83_87 V83 V87 -673.5229192723473
L83_87 V83 V87 1.2288064025496799e-12
C83_87 V83 V87 4.747675354178601e-19

R83_88 V83 V88 -1299.375541240937
L83_88 V83 V88 8.284801734303858e-12
C83_88 V83 V88 1.2755604250016145e-19

R83_89 V83 V89 -584.3025849587177
L83_89 V83 V89 2.237684345219742e-11
C83_89 V83 V89 6.160949713076338e-20

R83_90 V83 V90 451.31725836164253
L83_90 V83 V90 7.379008951836998e-12
C83_90 V83 V90 1.5370534800104988e-20

R83_91 V83 V91 328.4401382535978
L83_91 V83 V91 -3.1941267819528598e-12
C83_91 V83 V91 -5.618460627861653e-20

R83_92 V83 V92 1066.7430922749757
L83_92 V83 V92 3.4111082855691056e-11
C83_92 V83 V92 -8.688279371364365e-20

R83_93 V83 V93 379.86229624837983
L83_93 V83 V93 -2.137496744566366e-11
C83_93 V83 V93 -3.605841523646436e-20

R83_94 V83 V94 1311.5119530830798
L83_94 V83 V94 5.406977647300194e-12
C83_94 V83 V94 1.0203698126101649e-19

R83_95 V83 V95 1717.635502971916
L83_95 V83 V95 -2.3655358456230663e-12
C83_95 V83 V95 -3.389621332437505e-19

R83_96 V83 V96 1416.9146805153953
L83_96 V83 V96 -3.1662744974197657e-11
C83_96 V83 V96 -1.1228088677371246e-20

R83_97 V83 V97 9743.449949839713
L83_97 V83 V97 -6.464037649121334e-12
C83_97 V83 V97 -1.659535063800501e-19

R83_98 V83 V98 -414.09184726785014
L83_98 V83 V98 -3.961834051187329e-12
C83_98 V83 V98 -1.2678241902936562e-19

R83_99 V83 V99 -272.46309786136845
L83_99 V83 V99 1.4038522790142393e-12
C83_99 V83 V99 2.8312455341289452e-19

R83_100 V83 V100 -774.3309451110049
L83_100 V83 V100 3.6836965049022715e-11
C83_100 V83 V100 9.81545412425543e-20

R83_101 V83 V101 -678.4603691393435
L83_101 V83 V101 4.3285077024806904e-12
C83_101 V83 V101 1.7735458324289586e-19

R83_102 V83 V102 2715.97580967299
L83_102 V83 V102 -7.422276235595321e-12
C83_102 V83 V102 -1.1642931220087588e-19

R83_103 V83 V103 834.3144955100671
L83_103 V83 V103 -5.127217996816262e-12
C83_103 V83 V103 6.020458223157905e-20

R83_104 V83 V104 -2138.747915554296
L83_104 V83 V104 -8.733970300145011e-12
C83_104 V83 V104 -9.68492865424122e-20

R83_105 V83 V105 448.8342096802935
L83_105 V83 V105 -2.3924514477251094e-11
C83_105 V83 V105 -3.0280455298468424e-20

R83_106 V83 V106 -8539.658503670204
L83_106 V83 V106 2.1922689179206774e-12
C83_106 V83 V106 2.642874054879628e-19

R83_107 V83 V107 876.1768860176346
L83_107 V83 V107 -2.82278704839603e-12
C83_107 V83 V107 -1.8157490878619923e-19

R83_108 V83 V108 1806.79929279153
L83_108 V83 V108 9.33725119909691e-12
C83_108 V83 V108 5.228756023582503e-20

R83_109 V83 V109 23097.446025402187
L83_109 V83 V109 -5.809710800533026e-12
C83_109 V83 V109 -1.5340187070138155e-19

R83_110 V83 V110 10139.283259702413
L83_110 V83 V110 -9.859978749977018e-12
C83_110 V83 V110 -9.94955798048507e-21

R83_111 V83 V111 -628.2353663363358
L83_111 V83 V111 1.0789079850556137e-10
C83_111 V83 V111 -8.690469790546892e-20

R83_112 V83 V112 -2763.665947574233
L83_112 V83 V112 1.1427990858570108e-11
C83_112 V83 V112 6.759952632598834e-21

R83_113 V83 V113 16958.946170294545
L83_113 V83 V113 6.731545691828489e-12
C83_113 V83 V113 1.203481387957162e-19

R83_114 V83 V114 1789.5390313961084
L83_114 V83 V114 -3.202369889278205e-12
C83_114 V83 V114 -2.0922437197355606e-19

R83_115 V83 V115 4317.016644262469
L83_115 V83 V115 2.0340189502679282e-12
C83_115 V83 V115 1.67467162828631e-19

R83_116 V83 V116 -76495.08368814117
L83_116 V83 V116 -8.058388700541443e-12
C83_116 V83 V116 -7.176311972939543e-20

R83_117 V83 V117 1804.7691527936577
L83_117 V83 V117 -5.2608474805356716e-11
C83_117 V83 V117 -7.634426641200648e-21

R83_118 V83 V118 -663.9409540667143
L83_118 V83 V118 3.5129932392663943e-10
C83_118 V83 V118 -1.2122266735969948e-20

R83_119 V83 V119 -1365.6586321449427
L83_119 V83 V119 -2.218755891968073e-12
C83_119 V83 V119 3.745795925193226e-20

R83_120 V83 V120 -4637.398123131522
L83_120 V83 V120 4.385018439888982e-11
C83_120 V83 V120 6.97731912163341e-20

R83_121 V83 V121 7279.55623504484
L83_121 V83 V121 -4.6249787887429484e-11
C83_121 V83 V121 -4.4119847137061033e-20

R83_122 V83 V122 3186.2791009218486
L83_122 V83 V122 3.702177394451543e-12
C83_122 V83 V122 1.9193833524585623e-19

R83_123 V83 V123 3851.545121149036
L83_123 V83 V123 -5.2375057860611544e-12
C83_123 V83 V123 -2.5552380532881703e-19

R83_124 V83 V124 -39614.666668699865
L83_124 V83 V124 9.808012212279825e-12
C83_124 V83 V124 -3.494579060245163e-20

R83_125 V83 V125 1363.3959700577484
L83_125 V83 V125 -5.3552372011522236e-11
C83_125 V83 V125 1.0165690355263661e-20

R83_126 V83 V126 757.4514200312462
L83_126 V83 V126 1.468212486449426e-11
C83_126 V83 V126 4.937916904615901e-20

R83_127 V83 V127 518.828302303733
L83_127 V83 V127 1.7622099341723429e-12
C83_127 V83 V127 3.761640061697101e-20

R83_128 V83 V128 2755.5623644578222
L83_128 V83 V128 -6.690348755902797e-11
C83_128 V83 V128 4.085328008100622e-21

R83_129 V83 V129 2150.5706087863655
L83_129 V83 V129 5.064129033256912e-12
C83_129 V83 V129 6.349268569709092e-20

R83_130 V83 V130 -985.4807274723839
L83_130 V83 V130 -3.47567009037317e-12
C83_130 V83 V130 -1.9059834333738904e-19

R83_131 V83 V131 -350.879648282454
L83_131 V83 V131 -6.552270392615444e-12
C83_131 V83 V131 2.3780624767329225e-19

R83_132 V83 V132 -731.2826467249791
L83_132 V83 V132 -1.1074581556030994e-11
C83_132 V83 V132 5.602997393957141e-20

R83_133 V83 V133 -1007.9592383777397
L83_133 V83 V133 -4.404092735190615e-12
C83_133 V83 V133 -8.100710738379173e-20

R83_134 V83 V134 -54236.92723326813
L83_134 V83 V134 1.865529640645307e-10
C83_134 V83 V134 1.7118854966510529e-19

R83_135 V83 V135 7833.93829494844
L83_135 V83 V135 -3.2947664422540773e-12
C83_135 V83 V135 -2.358076369941154e-19

R83_136 V83 V136 7074.439154716785
L83_136 V83 V136 -3.5873354683080986e-11
C83_136 V83 V136 -1.0975818680158335e-19

R83_137 V83 V137 715.0975228912976
L83_137 V83 V137 -5.8067094226743745e-12
C83_137 V83 V137 -7.366455693396068e-20

R83_138 V83 V138 763.6923794850965
L83_138 V83 V138 6.392747382955891e-12
C83_138 V83 V138 -4.94195576365745e-20

R83_139 V83 V139 431.44760042919177
L83_139 V83 V139 6.2106146263440116e-12
C83_139 V83 V139 1.0485183942042634e-19

R83_140 V83 V140 601.0396100151651
L83_140 V83 V140 4.784191969714961e-12
C83_140 V83 V140 1.6520184125333127e-19

R83_141 V83 V141 -1019.3218073812599
L83_141 V83 V141 3.856682643517011e-12
C83_141 V83 V141 1.059179764692647e-19

R83_142 V83 V142 -740.3439899977279
L83_142 V83 V142 1.8810914179648286e-11
C83_142 V83 V142 -7.499568588188609e-20

R83_143 V83 V143 -387.1699511595229
L83_143 V83 V143 -1.8443107928040005e-11
C83_143 V83 V143 3.708566554339728e-20

R83_144 V83 V144 -559.2409841546346
L83_144 V83 V144 -6.155721967332295e-12
C83_144 V83 V144 -1.4965044820720992e-20

R83_145 V83 V145 -8485.976703165123
L83_145 V83 V145 1.3840810720641365e-11
C83_145 V83 V145 4.345841211132441e-20

R83_146 V83 V146 -596.835177820847
L83_146 V83 V146 -6.3765641560802254e-12
C83_146 V83 V146 5.584344565573745e-20

R83_147 V83 V147 1716.9406918608504
L83_147 V83 V147 2.9808154427185125e-12
C83_147 V83 V147 -8.762215749786075e-20

R83_148 V83 V148 6849.759471876493
L83_148 V83 V148 2.453853051847581e-11
C83_148 V83 V148 -1.0343468878093405e-19

R83_149 V83 V149 -2575.5367284681806
L83_149 V83 V149 -9.176797034189462e-12
C83_149 V83 V149 -1.106049025777142e-19

R83_150 V83 V150 733.5885347055281
L83_150 V83 V150 -5.920511958434937e-12
C83_150 V83 V150 6.94264113726434e-20

R83_151 V83 V151 727.2769643828651
L83_151 V83 V151 -2.978500991320447e-11
C83_151 V83 V151 -4.045918249932877e-20

R83_152 V83 V152 962.5132926965209
L83_152 V83 V152 5.9606934043513635e-12
C83_152 V83 V152 3.257538754075582e-20

R83_153 V83 V153 373.9306617553947
L83_153 V83 V153 -9.3395630099356e-12
C83_153 V83 V153 -5.792002720472392e-20

R83_154 V83 V154 674.0793147011308
L83_154 V83 V154 6.194989335909642e-12
C83_154 V83 V154 -1.2013063772097814e-19

R83_155 V83 V155 2169.1658026550176
L83_155 V83 V155 -6.407774709797631e-12
C83_155 V83 V155 1.8406490932400193e-19

R83_156 V83 V156 -1904.3429151135474
L83_156 V83 V156 1.741387679594506e-11
C83_156 V83 V156 3.7352223141946895e-20

R83_157 V83 V157 -5826.937111158184
L83_157 V83 V157 -1.012236072417899e-11
C83_157 V83 V157 4.9150063357719786e-20

R83_158 V83 V158 -481.8459946397486
L83_158 V83 V158 1.9552226597533208e-11
C83_158 V83 V158 5.71298979799808e-20

R83_159 V83 V159 -391.68615763295253
L83_159 V83 V159 -8.230929327222002e-12
C83_159 V83 V159 -1.8243691495114125e-19

R83_160 V83 V160 -712.103857765336
L83_160 V83 V160 -2.228786760405233e-12
C83_160 V83 V160 -5.583620719103552e-20

R83_161 V83 V161 1086.7431415658098
L83_161 V83 V161 2.9287717654779605e-12
C83_161 V83 V161 1.2866848117422898e-19

R83_162 V83 V162 -3979.448325470571
L83_162 V83 V162 -2.2087472953707512e-11
C83_162 V83 V162 -5.068331742354874e-21

R83_163 V83 V163 633.2057104065295
L83_163 V83 V163 1.0598538468828484e-12
C83_163 V83 V163 1.2918662594937117e-19

R83_164 V83 V164 818.438383513336
L83_164 V83 V164 2.7041649976994166e-12
C83_164 V83 V164 5.868275073204105e-20

R83_165 V83 V165 1210.8887448325572
L83_165 V83 V165 1.8702227415946044e-10
C83_165 V83 V165 -1.2002561758375003e-19

R83_166 V83 V166 574.7816918821159
L83_166 V83 V166 6.994509023195332e-12
C83_166 V83 V166 -4.57749694656343e-20

R83_167 V83 V167 -2104.9792599109146
L83_167 V83 V167 -9.838720068146595e-13
C83_167 V83 V167 -2.2764418579456478e-20

R83_168 V83 V168 -4303.527531938497
L83_168 V83 V168 2.635959398620281e-12
C83_168 V83 V168 7.693106324258335e-20

R83_169 V83 V169 -1436.2271566272398
L83_169 V83 V169 -1.079691420990393e-11
C83_169 V83 V169 -5.0115517618420234e-20

R83_170 V83 V170 -655.715280230293
L83_170 V83 V170 1.3211363450853276e-11
C83_170 V83 V170 9.916701483817466e-21

R83_171 V83 V171 -1268.975439261654
L83_171 V83 V171 -8.604746869308056e-12
C83_171 V83 V171 -1.4139107704391596e-20

R83_172 V83 V172 -978.8983358319493
L83_172 V83 V172 -3.055084643056141e-12
C83_172 V83 V172 -5.652065748455192e-20

R83_173 V83 V173 1386.514602529921
L83_173 V83 V173 -3.902305647705146e-11
C83_173 V83 V173 2.464091809771436e-21

R83_174 V83 V174 -919.3943288815819
L83_174 V83 V174 -3.545061706102231e-12
C83_174 V83 V174 -7.989707287513974e-21

R83_175 V83 V175 1828.5824373960481
L83_175 V83 V175 1.03507591391194e-12
C83_175 V83 V175 2.4540256615765312e-20

R83_176 V83 V176 1213.416451751492
L83_176 V83 V176 -2.961395640083864e-11
C83_176 V83 V176 -1.074770422501285e-20

R83_177 V83 V177 4534.037298208234
L83_177 V83 V177 -4.980393003332872e-12
C83_177 V83 V177 -3.285564176321582e-20

R83_178 V83 V178 513.9675246991906
L83_178 V83 V178 -2.4864342010154325e-11
C83_178 V83 V178 3.1892849223891867e-20

R83_179 V83 V179 1106.9867002296482
L83_179 V83 V179 -3.818771988238095e-12
C83_179 V83 V179 -1.4804422993172555e-20

R83_180 V83 V180 1881.2530136881517
L83_180 V83 V180 1.8669469351350086e-11
C83_180 V83 V180 4.935007758388124e-21

R83_181 V83 V181 -956.3837015211959
L83_181 V83 V181 2.0182582892650646e-11
C83_181 V83 V181 9.983362598217473e-20

R83_182 V83 V182 -1635.6088856559054
L83_182 V83 V182 1.2618202758090538e-11
C83_182 V83 V182 -2.916901146888583e-20

R83_183 V83 V183 -673.6849766524311
L83_183 V83 V183 -1.656959479551106e-12
C83_183 V83 V183 1.793510128560292e-20

R83_184 V83 V184 -946.1542110528968
L83_184 V83 V184 -8.636000390895495e-12
C83_184 V83 V184 4.090168945746949e-20

R83_185 V83 V185 899.0929954866447
L83_185 V83 V185 2.8956019527796615e-12
C83_185 V83 V185 -3.1350775992012866e-20

R83_186 V83 V186 -600.3102047254273
L83_186 V83 V186 7.988933881654493e-12
C83_186 V83 V186 1.319077911719736e-20

R83_187 V83 V187 2453.7540091841706
L83_187 V83 V187 1.7579976233854259e-12
C83_187 V83 V187 7.735040879898641e-20

R83_188 V83 V188 825.9215718243264
L83_188 V83 V188 4.136602672389628e-12
C83_188 V83 V188 4.805164735591984e-21

R83_189 V83 V189 -1549.672044298918
L83_189 V83 V189 -5.867778808594687e-12
C83_189 V83 V189 -1.0570647604729591e-19

R83_190 V83 V190 1185.5341894454164
L83_190 V83 V190 -5.878237742346563e-12
C83_190 V83 V190 1.9619157144189727e-20

R83_191 V83 V191 493.5298808706037
L83_191 V83 V191 3.0990132793430573e-12
C83_191 V83 V191 -1.6994752053644443e-19

R83_192 V83 V192 909.8433248184651
L83_192 V83 V192 1.1468492423257809e-11
C83_192 V83 V192 -1.4091445825439408e-19

R83_193 V83 V193 -2681.9110037290843
L83_193 V83 V193 -3.177549731350487e-12
C83_193 V83 V193 1.5278530826255355e-20

R83_194 V83 V194 1847.270698445255
L83_194 V83 V194 1.9334512935004284e-11
C83_194 V83 V194 -4.7934730364246147e-20

R83_195 V83 V195 -632.3400851814334
L83_195 V83 V195 -2.8632307438463584e-12
C83_195 V83 V195 1.6249784406279678e-19

R83_196 V83 V196 -925.7381324457482
L83_196 V83 V196 -3.7486358830726035e-12
C83_196 V83 V196 1.1085188500624902e-19

R83_197 V83 V197 1735.781375125543
L83_197 V83 V197 5.174891017400548e-12
C83_197 V83 V197 1.1947535180679892e-19

R83_198 V83 V198 -839.0139268041693
L83_198 V83 V198 1.9589666596101787e-11
C83_198 V83 V198 -5.267625412824943e-20

R83_199 V83 V199 -652.2256682238882
L83_199 V83 V199 -5.758741917246405e-12
C83_199 V83 V199 9.643924723822419e-20

R83_200 V83 V200 -1039.3250664314035
L83_200 V83 V200 -2.6543490149314147e-11
C83_200 V83 V200 1.0220441579296364e-19

R84_84 V84 0 1391.017205619349
L84_84 V84 0 2.571891041751061e-13
C84_84 V84 0 1.6593862564854512e-18

R84_85 V84 V85 -1912.9793483672574
L84_85 V84 V85 -4.0554514221034576e-11
C84_85 V84 V85 -9.882631069041538e-21

R84_86 V84 V86 -515.8188898683787
L84_86 V84 V86 -8.10139998263631e-12
C84_86 V84 V86 -1.9077218875611686e-20

R84_87 V84 V87 -2177.4957729744597
L84_87 V84 V87 3.166573327133828e-12
C84_87 V84 V87 1.572040836931563e-19

R84_88 V84 V88 -702.0440274086803
L84_88 V84 V88 8.096807166045148e-13
C84_88 V84 V88 6.032696623036382e-19

R84_89 V84 V89 -796.4965863854003
L84_89 V84 V89 2.6889029031358018e-12
C84_89 V84 V89 1.6879396595142976e-19

R84_90 V84 V90 533.5642991668927
L84_90 V84 V90 1.3354030849641196e-12
C84_90 V84 V90 2.422247377856558e-19

R84_91 V84 V91 1183.4527264581398
L84_91 V84 V91 -2.127102545357248e-12
C84_91 V84 V91 -1.9734826957456353e-19

R84_92 V84 V92 406.00915803631983
L84_92 V84 V92 -2.3281895864949188e-12
C84_92 V84 V92 -1.1312055290705944e-20

R84_93 V84 V93 497.72384606058506
L84_93 V84 V93 -2.378860300555734e-11
C84_93 V84 V93 -2.231807491268275e-20

R84_94 V84 V94 2825.3541353329033
L84_94 V84 V94 -9.554790103131673e-12
C84_94 V84 V94 -3.926505077964301e-20

R84_95 V84 V95 3906.6527131446155
L84_95 V84 V95 -3.7042300458638025e-11
C84_95 V84 V95 -2.4799711207926196e-20

R84_96 V84 V96 1079.3454861731316
L84_96 V84 V96 -2.1637258155909725e-12
C84_96 V84 V96 -4.443232212184614e-19

R84_97 V84 V97 2949.380758986655
L84_97 V84 V97 -1.6117450991871511e-12
C84_97 V84 V97 -3.2029596607721887e-19

R84_98 V84 V98 -552.2580648330453
L84_98 V84 V98 -1.6875094215495682e-12
C84_98 V84 V98 -2.6297947052288258e-19

R84_99 V84 V99 -903.8937815599758
L84_99 V84 V99 1.4950065113535034e-12
C84_99 V84 V99 2.1384726005769845e-19

R84_100 V84 V100 -293.45768906211777
L84_100 V84 V100 1.3231684211503253e-12
C84_100 V84 V100 3.840760315272567e-19

R84_101 V84 V101 -670.7424237748623
L84_101 V84 V101 1.8957044007989492e-12
C84_101 V84 V101 2.3716138762816665e-19

R84_102 V84 V102 1426.0570147799212
L84_102 V84 V102 3.4306223999615296e-12
C84_102 V84 V102 9.427782999594423e-20

R84_103 V84 V103 -10083.569126911481
L84_103 V84 V103 -3.783833701773234e-12
C84_103 V84 V103 -7.121345444970246e-20

R84_104 V84 V104 1285.865856385876
L84_104 V84 V104 -3.0871875092775237e-12
C84_104 V84 V104 5.103647754532167e-20

R84_105 V84 V105 564.8447544428294
L84_105 V84 V105 6.78903255317777e-12
C84_105 V84 V105 2.767571272437687e-21

R84_106 V84 V106 -1016.0086331757395
L84_106 V84 V106 1.8090757127246231e-12
C84_106 V84 V106 2.4593359498819023e-19

R84_107 V84 V107 5482.715997603693
L84_107 V84 V107 -3.172429442013054e-12
C84_107 V84 V107 -1.4062767994064057e-19

R84_108 V84 V108 685.0443074322621
L84_108 V84 V108 -2.4638461949639602e-11
C84_108 V84 V108 -1.4696597231078615e-19

R84_109 V84 V109 1577.2836603507071
L84_109 V84 V109 -1.894485978508468e-12
C84_109 V84 V109 -2.8403175095524733e-19

R84_110 V84 V110 1712.0378702941348
L84_110 V84 V110 -3.79144964384441e-12
C84_110 V84 V110 -1.062313957612904e-19

R84_111 V84 V111 -1757.7048805455945
L84_111 V84 V111 2.1035609830299605e-11
C84_111 V84 V111 6.281126290176727e-20

R84_112 V84 V112 -531.6397304886041
L84_112 V84 V112 -2.458684600063004e-12
C84_112 V84 V112 -2.250001628540522e-19

R84_113 V84 V113 -4074.2222858361542
L84_113 V84 V113 2.0219695737284414e-11
C84_113 V84 V113 1.0846574731834796e-19

R84_114 V84 V114 1052.8312757386866
L84_114 V84 V114 -2.1384894941307826e-12
C84_114 V84 V114 -2.0451009786448394e-19

R84_115 V84 V115 1332.1868228529327
L84_115 V84 V115 2.941904111934239e-12
C84_115 V84 V115 6.029847154395321e-20

R84_116 V84 V116 5510.206380978022
L84_116 V84 V116 1.6006798123714866e-12
C84_116 V84 V116 2.2922762560477243e-19

R84_117 V84 V117 16318.50612792871
L84_117 V84 V117 3.998679602979027e-12
C84_117 V84 V117 1.0832616793491814e-19

R84_118 V84 V118 -487.26859111101544
L84_118 V84 V118 3.1028785517000736e-12
C84_118 V84 V118 1.2269487686866582e-19

R84_119 V84 V119 -2319.364715235088
L84_119 V84 V119 1.811494669018294e-11
C84_119 V84 V119 2.365867459956779e-20

R84_120 V84 V120 6376.652933391968
L84_120 V84 V120 -2.3040213397513834e-11
C84_120 V84 V120 1.6876632051509012e-19

R84_121 V84 V121 1185.3909408792608
L84_121 V84 V121 1.405850560397367e-11
C84_121 V84 V121 -6.317732365064525e-20

R84_122 V84 V122 2048.7374333476287
L84_122 V84 V122 6.605045332793562e-12
C84_122 V84 V122 9.24044514483067e-20

R84_123 V84 V123 -2020.3970368762382
L84_123 V84 V123 -3.740068438359115e-12
C84_123 V84 V123 -6.56684794191609e-21

R84_124 V84 V124 -2053.858358764108
L84_124 V84 V124 -1.1853410968990028e-12
C84_124 V84 V124 -4.80683841713613e-19

R84_125 V84 V125 1512.7455816504894
L84_125 V84 V125 -3.997027429237306e-12
C84_125 V84 V125 -8.444132073395113e-20

R84_126 V84 V126 775.8245349093045
L84_126 V84 V126 -3.629705343113491e-12
C84_126 V84 V126 -3.603321676690884e-20

R84_127 V84 V127 1179.8008846752614
L84_127 V84 V127 -1.0730391067100482e-11
C84_127 V84 V127 -5.487496959267182e-20

R84_128 V84 V128 939.6332467552406
L84_128 V84 V128 1.5413463121197398e-12
C84_128 V84 V128 4.90308933688626e-20

R84_129 V84 V129 -5064.832078103748
L84_129 V84 V129 -2.3876858891383985e-11
C84_129 V84 V129 -7.617974116394036e-20

R84_130 V84 V130 -1132.2609333809976
L84_130 V84 V130 6.285629407901191e-12
C84_130 V84 V130 3.6903846271683125e-23

R84_131 V84 V131 -1031.9898174126663
L84_131 V84 V131 8.31926803015814e-12
C84_131 V84 V131 4.580014526325094e-20

R84_132 V84 V132 -456.4673943462534
L84_132 V84 V132 2.577098130408869e-11
C84_132 V84 V132 2.9552451516478617e-19

R84_133 V84 V133 -1730.727639902025
L84_133 V84 V133 4.897232883730145e-12
C84_133 V84 V133 1.6783916469959487e-19

R84_134 V84 V134 129225.05297418522
L84_134 V84 V134 -6.693946943744543e-12
C84_134 V84 V134 1.7143294712351685e-20

R84_135 V84 V135 2377.4618984261288
L84_135 V84 V135 -2.885861969236988e-11
C84_135 V84 V135 -1.1347488819710795e-20

R84_136 V84 V136 -3000.643634465517
L84_136 V84 V136 -2.034490056437814e-12
C84_136 V84 V136 -2.5086517542086446e-19

R84_137 V84 V137 674.3935427488728
L84_137 V84 V137 -5.126766349406679e-11
C84_137 V84 V137 6.517412775885731e-20

R84_138 V84 V138 930.6809936391973
L84_138 V84 V138 1.0541418261198757e-10
C84_138 V84 V138 2.4029578300231826e-20

R84_139 V84 V139 937.7203171154368
L84_139 V84 V139 2.4767650611104522e-12
C84_139 V84 V139 1.4201010377538451e-19

R84_140 V84 V140 345.0812568554158
L84_140 V84 V140 2.5975880766867555e-12
C84_140 V84 V140 1.7319893288255124e-19

R84_141 V84 V141 -1094.0180499970852
L84_141 V84 V141 -2.989627080380477e-12
C84_141 V84 V141 -2.6392566191496654e-19

R84_142 V84 V142 -991.9100417781435
L84_142 V84 V142 3.597023035307476e-12
C84_142 V84 V142 -1.8081730729475302e-20

R84_143 V84 V143 -491.9653590979795
L84_143 V84 V143 -2.5463261290323034e-12
C84_143 V84 V143 -9.788212544154302e-20

R84_144 V84 V144 -459.7133143009898
L84_144 V84 V144 -1.2742245409543053e-11
C84_144 V84 V144 -7.340816551489873e-21

R84_145 V84 V145 -1582.4606291335208
L84_145 V84 V145 -6.7135670424265e-12
C84_145 V84 V145 -8.283821638552961e-20

R84_146 V84 V146 -460.7953603953902
L84_146 V84 V146 -3.681958649587007e-12
C84_146 V84 V146 2.6636624114606978e-20

R84_147 V84 V147 2865.341325963544
L84_147 V84 V147 -3.3016591795389656e-12
C84_147 V84 V147 -1.5456646400456014e-19

R84_148 V84 V148 -963.8525339648033
L84_148 V84 V148 -4.6982953668088065e-12
C84_148 V84 V148 -1.119241465635496e-19

R84_149 V84 V149 -7464.488691502071
L84_149 V84 V149 9.841827122747622e-13
C84_149 V84 V149 3.422742001855325e-19

R84_150 V84 V150 705.6733300156692
L84_150 V84 V150 -2.780823301887912e-12
C84_150 V84 V150 -2.2263470340384255e-19

R84_151 V84 V151 801.4269720374715
L84_151 V84 V151 2.420722062534421e-12
C84_151 V84 V151 8.974114850200253e-20

R84_152 V84 V152 406.4091048751035
L84_152 V84 V152 1.8060764067791638e-12
C84_152 V84 V152 -6.502393921194159e-21

R84_153 V84 V153 334.1377661662538
L84_153 V84 V153 -6.09455836828442e-11
C84_153 V84 V153 2.728140935862324e-20

R84_154 V84 V154 436.45765096212426
L84_154 V84 V154 2.3238344505536685e-12
C84_154 V84 V154 1.1800043768385789e-19

R84_155 V84 V155 1941.8563887576247
L84_155 V84 V155 2.009857799757136e-12
C84_155 V84 V155 1.1755327929028538e-19

R84_156 V84 V156 -1657.9188545896284
L84_156 V84 V156 -1.0579840027997658e-12
C84_156 V84 V156 1.1694078384848862e-19

R84_157 V84 V157 15376.545827177908
L84_157 V84 V157 -7.760471733665746e-13
C84_157 V84 V157 -3.81788353027703e-19

R84_158 V84 V158 -392.69134734233927
L84_158 V84 V158 2.0222715890239837e-11
C84_158 V84 V158 3.5135730994200717e-20

R84_159 V84 V159 -506.57749464128193
L84_159 V84 V159 -1.5982189908981693e-12
C84_159 V84 V159 -6.413062135433319e-20

R84_160 V84 V160 -426.4687903043282
L84_160 V84 V160 4.321094268201829e-12
C84_160 V84 V160 2.3845826280982895e-20

R84_161 V84 V161 3253.7861781597776
L84_161 V84 V161 2.1730328134565557e-12
C84_161 V84 V161 3.278222881947329e-20

R84_162 V84 V162 -1491.578952301939
L84_162 V84 V162 9.07754679407005e-12
C84_162 V84 V162 3.73130712162822e-20

R84_163 V84 V163 2259.6954084921435
L84_163 V84 V163 -8.993732610876269e-12
C84_163 V84 V163 -3.276127031853814e-20

R84_164 V84 V164 2155.408150729514
L84_164 V84 V164 1.5104953907570586e-12
C84_164 V84 V164 1.3884766358597317e-20

R84_165 V84 V165 4636.331185702789
L84_165 V84 V165 3.5887713535619627e-12
C84_165 V84 V165 7.398456193394548e-20

R84_166 V84 V166 500.61191747122416
L84_166 V84 V166 6.64446343918197e-11
C84_166 V84 V166 -1.3910223050295573e-19

R84_167 V84 V167 -1882.6094462746785
L84_167 V84 V167 2.416721632840974e-12
C84_167 V84 V167 -1.702341752206003e-20

R84_168 V84 V168 688.0285006003079
L84_168 V84 V168 -1.3351242244673879e-12
C84_168 V84 V168 -3.4875338588534745e-20

R84_169 V84 V169 -3405.5755146359948
L84_169 V84 V169 -9.717622157878375e-12
C84_169 V84 V169 -2.9716465286986896e-20

R84_170 V84 V170 -697.0466507646693
L84_170 V84 V170 3.657742552144781e-11
C84_170 V84 V170 1.0092931975824789e-19

R84_171 V84 V171 7556.206177696825
L84_171 V84 V171 4.3672708340713876e-12
C84_171 V84 V171 8.071157400785124e-20

R84_172 V84 V172 -655.6296136429082
L84_172 V84 V172 -3.046879061545461e-12
C84_172 V84 V172 9.367857711047833e-20

R84_173 V84 V173 1469.6427065666355
L84_173 V84 V173 -9.457064414903094e-12
C84_173 V84 V173 -3.4623795237027015e-20

R84_174 V84 V174 -1185.2370248786433
L84_174 V84 V174 -5.835800288439381e-12
C84_174 V84 V174 -3.503321311405216e-20

R84_175 V84 V175 15910.455769263108
L84_175 V84 V175 -9.196396206469237e-12
C84_175 V84 V175 7.432400426746022e-20

R84_176 V84 V176 5553.652027363341
L84_176 V84 V176 1.0649073036645238e-12
C84_176 V84 V176 1.4503852612464464e-19

R84_177 V84 V177 -48929.42154670717
L84_177 V84 V177 -2.990886187050117e-12
C84_177 V84 V177 -3.783626651935939e-20

R84_178 V84 V178 716.3874035789054
L84_178 V84 V178 -5.3326302013246835e-12
C84_178 V84 V178 -6.030356147082767e-20

R84_179 V84 V179 -10669.149483381336
L84_179 V84 V179 -2.083490062865753e-12
C84_179 V84 V179 -1.6020969377954282e-19

R84_180 V84 V180 798.7789425532375
L84_180 V84 V180 -2.468380343619851e-12
C84_180 V84 V180 -2.3711790645548993e-19

R84_181 V84 V181 -1020.542776109113
L84_181 V84 V181 1.3650921330741096e-11
C84_181 V84 V181 -1.3117802091900582e-20

R84_182 V84 V182 -4869.529357233942
L84_182 V84 V182 2.2120090154728134e-12
C84_182 V84 V182 1.0202938936530623e-19

R84_183 V84 V183 -1732.5329028234783
L84_183 V84 V183 -3.1148747521514895e-12
C84_183 V84 V183 -1.9483282104562234e-20

R84_184 V84 V184 -698.9897805690177
L84_184 V84 V184 -1.104588979843732e-12
C84_184 V84 V184 2.7650165644903645e-20

R84_185 V84 V185 899.048243258691
L84_185 V84 V185 2.459941699387779e-12
C84_185 V84 V185 4.7855477283913176e-20

R84_186 V84 V186 -809.6435701765736
L84_186 V84 V186 -7.143312737809947e-12
C84_186 V84 V186 -4.2363774681462517e-20

R84_187 V84 V187 1780.1143099553824
L84_187 V84 V187 2.3241848549295536e-12
C84_187 V84 V187 1.2550364325809358e-19

R84_188 V84 V188 636.3594627172189
L84_188 V84 V188 6.22928737814142e-13
C84_188 V84 V188 1.9112573077340964e-19

R84_189 V84 V189 -1675.0053264033218
L84_189 V84 V189 -8.262941011909387e-12
C84_189 V84 V189 1.0088937593062548e-20

R84_190 V84 V190 3134.1283014350233
L84_190 V84 V190 -3.64484464163847e-12
C84_190 V84 V190 -1.1478912593863099e-19

R84_191 V84 V191 738.6813795967504
L84_191 V84 V191 1.51105219885387e-12
C84_191 V84 V191 6.211511402776184e-21

R84_192 V84 V192 1089.5978092458656
L84_192 V84 V192 -2.3562846411007405e-11
C84_192 V84 V192 -1.2436470734492008e-19

R84_193 V84 V193 -5585.789697799139
L84_193 V84 V193 -2.5456831164928896e-12
C84_193 V84 V193 -3.7154841587074807e-20

R84_194 V84 V194 2932.493975832893
L84_194 V84 V194 3.870016126094914e-11
C84_194 V84 V194 -4.491559637544428e-20

R84_195 V84 V195 -870.7596903114445
L84_195 V84 V195 -1.210971493004571e-12
C84_195 V84 V195 -1.444317550371367e-19

R84_196 V84 V196 -636.4303113000414
L84_196 V84 V196 -1.6565782960530528e-12
C84_196 V84 V196 8.958647343038924e-20

R84_197 V84 V197 2239.7496170093577
L84_197 V84 V197 -2.5980216597469932e-11
C84_197 V84 V197 -2.4581203969018783e-20

R84_198 V84 V198 -1572.5497535609416
L84_198 V84 V198 -4.54604431526985e-11
C84_198 V84 V198 -6.970426602821455e-20

R84_199 V84 V199 -676.3414754384179
L84_199 V84 V199 -2.3045169966863418e-12
C84_199 V84 V199 -6.791064376459368e-20

R84_200 V84 V200 -95477.57871133016
L84_200 V84 V200 -5.4593173530810296e-12
C84_200 V84 V200 7.053523189835036e-20

R85_85 V85 0 -834.1303635805851
L85_85 V85 0 5.297170272259897e-13
C85_85 V85 0 6.270621339940209e-19

R85_86 V85 V86 -708.454531825036
L85_86 V85 V86 -6.551575396386471e-12
C85_86 V85 V86 -1.7108866867846235e-19

R85_87 V85 V87 -5391.826294498321
L85_87 V85 V87 4.0209128761186436e-12
C85_87 V85 V87 1.0632111732346935e-19

R85_88 V85 V88 -5352.138069898675
L85_88 V85 V88 4.023440966213554e-12
C85_88 V85 V88 7.914978764055362e-20

R85_89 V85 V89 -803.2590749116815
L85_89 V85 V89 1.8208264855443047e-12
C85_89 V85 V89 3.3688171739474643e-19

R85_90 V85 V90 610.7475877803076
L85_90 V85 V90 8.868562539096541e-12
C85_90 V85 V90 1.7357723444757848e-21

R85_91 V85 V91 981.679859938446
L85_91 V85 V91 -1.7046252822662932e-12
C85_91 V85 V91 -2.855984933490238e-19

R85_92 V85 V92 1916.167088995526
L85_92 V85 V92 -2.0289109747443093e-12
C85_92 V85 V92 -1.8276206051824116e-19

R85_93 V85 V93 379.73624028862594
L85_93 V85 V93 1.495580639653321e-12
C85_93 V85 V93 4.076164475639925e-19

R85_94 V85 V94 6388.580467383832
L85_94 V85 V94 7.633625909009863e-12
C85_94 V85 V94 1.893174523004783e-19

R85_95 V85 V95 -3920.3699328842135
L85_95 V85 V95 1.6603361157736413e-11
C85_95 V85 V95 -2.512357192828647e-21

R85_96 V85 V96 -7299.55243857809
L85_96 V85 V96 6.1643386560591675e-12
C85_96 V85 V96 2.0747458676230085e-20

R85_97 V85 V97 -1810.680528983859
L85_97 V85 V97 -1.4458022474867353e-12
C85_97 V85 V97 -2.5812318369729634e-19

R85_98 V85 V98 -684.5766684360017
L85_98 V85 V98 -4.497703108079348e-12
C85_98 V85 V98 -1.599365740296251e-19

R85_99 V85 V99 -1296.4501780808032
L85_99 V85 V99 1.5867073135963959e-12
C85_99 V85 V99 3.535943375783601e-19

R85_100 V85 V100 -3617.1388540501875
L85_100 V85 V100 2.869367980181516e-12
C85_100 V85 V100 2.41302064430153e-19

R85_101 V85 V101 -550.3864858103715
L85_101 V85 V101 4.008432442220609e-12
C85_101 V85 V101 4.266983127824495e-20

R85_102 V85 V102 1792.7933835851084
L85_102 V85 V102 -2.5020992289378065e-10
C85_102 V85 V102 -9.328012691112392e-20

R85_103 V85 V103 2737.6183999405393
L85_103 V85 V103 -4.073487855638795e-12
C85_103 V85 V103 -1.5882940243802965e-19

R85_104 V85 V104 13548.14000518475
L85_104 V85 V104 -4.77819430822736e-12
C85_104 V85 V104 -1.399658644881739e-19

R85_105 V85 V105 421.70289818017227
L85_105 V85 V105 -1.1136168889797302e-11
C85_105 V85 V105 -1.6541055075646026e-19

R85_106 V85 V106 3315.428139658001
L85_106 V85 V106 3.031574746397843e-12
C85_106 V85 V106 3.0247284467698653e-19

R85_107 V85 V107 -155290.6478206753
L85_107 V85 V107 -3.658965278600561e-12
C85_107 V85 V107 -1.5537452530990636e-19

R85_108 V85 V108 -4830.381611660636
L85_108 V85 V108 -1.2371857442383997e-11
C85_108 V85 V108 -9.018620049903182e-20

R85_109 V85 V109 2860.8753605587785
L85_109 V85 V109 -3.2215919126825675e-12
C85_109 V85 V109 -1.0637399857574509e-19

R85_110 V85 V110 -1793.9621178168043
L85_110 V85 V110 -1.482471146580874e-11
C85_110 V85 V110 -1.1939287040871352e-19

R85_111 V85 V111 -10420.238850006423
L85_111 V85 V111 -2.010715553657404e-11
C85_111 V85 V111 3.768998608138878e-20

R85_112 V85 V112 10162.369698402694
L85_112 V85 V112 -7.175199829493231e-12
C85_112 V85 V112 5.4771757507136026e-21

R85_113 V85 V113 -571.6004319633312
L85_113 V85 V113 1.852528180651767e-11
C85_113 V85 V113 2.9242363001685833e-19

R85_114 V85 V114 6130.436884364019
L85_114 V85 V114 -2.821717177453324e-12
C85_114 V85 V114 -1.7704707605681842e-19

R85_115 V85 V115 10743.416096364674
L85_115 V85 V115 2.537157163981587e-12
C85_115 V85 V115 1.138832699301895e-19

R85_116 V85 V116 6517.927971935922
L85_116 V85 V116 2.9314735516482776e-12
C85_116 V85 V116 1.398308937767852e-19

R85_117 V85 V117 1562.3100498941976
L85_117 V85 V117 2.171688453808669e-12
C85_117 V85 V117 1.3259269347684587e-20

R85_118 V85 V118 -5570.556015098401
L85_118 V85 V118 4.532705412561929e-12
C85_118 V85 V118 1.0220968443878954e-19

R85_119 V85 V119 -4050.98288028235
L85_119 V85 V119 2.7058582897148906e-11
C85_119 V85 V119 2.7393042255514264e-20

R85_120 V85 V120 -3358.505524030764
L85_120 V85 V120 8.59714884585501e-12
C85_120 V85 V120 4.2684907356947e-20

R85_121 V85 V121 961.1565584607777
L85_121 V85 V121 -2.001938925557856e-12
C85_121 V85 V121 -2.6738377130765e-19

R85_122 V85 V122 5143.17954421082
L85_122 V85 V122 7.632982080376006e-12
C85_122 V85 V122 1.0391002159091889e-19

R85_123 V85 V123 5199.395160324435
L85_123 V85 V123 -2.597775891480134e-12
C85_123 V85 V123 -1.8060134991908217e-19

R85_124 V85 V124 3945.108943074807
L85_124 V85 V124 -1.9004840029453356e-12
C85_124 V85 V124 -2.6937450309238277e-19

R85_125 V85 V125 2643.268570712187
L85_125 V85 V125 2.5619593627656503e-12
C85_125 V85 V125 2.325067718075106e-19

R85_126 V85 V126 5411.300496548896
L85_126 V85 V126 -3.8480800678313934e-12
C85_126 V85 V126 -8.248087117744756e-20

R85_127 V85 V127 55601.84691561574
L85_127 V85 V127 1.671843819883152e-11
C85_127 V85 V127 2.4767961677186687e-20

R85_128 V85 V128 -5733.850227334437
L85_128 V85 V128 9.356714923704981e-12
C85_128 V85 V128 4.0171344769719426e-20

R85_129 V85 V129 -1129.3877412586219
L85_129 V85 V129 -2.772389202586975e-12
C85_129 V85 V129 -3.3244442204611085e-19

R85_130 V85 V130 -1388.5652710429779
L85_130 V85 V130 6.715245553684884e-11
C85_130 V85 V130 -1.0117575864877356e-19

R85_131 V85 V131 -2391.3412236366853
L85_131 V85 V131 5.217571411889814e-12
C85_131 V85 V131 1.0188632874745334e-19

R85_132 V85 V132 -2496.277175213637
L85_132 V85 V132 2.9298326197309748e-12
C85_132 V85 V132 1.5620706391781286e-19

R85_133 V85 V133 -1470.5076559186589
L85_133 V85 V133 1.890234857246468e-11
C85_133 V85 V133 3.7702662461284167e-19

R85_134 V85 V134 1318.629454561566
L85_134 V85 V134 8.887447731047537e-12
C85_134 V85 V134 2.3673319961621767e-19

R85_135 V85 V135 1199.5563409658037
L85_135 V85 V135 -5.531835402452265e-12
C85_135 V85 V135 -1.2358204197169256e-19

R85_136 V85 V136 980.3826236163302
L85_136 V85 V136 -5.621784480993171e-12
C85_136 V85 V136 -8.542088358319194e-20

R85_137 V85 V137 475.700695987615
L85_137 V85 V137 2.46822161362999e-12
C85_137 V85 V137 4.3810185991406804e-20

R85_138 V85 V138 6331.361442053295
L85_138 V85 V138 -2.473322947217522e-11
C85_138 V85 V138 -1.2598346692830779e-19

R85_139 V85 V139 -3134.1342458535523
L85_139 V85 V139 4.122096393822431e-12
C85_139 V85 V139 1.8101794236494324e-19

R85_140 V85 V140 -3993.180268041968
L85_140 V85 V140 8.080989658478859e-12
C85_140 V85 V140 1.6602144532197523e-19

R85_141 V85 V141 8839.659859612662
L85_141 V85 V141 -1.5389871642570543e-12
C85_141 V85 V141 -2.7879921693673706e-19

R85_142 V85 V142 -620.0813178617547
L85_142 V85 V142 -4.346877330759858e-12
C85_142 V85 V142 -1.142327356417021e-19

R85_143 V85 V143 -849.4026402414967
L85_143 V85 V143 -5.686485706728041e-12
C85_143 V85 V143 -9.283300418785813e-21

R85_144 V85 V144 -568.4118792515662
L85_144 V85 V144 -8.626145801425458e-12
C85_144 V85 V144 -9.380238456260204e-20

R85_145 V85 V145 -420.3743907146937
L85_145 V85 V145 7.539667818867616e-12
C85_145 V85 V145 1.0950160590671514e-19

R85_146 V85 V146 -1671.8867936219854
L85_146 V85 V146 9.2916345613584e-12
C85_146 V85 V146 9.165906240137626e-20

R85_147 V85 V147 5371.666536453669
L85_147 V85 V147 -7.356838915527445e-12
C85_147 V85 V147 -2.2610658847808523e-19

R85_148 V85 V148 843.7041847685566
L85_148 V85 V148 -2.9015794050339073e-12
C85_148 V85 V148 -1.3875626640650733e-19

R85_149 V85 V149 2386.8392414838795
L85_149 V85 V149 2.0849712694283284e-12
C85_149 V85 V149 -7.641075966818054e-20

R85_150 V85 V150 387.9339786066368
L85_150 V85 V150 -3.29242560940123e-11
C85_150 V85 V150 7.054085054447997e-22

R85_151 V85 V151 574.8568056271914
L85_151 V85 V151 3.3473315741156255e-11
C85_151 V85 V151 3.6865196340276425e-20

R85_152 V85 V152 1003.3987967324083
L85_152 V85 V152 3.98566133532547e-12
C85_152 V85 V152 7.31910333095674e-20

R85_153 V85 V153 412.17117692758137
L85_153 V85 V153 -5.297398696775351e-12
C85_153 V85 V153 -4.1304284639358396e-20

R85_154 V85 V154 1139.1861354836071
L85_154 V85 V154 7.134636897629296e-12
C85_154 V85 V154 -4.432514189849724e-20

R85_155 V85 V155 -683.1241216873754
L85_155 V85 V155 2.857882432432767e-12
C85_155 V85 V155 1.0071098701554684e-19

R85_156 V85 V156 -33736.68062144283
L85_156 V85 V156 9.596562865959528e-11
C85_156 V85 V156 1.075164245301833e-19

R85_157 V85 V157 1402.1958780559319
L85_157 V85 V157 -3.932521095701907e-12
C85_157 V85 V157 1.9734596982485257e-19

R85_158 V85 V158 -485.2263696962113
L85_158 V85 V158 -2.1704506340855126e-11
C85_158 V85 V158 7.991484931638568e-20

R85_159 V85 V159 -2801.4361265289504
L85_159 V85 V159 -4.8441966998361e-12
C85_159 V85 V159 -3.5010634093866696e-20

R85_160 V85 V160 -513.9971574881317
L85_160 V85 V160 -2.333865116488306e-11
C85_160 V85 V160 -3.859229738503995e-20

R85_161 V85 V161 -1343.0754205872242
L85_161 V85 V161 3.4918494016824837e-12
C85_161 V85 V161 -5.0051101049454704e-20

R85_162 V85 V162 -1948.4659962245748
L85_162 V85 V162 6.0769830122249474e-12
C85_162 V85 V162 5.904636578730395e-20

R85_163 V85 V163 2313.2379040227424
L85_163 V85 V163 6.676984896289703e-12
C85_163 V85 V163 8.387677266709484e-20

R85_164 V85 V164 866.6822911661407
L85_164 V85 V164 4.7287439780212154e-11
C85_164 V85 V164 1.446824868828893e-20

R85_165 V85 V165 2601.6315794912566
L85_165 V85 V165 -8.04697252985693e-12
C85_165 V85 V165 -5.0183770836246507e-20

R85_166 V85 V166 356.5248804507237
L85_166 V85 V166 -4.327097675582583e-12
C85_166 V85 V166 -1.229240946570839e-19

R85_167 V85 V167 12671.661481893207
L85_167 V85 V167 -1.5572908703747916e-11
C85_167 V85 V167 -2.81671648738456e-20

R85_168 V85 V168 -1661.241786755684
L85_168 V85 V168 9.101135627941535e-12
C85_168 V85 V168 -4.665869995991468e-20

R85_169 V85 V169 1558.4819092570403
L85_169 V85 V169 -3.7971452028470336e-12
C85_169 V85 V169 -6.189758382589269e-20

R85_170 V85 V170 -662.0568177481103
L85_170 V85 V170 3.012272000747188e-12
C85_170 V85 V170 -9.879160531675244e-21

R85_171 V85 V171 -1648.582850174501
L85_171 V85 V171 -2.4078137763676994e-11
C85_171 V85 V171 -1.413619817674365e-19

R85_172 V85 V172 -1500.6902591453654
L85_172 V85 V172 -3.6263166029218333e-12
C85_172 V85 V172 -7.134278359772716e-20

R85_173 V85 V173 -2439.725855832354
L85_173 V85 V173 1.5667438781863612e-12
C85_173 V85 V173 1.699706626360268e-19

R85_174 V85 V174 -552.1281064765819
L85_174 V85 V174 1.3016440499581058e-10
C85_174 V85 V174 9.691248448066505e-20

R85_175 V85 V175 1861.9768414605435
L85_175 V85 V175 8.905928300644842e-12
C85_175 V85 V175 1.7836820417715981e-19

R85_176 V85 V176 1122.5676474219533
L85_176 V85 V176 3.4851407169059947e-12
C85_176 V85 V176 2.184280308954232e-19

R85_177 V85 V177 2955.5836148511344
L85_177 V85 V177 -1.2626222187391111e-12
C85_177 V85 V177 -2.678767897389693e-19

R85_178 V85 V178 549.6306069426065
L85_178 V85 V178 -2.5122638708338276e-12
C85_178 V85 V178 7.75363510521157e-22

R85_179 V85 V179 -3553.4788067359964
L85_179 V85 V179 -2.7835856009403124e-11
C85_179 V85 V179 -2.1938600588202096e-20

R85_180 V85 V180 -12915.50904983846
L85_180 V85 V180 -8.463990159279889e-12
C85_180 V85 V180 -8.65792605852607e-20

R85_181 V85 V181 -22823.55382317692
L85_181 V85 V181 1.4462842703408547e-12
C85_181 V85 V181 1.1023081093568372e-19

R85_182 V85 V182 11541.86926023117
L85_182 V85 V182 3.920610828620747e-12
C85_182 V85 V182 -1.2381055957762473e-20

R85_183 V85 V183 -8510.895155855502
L85_183 V85 V183 -5.6019762728035865e-12
C85_183 V85 V183 -3.4769164508636094e-20

R85_184 V85 V184 -2121.2626743764795
L85_184 V85 V184 -4.204441051790725e-12
C85_184 V85 V184 -5.529120574387184e-20

R85_185 V85 V185 -12654.99288646102
L85_185 V85 V185 1.0720378505448889e-11
C85_185 V85 V185 1.789483450041019e-19

R85_186 V85 V186 -964.7530552831673
L85_186 V85 V186 -5.763022989869929e-12
C85_186 V85 V186 -1.4549249393756814e-19

R85_187 V85 V187 11530.613140801337
L85_187 V85 V187 2.191639695364904e-11
C85_187 V85 V187 5.461021656232928e-20

R85_188 V85 V188 2038.9712639854185
L85_188 V85 V188 2.464855268464088e-12
C85_188 V85 V188 5.356484602790977e-20

R85_189 V85 V189 -110583.28028086598
L85_189 V85 V189 -1.1800370315176884e-12
C85_189 V85 V189 -1.551125956634808e-19

R85_190 V85 V190 2102.8378160516595
L85_190 V85 V190 -2.4475805354543072e-11
C85_190 V85 V190 6.754441841614514e-20

R85_191 V85 V191 1622.404363455569
L85_191 V85 V191 2.3689676460872633e-11
C85_191 V85 V191 -1.111377733041709e-19

R85_192 V85 V192 4770.252198488601
L85_192 V85 V192 -3.4076882292883226e-12
C85_192 V85 V192 -1.0923348046052078e-19

R85_193 V85 V193 46302.262026496486
L85_193 V85 V193 1.0982161929523404e-12
C85_193 V85 V193 7.14966736483416e-20

R85_194 V85 V194 -4884.953416325648
L85_194 V85 V194 -5.3165191615368935e-12
C85_194 V85 V194 -2.800485801399082e-20

R85_195 V85 V195 -1898.0064754927528
L85_195 V85 V195 -3.939124921818126e-12
C85_195 V85 V195 9.819122728208571e-20

R85_196 V85 V196 -14994.376373028163
L85_196 V85 V196 -5.788929416715508e-11
C85_196 V85 V196 1.9531405866935996e-19

R85_197 V85 V197 -4674.488573571992
L85_197 V85 V197 -2.0786527024515337e-12
C85_197 V85 V197 -1.5807204598556927e-19

R85_198 V85 V198 3278.9089756985018
L85_198 V85 V198 1.0879488911099766e-11
C85_198 V85 V198 -7.539183451079929e-20

R85_199 V85 V199 5853.127407358731
L85_199 V85 V199 4.80138766016522e-12
C85_199 V85 V199 8.687636965845796e-20

R85_200 V85 V200 -1929.527970817215
L85_200 V85 V200 6.900136600264266e-12
C85_200 V85 V200 -3.917344370558796e-20

R86_86 V86 0 96.35713435582792
L86_86 V86 0 3.958052880818357e-12
C86_86 V86 0 -3.0827314753663715e-19

R86_87 V86 V87 -443.49578275956645
L86_87 V86 V87 2.7489889266173386e-12
C86_87 V86 V87 2.20690267593677e-19

R86_88 V86 V88 -371.0317220405744
L86_88 V86 V88 3.0584916496275058e-12
C86_88 V86 V88 2.0434392974053174e-19

R86_89 V86 V89 -277.0905680585763
L86_89 V86 V89 -3.746556879533384e-11
C86_89 V86 V89 7.147915409219267e-20

R86_90 V86 V90 97.59637794765986
L86_90 V86 V90 9.072573973751973e-13
C86_90 V86 V90 5.257354956157973e-19

R86_91 V86 V91 216.04173344538341
L86_91 V86 V91 -1.6747593982835333e-12
C86_91 V86 V91 -3.327680828791827e-19

R86_92 V86 V92 322.6233047220218
L86_92 V86 V92 -1.538185383418802e-12
C86_92 V86 V92 -3.10599526817984e-19

R86_93 V86 V93 202.63711190896646
L86_93 V86 V93 3.4553013923844943e-12
C86_93 V86 V93 1.5144765167077392e-19

R86_94 V86 V94 367.9132846264121
L86_94 V86 V94 1.7611352605233126e-12
C86_94 V86 V94 2.726499979100036e-19

R86_95 V86 V95 1516.2149787696985
L86_95 V86 V95 2.6644427116685588e-11
C86_95 V86 V95 -6.335562038043263e-20

R86_96 V86 V96 614.063478405972
L86_96 V86 V96 4.4077480566990706e-12
C86_96 V86 V96 -2.5018571670494182e-20

R86_97 V86 V97 4993.207039615938
L86_97 V86 V97 -1.460670551841127e-11
C86_97 V86 V97 -1.7254880884620106e-19

R86_98 V86 V98 -117.86867865853444
L86_98 V86 V98 -9.078338028736146e-13
C86_98 V86 V98 -4.702070221875465e-19

R86_99 V86 V99 -277.02329204168
L86_99 V86 V99 1.4051170292637918e-12
C86_99 V86 V99 3.9378461165564546e-19

R86_100 V86 V100 -442.900571215298
L86_100 V86 V100 1.858471411819206e-12
C86_100 V86 V100 4.2494360486440992e-19

R86_101 V86 V101 -968.6401685999615
L86_101 V86 V101 8.675909069647638e-12
C86_101 V86 V101 8.882104040253512e-20

R86_102 V86 V102 565.4845532827965
L86_102 V86 V102 -1.748560288142397e-11
C86_102 V86 V102 -7.028096327811532e-20

R86_103 V86 V103 -521.79933048239
L86_103 V86 V103 -1.6774533707386581e-12
C86_103 V86 V103 -2.6727741324940033e-19

R86_104 V86 V104 -284.7045890572622
L86_104 V86 V104 -1.703701277534838e-12
C86_104 V86 V104 -2.549584934998945e-19

R86_105 V86 V105 722.1498025475743
L86_105 V86 V105 -5.751278796990626e-12
C86_105 V86 V105 -1.5021593887400958e-19

R86_106 V86 V106 -426.77863329361475
L86_106 V86 V106 1.3656647115728319e-12
C86_106 V86 V106 4.253976807257766e-19

R86_107 V86 V107 293.339865052457
L86_107 V86 V107 4.041300381612214e-11
C86_107 V86 V107 -7.884789557702782e-20

R86_108 V86 V108 343.222704229845
L86_108 V86 V108 8.39824972877364e-12
C86_108 V86 V108 -8.064642202696055e-20

R86_109 V86 V109 -2403.8643132339243
L86_109 V86 V109 -3.928241729984146e-11
C86_109 V86 V109 -1.0822172711530288e-19

R86_110 V86 V110 204.1711622228887
L86_110 V86 V110 -6.466126635929772e-12
C86_110 V86 V110 2.917373568644649e-20

R86_111 V86 V111 1124.2563646908309
L86_111 V86 V111 1.1932828764573949e-11
C86_111 V86 V111 7.059036263176499e-20

R86_112 V86 V112 653.5855885849516
L86_112 V86 V112 -7.90387398487641e-12
C86_112 V86 V112 -6.934105631899107e-20

R86_113 V86 V113 223.56110545142846
L86_113 V86 V113 2.3758661158594065e-12
C86_113 V86 V113 3.6128066446448383e-19

R86_114 V86 V114 406.20561027387697
L86_114 V86 V114 -1.5487352401501385e-12
C86_114 V86 V114 -4.835321096520505e-19

R86_115 V86 V115 -312.10098595844227
L86_115 V86 V115 1.2585292421945911e-11
C86_115 V86 V115 3.165120405923776e-22

R86_116 V86 V116 -321.51290988773917
L86_116 V86 V116 4.674199014410834e-12
C86_116 V86 V116 1.1720936126977872e-19

R86_117 V86 V117 831.4551228217099
L86_117 V86 V117 1.1436837641838325e-09
C86_117 V86 V117 -8.729491537762148e-20

R86_118 V86 V118 -73.54887107154035
L86_118 V86 V118 6.050130555008827e-12
C86_118 V86 V118 1.9462217106579472e-19

R86_119 V86 V119 -616.1561716667561
L86_119 V86 V119 9.721597499132087e-12
C86_119 V86 V119 1.1363332689777e-19

R86_120 V86 V120 -1395.8994005618567
L86_120 V86 V120 5.768162150793646e-12
C86_120 V86 V120 1.7854149357178926e-19

R86_121 V86 V121 -216.02498500606018
L86_121 V86 V121 -2.778936211559167e-12
C86_121 V86 V121 -3.289869754164426e-19

R86_122 V86 V122 192.69022808843698
L86_122 V86 V122 2.2230817499985913e-12
C86_122 V86 V122 3.4707887873681733e-19

R86_123 V86 V123 490.2386858530692
L86_123 V86 V123 -2.0165532877239153e-12
C86_123 V86 V123 -2.742792269072681e-19

R86_124 V86 V124 519.5765063544641
L86_124 V86 V124 -1.459298963155363e-12
C86_124 V86 V124 -4.754394468715008e-19

R86_125 V86 V125 50513.766805265564
L86_125 V86 V125 5.279042825853444e-12
C86_125 V86 V125 2.3569322851386274e-19

R86_126 V86 V126 78.09964051039508
L86_126 V86 V126 -3.814969046081657e-12
C86_126 V86 V126 -3.4912962361663063e-19

R86_127 V86 V127 226.0098832833717
L86_127 V86 V127 4.801027757660831e-12
C86_127 V86 V127 1.0093836926840497e-19

R86_128 V86 V128 309.13578724309303
L86_128 V86 V128 4.0685483214712765e-12
C86_128 V86 V128 1.2077284124266612e-19

R86_129 V86 V129 126.38573898506068
L86_129 V86 V129 2.105147831245553e-12
C86_129 V86 V129 1.4075437446220466e-19

R86_130 V86 V130 -98.27804565380883
L86_130 V86 V130 -2.5691443840136056e-12
C86_130 V86 V130 -4.367290848813021e-20

R86_131 V86 V131 -136.59421612238845
L86_131 V86 V131 6.3571285076487714e-12
C86_131 V86 V131 1.5328096049023746e-19

R86_132 V86 V132 -114.60837175413137
L86_132 V86 V132 4.325059317916264e-12
C86_132 V86 V132 2.4198775309174522e-19

R86_133 V86 V133 -353.74500784196937
L86_133 V86 V133 -1.587152516112587e-12
C86_133 V86 V133 -2.590678666237758e-19

R86_134 V86 V134 -241.41916051179427
L86_134 V86 V134 1.334784091025125e-12
C86_134 V86 V134 5.640665634698737e-19

R86_135 V86 V135 -964.3709803629822
L86_135 V86 V135 -1.966188414843097e-12
C86_135 V86 V135 -3.6996501520432713e-19

R86_136 V86 V136 -374.0694113307418
L86_136 V86 V136 -2.237821461226348e-12
C86_136 V86 V136 -4.0306178115412713e-19

R86_137 V86 V137 -262.64655136584014
L86_137 V86 V137 -1.028033024865457e-11
C86_137 V86 V137 -6.350164807778167e-20

R86_138 V86 V138 123.42820929662993
L86_138 V86 V138 -1.51886725140139e-12
C86_138 V86 V138 -5.477041576078831e-19

R86_139 V86 V139 141.31564080764696
L86_139 V86 V139 1.790870859752748e-12
C86_139 V86 V139 3.643170909787561e-19

R86_140 V86 V140 91.17138536967481
L86_140 V86 V140 2.0319315318327306e-12
C86_140 V86 V140 4.472662733969132e-19

R86_141 V86 V141 -392.2997268860706
L86_141 V86 V141 2.363294561772289e-12
C86_141 V86 V141 2.509327620552556e-19

R86_142 V86 V142 382.3250437358149
L86_142 V86 V142 -1.6256855697554095e-12
C86_142 V86 V142 -4.791698841701611e-20

R86_143 V86 V143 -230.77356187388938
L86_143 V86 V143 -7.389282778591617e-12
C86_143 V86 V143 5.965371884291102e-20

R86_144 V86 V144 -221.79216717233473
L86_144 V86 V144 -7.1773224437780486e-12
C86_144 V86 V144 -1.9673523703549162e-20

R86_145 V86 V145 149.96508331004293
L86_145 V86 V145 -1.1470633531813643e-11
C86_145 V86 V145 2.1227781849942227e-20

R86_146 V86 V146 -135.36540004391637
L86_146 V86 V146 9.907905409123823e-13
C86_146 V86 V146 2.251230184055158e-19

R86_147 V86 V147 2153.231890403375
L86_147 V86 V147 -2.9660170910097446e-12
C86_147 V86 V147 -3.8379545157951028e-19

R86_148 V86 V148 -754.0290220895354
L86_148 V86 V148 -2.1007710455500494e-12
C86_148 V86 V148 -3.3263591354725526e-19

R86_149 V86 V149 894.934574667936
L86_149 V86 V149 -4.295781057217521e-12
C86_149 V86 V149 -3.7240520385725746e-19

R86_150 V86 V150 -130.67590854206043
L86_150 V86 V150 -9.464867997091059e-12
C86_150 V86 V150 1.6954494236852331e-19

R86_151 V86 V151 354.40380630700787
L86_151 V86 V151 7.532057138047456e-12
C86_151 V86 V151 1.808570194193337e-20

R86_152 V86 V152 142.16117967615938
L86_152 V86 V152 2.4171530452329284e-12
C86_152 V86 V152 1.155092258898793e-19

R86_153 V86 V153 -419.1621860345779
L86_153 V86 V153 1.4931764771831787e-11
C86_153 V86 V153 3.108199792655033e-20

R86_154 V86 V154 271.6681024933599
L86_154 V86 V154 -3.1160621502411288e-12
C86_154 V86 V154 -3.3431233486944214e-19

R86_155 V86 V155 -1528.3711957604698
L86_155 V86 V155 2.757276823096745e-12
C86_155 V86 V155 1.7879070517477504e-19

R86_156 V86 V156 -133.0896567169758
L86_156 V86 V156 -1.0552684876500641e-11
C86_156 V86 V156 1.7640157557013361e-19

R86_157 V86 V157 -166.73702622964376
L86_157 V86 V157 1.1152133159967073e-11
C86_157 V86 V157 2.85372865052206e-19

R86_158 V86 V158 292.17341768973847
L86_158 V86 V158 8.518794842710669e-12
C86_158 V86 V158 2.1289408478881185e-19

R86_159 V86 V159 -146.9595113143111
L86_159 V86 V159 -2.205589216744562e-12
C86_159 V86 V159 -1.8342383737033605e-19

R86_160 V86 V160 -154.23312648760506
L86_160 V86 V160 -3.1434044158770358e-12
C86_160 V86 V160 -1.8268885121813295e-19

R86_161 V86 V161 98.93242043718831
L86_161 V86 V161 2.624924240547578e-12
C86_161 V86 V161 9.527199621673661e-20

R86_162 V86 V162 196.60696347850015
L86_162 V86 V162 -4.99803156636758e-10
C86_162 V86 V162 -4.0476846834213413e-20

R86_163 V86 V163 117.12910931044594
L86_163 V86 V163 2.226307564595823e-12
C86_163 V86 V163 2.22169900165919e-19

R86_164 V86 V164 81.12541378787495
L86_164 V86 V164 3.68116983599058e-12
C86_164 V86 V164 1.2490037499917459e-19

R86_165 V86 V165 272.3769918101223
L86_165 V86 V165 -3.615976513946907e-12
C86_165 V86 V165 -3.272427326293131e-19

R86_166 V86 V166 -110.42448630732935
L86_166 V86 V166 -3.850159769355468e-12
C86_166 V86 V166 -1.6063913229378569e-19

R86_167 V86 V167 1383.4790642341168
L86_167 V86 V167 1.19150668574413e-11
C86_167 V86 V167 3.523334541532628e-20

R86_168 V86 V168 560.0738547145726
L86_168 V86 V168 2.5308990379674793e-12
C86_168 V86 V168 1.0995604795661237e-19

R86_169 V86 V169 -88.9469724173699
L86_169 V86 V169 -3.044804926182935e-12
C86_169 V86 V169 -7.639073992696649e-20

R86_170 V86 V170 -226.07700557534653
L86_170 V86 V170 7.157536029051617e-12
C86_170 V86 V170 -2.0082700965744966e-20

R86_171 V86 V171 -142.6785935773923
L86_171 V86 V171 -1.6517551037616772e-12
C86_171 V86 V171 -3.3761378416547044e-19

R86_172 V86 V172 -109.25345602446556
L86_172 V86 V172 -1.1908135820090748e-12
C86_172 V86 V172 -2.246769045645546e-19

R86_173 V86 V173 201.80067106609187
L86_173 V86 V173 2.5075742695050845e-12
C86_173 V86 V173 2.0198861727511633e-19

R86_174 V86 V174 103.47203726285028
L86_174 V86 V174 -8.517306942541315e-12
C86_174 V86 V174 1.4872539445975453e-19

R86_175 V86 V175 2059.2732880095905
L86_175 V86 V175 6.9095061411547335e-12
C86_175 V86 V175 1.507365059293024e-19

R86_176 V86 V176 480.9753541885146
L86_176 V86 V176 2.8617707099455562e-12
C86_176 V86 V176 2.0324833647113083e-19

R86_177 V86 V177 195.73131567735624
L86_177 V86 V177 5.629370753172088e-11
C86_177 V86 V177 -2.137619949086161e-19

R86_178 V86 V178 250.32886047470325
L86_178 V86 V178 5.772883319774244e-12
C86_178 V86 V178 5.768056231546024e-20

R86_179 V86 V179 280.85330713482153
L86_179 V86 V179 3.090604361051021e-12
C86_179 V86 V179 1.2666202144592927e-19

R86_180 V86 V180 213.17729935659764
L86_180 V86 V180 2.628808156218716e-12
C86_180 V86 V180 -1.7635600627287072e-20

R86_181 V86 V181 -156.9122768409149
L86_181 V86 V181 -4.342328402304826e-11
C86_181 V86 V181 1.324093792408694e-19

R86_182 V86 V182 -81.03614758511283
L86_182 V86 V182 -2.1106906992642254e-12
C86_182 V86 V182 -1.4834732237418437e-19

R86_183 V86 V183 -440.7021199408218
L86_183 V86 V183 -7.430364531588461e-12
C86_183 V86 V183 4.0083386685794015e-20

R86_184 V86 V184 -344.83872782563867
L86_184 V86 V184 -3.034609973872568e-12
C86_184 V86 V184 2.9733061845427106e-20

R86_185 V86 V185 -1394.9731058326634
L86_185 V86 V185 -7.542577428446472e-12
C86_185 V86 V185 9.252509177352108e-20

R86_186 V86 V186 -301.4168534799752
L86_186 V86 V186 -2.1406644518528e-12
C86_186 V86 V186 -5.747883942661533e-20

R86_187 V86 V187 773.3175064411835
L86_187 V86 V187 -1.3798917874979959e-11
C86_187 V86 V187 -1.8807659228671242e-20

R86_188 V86 V188 362.1008471567592
L86_188 V86 V188 3.198166854143415e-12
C86_188 V86 V188 -3.424221279271282e-20

R86_189 V86 V189 453.0028425030325
L86_189 V86 V189 -5.05891587167258e-12
C86_189 V86 V189 -3.232410541630154e-19

R86_190 V86 V190 116.66979483183123
L86_190 V86 V190 2.097288995347341e-12
C86_190 V86 V190 1.6367800259190012e-19

R86_191 V86 V191 304.01678893468113
L86_191 V86 V191 -8.60686439694872e-12
C86_191 V86 V191 -3.604399146027172e-19

R86_192 V86 V192 440.0414032471318
L86_192 V86 V192 -2.2329078829414e-12
C86_192 V86 V192 -3.7403623434709587e-19

R86_193 V86 V193 632.3537958764471
L86_193 V86 V193 2.6198999790054018e-12
C86_193 V86 V193 1.0827623300778963e-19

R86_194 V86 V194 -284.14063261960507
L86_194 V86 V194 -2.3211647856495765e-12
C86_194 V86 V194 -1.4977027020317955e-19

R86_195 V86 V195 -302.4576774604816
L86_195 V86 V195 4.837492219092168e-12
C86_195 V86 V195 4.338725421280334e-19

R86_196 V86 V196 -394.23260852797875
L86_196 V86 V196 1.549091206257814e-12
C86_196 V86 V196 6.287128813505902e-19

R86_197 V86 V197 -707.4849041897487
L86_197 V86 V197 4.1461613130311826e-12
C86_197 V86 V197 1.9630800438391613e-19

R86_198 V86 V198 -131.01931424815788
L86_198 V86 V198 -3.3681287463600775e-12
C86_198 V86 V198 -6.102913180577638e-20

R86_199 V86 V199 -334.6613786151392
L86_199 V86 V199 2.4123883585681212e-12
C86_199 V86 V199 2.3228288819036205e-19

R86_200 V86 V200 -4637.057053656828
L86_200 V86 V200 3.755759352076475e-12
C86_200 V86 V200 9.36657510795191e-20

R87_87 V87 0 193.0735936679275
L87_87 V87 0 -1.5118403092192174e-12
C87_87 V87 0 -4.1948468052493995e-19

R87_88 V87 V88 -557.5471915679393
L87_88 V87 V88 -5.013771237660843e-12
C87_88 V87 V88 -1.435965538511249e-19

R87_89 V87 V89 -722.8367085678199
L87_89 V87 V89 -2.1975495904225396e-12
C87_89 V87 V89 -2.381156607044943e-19

R87_90 V87 V90 1581.6362238907209
L87_90 V87 V90 -1.1932684564708866e-12
C87_90 V87 V90 -4.851266255588524e-19

R87_91 V87 V91 108.19136951629255
L87_91 V87 V91 4.520691101273824e-13
C87_91 V87 V91 1.0637359774962005e-18

R87_92 V87 V92 574.6218364553094
L87_92 V87 V92 3.8104110407870395e-11
C87_92 V87 V92 1.5180114763764276e-20

R87_93 V87 V93 2449.9522871812296
L87_93 V87 V93 -7.504761130883078e-12
C87_93 V87 V93 -4.7584371662707943e-20

R87_94 V87 V94 676.8022489534873
L87_94 V87 V94 -1.0169443632319763e-11
C87_94 V87 V94 -1.2765797469084394e-20

R87_95 V87 V95 226.24773840490923
L87_95 V87 V95 2.610563850823704e-12
C87_95 V87 V95 4.2932031369820037e-19

R87_96 V87 V96 635.8299839178046
L87_96 V87 V96 1.2053801580747761e-11
C87_96 V87 V96 9.587242222814216e-20

R87_97 V87 V97 755.6047589105805
L87_97 V87 V97 1.265446286533691e-12
C87_97 V87 V97 5.843068583102891e-19

R87_98 V87 V98 -778.87240511245
L87_98 V87 V98 1.377897707385041e-12
C87_98 V87 V98 4.333089108064267e-19

R87_99 V87 V99 -78.16174114250003
L87_99 V87 V99 -4.021193805170079e-13
C87_99 V87 V99 -1.2791277646076537e-18

R87_100 V87 V100 -466.7566854730183
L87_100 V87 V100 -8.99480934255132e-12
C87_100 V87 V100 -9.642867051321374e-20

R87_101 V87 V101 715.1099115376666
L87_101 V87 V101 -3.187855278298162e-12
C87_101 V87 V101 -3.2594940648863913e-19

R87_102 V87 V102 -855.9728392412499
L87_102 V87 V102 -1.4500053702806689e-11
C87_102 V87 V102 -2.4173925881329996e-20

R87_103 V87 V103 412.125150814814
L87_103 V87 V103 8.312888477496437e-13
C87_103 V87 V103 4.229071243898354e-19

R87_104 V87 V104 -832.9134940371487
L87_104 V87 V104 4.3798312895768505e-12
C87_104 V87 V104 1.2564595908539684e-19

R87_105 V87 V105 -364.71419142265546
L87_105 V87 V105 -2.790991372789889e-12
C87_105 V87 V105 -2.307904648590547e-19

R87_106 V87 V106 -1536.340545851861
L87_106 V87 V106 -1.0312483616149322e-12
C87_106 V87 V106 -6.146949664278444e-19

R87_107 V87 V107 120.89386300193769
L87_107 V87 V107 1.208185241350281e-12
C87_107 V87 V107 4.05337192813491e-19

R87_108 V87 V108 584.1820373857366
L87_108 V87 V108 -6.016109884850245e-12
C87_108 V87 V108 -1.3754943435732291e-19

R87_109 V87 V109 -497.7133620655427
L87_109 V87 V109 3.702838909024484e-12
C87_109 V87 V109 3.493333687676703e-19

R87_110 V87 V110 602.4201458820248
L87_110 V87 V110 2.3513814341999763e-12
C87_110 V87 V110 2.4750540108035605e-19

R87_111 V87 V111 -148.0078512023352
L87_111 V87 V111 -4.349708404070921e-12
C87_111 V87 V111 1.0107949645875215e-19

R87_112 V87 V112 -1344.7286597084596
L87_112 V87 V112 -3.0738555010412934e-12
C87_112 V87 V112 -1.6396587057663774e-19

R87_113 V87 V113 144.61048686718192
L87_113 V87 V113 3.5553327310916843e-12
C87_113 V87 V113 7.039887994848375e-20

R87_114 V87 V114 937.496901565677
L87_114 V87 V114 1.1730063178632395e-12
C87_114 V87 V114 5.485243155905093e-19

R87_115 V87 V115 -312.558156900596
L87_115 V87 V115 -7.876925656987716e-13
C87_115 V87 V115 -4.997150173893346e-19

R87_116 V87 V116 -890.425744068335
L87_116 V87 V116 3.124190865285754e-12
C87_116 V87 V116 2.9771262127499757e-19

R87_117 V87 V117 807.9781760987254
L87_117 V87 V117 -5.5603208447393276e-12
C87_117 V87 V117 -1.1281795219830252e-19

R87_118 V87 V118 -345.89759016333875
L87_118 V87 V118 -1.430361323986079e-12
C87_118 V87 V118 -4.321123813038291e-19

R87_119 V87 V119 174.75672988781892
L87_119 V87 V119 2.1799415030230436e-12
C87_119 V87 V119 -1.060989524290475e-19

R87_120 V87 V120 743.0088280218939
L87_120 V87 V120 -9.64197761881338e-12
C87_120 V87 V120 -1.9895154211831514e-19

R87_121 V87 V121 -162.10947098159326
L87_121 V87 V121 -6.326063438665874e-11
C87_121 V87 V121 9.223176735118708e-21

R87_122 V87 V122 13232.822322501344
L87_122 V87 V122 -4.345374408325153e-12
C87_122 V87 V122 -1.4399313592591071e-19

R87_123 V87 V123 -270.09621116234825
L87_123 V87 V123 7.628987974127238e-13
C87_123 V87 V123 9.7019094296814e-19

R87_124 V87 V124 -984.2581212094026
L87_124 V87 V124 -6.305365999927691e-12
C87_124 V87 V124 -8.338625708486058e-20

R87_125 V87 V125 -868.8633497899632
L87_125 V87 V125 -9.431456381905063e-12
C87_125 V87 V125 -1.0439664579120243e-19

R87_126 V87 V126 361.5796006512452
L87_126 V87 V126 1.4689195521739152e-12
C87_126 V87 V126 3.019948762476228e-19

R87_127 V87 V127 932.2191315323712
L87_127 V87 V127 -7.692682614222075e-13
C87_127 V87 V127 -5.882413232206991e-19

R87_128 V87 V128 -10137.800628264673
L87_128 V87 V128 4.6602581261644275e-12
C87_128 V87 V128 2.4060929713567015e-19

R87_129 V87 V129 148.362617618987
L87_129 V87 V129 7.461526843794661e-12
C87_129 V87 V129 1.823758338907475e-19

R87_130 V87 V130 -1387.496293046949
L87_130 V87 V130 -6.878023756017542e-12
C87_130 V87 V130 -5.2339926298684705e-21

R87_131 V87 V131 -2164.191598449112
L87_131 V87 V131 6.664991056525194e-12
C87_131 V87 V131 -1.9644408073287114e-19

R87_132 V87 V132 4860.367749747501
L87_132 V87 V132 -2.750491909538106e-12
C87_132 V87 V132 -3.8684098438913116e-19

R87_133 V87 V133 887.7517763276152
L87_133 V87 V133 1.3701416570461494e-11
C87_133 V87 V133 -1.836710599168817e-20

R87_134 V87 V134 3503.7881876504202
L87_134 V87 V134 -7.692048896866863e-12
C87_134 V87 V134 -1.9971381572676743e-19

R87_135 V87 V135 -145.84806080035625
L87_135 V87 V135 7.516384283923536e-13
C87_135 V87 V135 1.1774665466489309e-18

R87_136 V87 V136 -788.1357254096573
L87_136 V87 V136 -6.981054567033522e-12
C87_136 V87 V136 -5.425843479019771e-20

R87_137 V87 V137 -162.2612845348441
L87_137 V87 V137 1.1879009342143615e-10
C87_137 V87 V137 1.7247817059450683e-20

R87_138 V87 V138 5026.593906708141
L87_138 V87 V138 2.5983632225911015e-12
C87_138 V87 V138 3.0141916239244317e-19

R87_139 V87 V139 99.35022822229922
L87_139 V87 V139 -5.518590191455683e-13
C87_139 V87 V139 -1.4862912110979638e-18

R87_140 V87 V140 273.9671613712443
L87_140 V87 V140 2.9086172071271656e-12
C87_140 V87 V140 1.7965705474815982e-19

R87_141 V87 V141 -308.54355105812
L87_141 V87 V141 1.2640293985483422e-11
C87_141 V87 V141 7.590801982201933e-20

R87_142 V87 V142 -4045.556908501473
L87_142 V87 V142 -1.3040572016751209e-11
C87_142 V87 V142 -1.6661273923177357e-21

R87_143 V87 V143 510.7389915758019
L87_143 V87 V143 1.5274030052097558e-12
C87_143 V87 V143 2.5012800431648796e-19

R87_144 V87 V144 -1051.489809080783
L87_144 V87 V144 -9.534985174631287e-11
C87_144 V87 V144 -1.0653386169597266e-19

R87_145 V87 V145 121.81281120827931
L87_145 V87 V145 3.1157462662148995e-11
C87_145 V87 V145 -1.2274373168252546e-21

R87_146 V87 V146 823.2334640211601
L87_146 V87 V146 -4.746576109965902e-12
C87_146 V87 V146 -1.6434353033398443e-19

R87_147 V87 V147 -150.63978328279964
L87_147 V87 V147 2.527701135948953e-12
C87_147 V87 V147 9.255158181295143e-19

R87_148 V87 V148 884.0823425452978
L87_148 V87 V148 -3.225189590487464e-12
C87_148 V87 V148 -1.5836236374652256e-20

R87_149 V87 V149 816.6156056061363
L87_149 V87 V149 -2.501045614816319e-12
C87_149 V87 V149 -2.943003937091575e-19

R87_150 V87 V150 -358.3415603821836
L87_150 V87 V150 8.04796822683364e-12
C87_150 V87 V150 -2.860691855838691e-20

R87_151 V87 V151 -105.20231434231323
L87_151 V87 V151 -2.0114672359137702e-12
C87_151 V87 V151 -4.547526447176733e-19

R87_152 V87 V152 -4145.714857070697
L87_152 V87 V152 4.440923804262983e-12
C87_152 V87 V152 6.719520730289406e-20

R87_153 V87 V153 -272.50764513349276
L87_153 V87 V153 4.118831215324203e-12
C87_153 V87 V153 2.3846044163114576e-19

R87_154 V87 V154 -434.38991370802466
L87_154 V87 V154 9.480438474312732e-12
C87_154 V87 V154 1.7835740844256651e-19

R87_155 V87 V155 75.56690252672618
L87_155 V87 V155 -1.0275347965606643e-12
C87_155 V87 V155 -5.5744864219428805e-19

R87_156 V87 V156 -553.9996593823527
L87_156 V87 V156 -1.6124260402304808e-11
C87_156 V87 V156 8.100056252158311e-20

R87_157 V87 V157 -167.84151794529998
L87_157 V87 V157 5.843326804130802e-12
C87_157 V87 V157 1.7475171926303637e-19

R87_158 V87 V158 10123.3196684391
L87_158 V87 V158 -3.835851993323719e-12
C87_158 V87 V158 -1.4577875123689191e-19

R87_159 V87 V159 269.28953208038837
L87_159 V87 V159 7.052116539762024e-13
C87_159 V87 V159 6.906968621662417e-19

R87_160 V87 V160 -633.5281785148693
L87_160 V87 V160 2.442788494145507e-11
C87_160 V87 V160 -6.582965807935494e-20

R87_161 V87 V161 232.0404405882102
L87_161 V87 V161 -2.455603316120039e-12
C87_161 V87 V161 -3.1473895569810377e-19

R87_162 V87 V162 436.6712305320679
L87_162 V87 V162 -3.8600122767048515e-12
C87_162 V87 V162 -1.2818963237032987e-19

R87_163 V87 V163 -16411.301068341014
L87_163 V87 V163 -1.3989840564665205e-12
C87_163 V87 V163 -3.4086074062884864e-19

R87_164 V87 V164 288.57958313495845
L87_164 V87 V164 -1.4796452329296954e-11
C87_164 V87 V164 -8.333880078720827e-20

R87_165 V87 V165 219.31499685883787
L87_165 V87 V165 4.407050777912234e-12
C87_165 V87 V165 1.0169741642686448e-19

R87_166 V87 V166 -1805.457185218029
L87_166 V87 V166 1.4338559351811134e-11
C87_166 V87 V166 5.3505276171323307e-20

R87_167 V87 V167 -129.95664257308826
L87_167 V87 V167 7.545899380259766e-12
C87_167 V87 V167 -6.687581371329265e-20

R87_168 V87 V168 562.6705178932177
L87_168 V87 V168 -3.161805759397958e-12
C87_168 V87 V168 -1.4495664710750785e-19

R87_169 V87 V169 -249.19832009711638
L87_169 V87 V169 2.0736587941059423e-12
C87_169 V87 V169 3.6232832879172667e-19

R87_170 V87 V170 -1173.6297490467446
L87_170 V87 V170 3.20326583583665e-11
C87_170 V87 V170 -1.001888905303959e-20

R87_171 V87 V171 705.8736871519715
L87_171 V87 V171 2.965575887598022e-12
C87_171 V87 V171 1.8519846800106898e-19

R87_172 V87 V172 -519.2293099045473
L87_172 V87 V172 5.1759519692734814e-12
C87_172 V87 V172 1.3373346901997606e-19

R87_173 V87 V173 -687.1247490753864
L87_173 V87 V173 -1.803309371280882e-12
C87_173 V87 V173 -1.881246367844654e-19

R87_174 V87 V174 -5639.723623168007
L87_174 V87 V174 5.079631444051226e-12
C87_174 V87 V174 1.3701030701621943e-19

R87_175 V87 V175 253.3454430949532
L87_175 V87 V175 -9.517604724818835e-13
C87_175 V87 V175 -4.6482402786247565e-19

R87_176 V87 V176 1752.663183603289
L87_176 V87 V176 5.528230555377635e-12
C87_176 V87 V176 1.5034980593940872e-19

R87_177 V87 V177 450.477725708757
L87_177 V87 V177 2.3345694570545274e-12
C87_177 V87 V177 -8.611368662301513e-21

R87_178 V87 V178 -4421.965748740096
L87_178 V87 V178 2.0933093029549303e-11
C87_178 V87 V178 -2.009559842587763e-20

R87_179 V87 V179 241.59759286056277
L87_179 V87 V179 2.364297340437795e-12
C87_179 V87 V179 3.8363999424914275e-19

R87_180 V87 V180 9284.722967356493
L87_180 V87 V180 -1.1025766055078583e-10
C87_180 V87 V180 -4.7574866646907204e-20

R87_181 V87 V181 -1043.4722463407459
L87_181 V87 V181 -3.823725158423311e-12
C87_181 V87 V181 -1.0227959054960136e-19

R87_182 V87 V182 4310.933065122854
L87_182 V87 V182 -2.8792038379258682e-12
C87_182 V87 V182 -1.2410935840069504e-19

R87_183 V87 V183 -137.67308318040176
L87_183 V87 V183 1.62766180418867e-12
C87_183 V87 V183 1.5161246811436511e-21

R87_184 V87 V184 -3216.463878511474
L87_184 V87 V184 4.693510397722495e-12
C87_184 V87 V184 5.3885515643423074e-20

R87_185 V87 V185 -672.1815870903412
L87_185 V87 V185 -1.975118773798466e-12
C87_185 V87 V185 3.813591219219171e-20

R87_186 V87 V186 1894.3921255213013
L87_186 V87 V186 4.756660053972182e-12
C87_186 V87 V186 9.010131282134348e-20

R87_187 V87 V187 5510.181442782569
L87_187 V87 V187 -7.980692653406612e-13
C87_187 V87 V187 -4.750609860665779e-19

R87_188 V87 V188 800.8060512070566
L87_188 V87 V188 -2.721928143568678e-12
C87_188 V87 V188 -1.2596507540285077e-19

R87_189 V87 V189 1118.813763686809
L87_189 V87 V189 1.6059036804811943e-12
C87_189 V87 V189 1.877561380530799e-19

R87_190 V87 V190 -1833.3807293470106
L87_190 V87 V190 9.654015106313651e-12
C87_190 V87 V190 1.1432346548299767e-20

R87_191 V87 V191 197.07195963329454
L87_191 V87 V191 7.895700819905988e-12
C87_191 V87 V191 4.559135811037557e-19

R87_192 V87 V192 3972.2935116832414
L87_192 V87 V192 -3.4937350048112508e-12
C87_192 V87 V192 8.520110165510452e-20

R87_193 V87 V193 809.3219023673191
L87_193 V87 V193 6.240489612068728e-12
C87_193 V87 V193 -9.948189715095775e-21

R87_194 V87 V194 -1190.3470182682836
L87_194 V87 V194 7.809374248890356e-12
C87_194 V87 V194 2.3208945613324944e-19

R87_195 V87 V195 -265.40074618092945
L87_195 V87 V195 -6.851622481498615e-12
C87_195 V87 V195 -6.590545644537648e-19

R87_196 V87 V196 -465.98238554035953
L87_196 V87 V196 1.1317645477210312e-12
C87_196 V87 V196 2.996301210423912e-19

R87_197 V87 V197 -617.7365452428335
L87_197 V87 V197 -2.7949809519361843e-12
C87_197 V87 V197 -1.849997901361254e-19

R87_198 V87 V198 -1522.8079847837366
L87_198 V87 V198 -1.8179487174039163e-11
C87_198 V87 V198 -2.893298978765725e-20

R87_199 V87 V199 -366.6468326600806
L87_199 V87 V199 -1.0550137410584993e-11
C87_199 V87 V199 -5.031215672689951e-20

R87_200 V87 V200 -10087.84500057011
L87_200 V87 V200 -3.3855754012434794e-12
C87_200 V87 V200 -2.999321794650814e-19

R88_88 V88 0 71.5661067104162
L88_88 V88 0 -2.2360890463384523e-13
C88_88 V88 0 -2.5331959486091226e-18

R88_89 V88 V89 -459.94397012670737
L88_89 V88 V89 -1.0666537484555393e-12
C88_89 V88 V89 -4.153765400091198e-19

R88_90 V88 V90 917.9642091012917
L88_90 V88 V90 -7.704994782810957e-13
C88_90 V88 V90 -6.681200114297946e-19

R88_91 V88 V91 512.5126758935862
L88_91 V88 V91 3.642118792688475e-12
C88_91 V88 V91 1.5963109057265074e-19

R88_92 V88 V92 87.5971452056967
L88_92 V88 V92 4.023506156753168e-13
C88_92 V88 V92 9.558782814386276e-19

R88_93 V88 V93 2148.280997645795
L88_93 V88 V93 -1.9786180300232127e-11
C88_93 V88 V93 3.325646171319138e-20

R88_94 V88 V94 1041.7250375660756
L88_94 V88 V94 9.096711141294956e-12
C88_94 V88 V94 1.5076947347318962e-19

R88_95 V88 V95 748.1708469057673
L88_95 V88 V95 7.294018466690992e-12
C88_95 V88 V95 9.477108233362474e-20

R88_96 V88 V96 199.6732749370842
L88_96 V88 V96 4.817102396873665e-12
C88_96 V88 V96 4.887419343953345e-19

R88_97 V88 V97 662.5818195146345
L88_97 V88 V97 7.627218606965753e-13
C88_97 V88 V97 8.8023733294244e-19

R88_98 V88 V98 -1012.7764169326647
L88_98 V88 V98 9.435059113310845e-13
C88_98 V88 V98 5.60088423437837e-19

R88_99 V88 V99 -323.0659714397978
L88_99 V88 V99 -1.4088103233109347e-12
C88_99 V88 V99 -2.4768802978269927e-19

R88_100 V88 V100 -64.70136830428042
L88_100 V88 V100 -4.624918191432051e-13
C88_100 V88 V100 -1.2024337599104235e-18

R88_101 V88 V101 772.9950534171803
L88_101 V88 V101 -1.4975731146281403e-12
C88_101 V88 V101 -4.648030078756817e-19

R88_102 V88 V102 -906.7455824079996
L88_102 V88 V102 -2.5557907077377633e-12
C88_102 V88 V102 -2.0693746078714903e-19

R88_103 V88 V103 -920.2793827040595
L88_103 V88 V103 5.8723890438567e-12
C88_103 V88 V103 1.0429068200224448e-19

R88_104 V88 V104 582.6759534596702
L88_104 V88 V104 7.807260497474421e-13
C88_104 V88 V104 4.2344155832570797e-19

R88_105 V88 V105 -328.90169234039865
L88_105 V88 V105 -1.5517334314679333e-12
C88_105 V88 V105 -3.241322751039961e-19

R88_106 V88 V106 -690.5755372628523
L88_106 V88 V106 -1.114843873269505e-12
C88_106 V88 V106 -5.287076074580237e-19

R88_107 V88 V107 408.6805480598344
L88_107 V88 V107 2.6641670967875006e-12
C88_107 V88 V107 1.3770911699078175e-19

R88_108 V88 V108 87.15935888407805
L88_108 V88 V108 -1.7364373885059415e-11
C88_108 V88 V108 3.1959416104122137e-20

R88_109 V88 V109 -721.1759948959062
L88_109 V88 V109 1.8042121013557533e-12
C88_109 V88 V109 5.382719061079515e-19

R88_110 V88 V110 328.1892626371014
L88_110 V88 V110 2.8995919335861946e-12
C88_110 V88 V110 1.729713102490883e-19

R88_111 V88 V111 -2280.91787162149
L88_111 V88 V111 -3.639672902308293e-12
C88_111 V88 V111 -1.9035119179262553e-19

R88_112 V88 V112 -142.58842334771091
L88_112 V88 V112 1.2731132164943722e-12
C88_112 V88 V112 6.051116639609509e-19

R88_113 V88 V113 133.57275079191064
L88_113 V88 V113 1.9221705951683597e-12
C88_113 V88 V113 1.4910936924356874e-19

R88_114 V88 V114 1004.4266484492889
L88_114 V88 V114 9.556580733321156e-13
C88_114 V88 V114 5.715404883077616e-19

R88_115 V88 V115 -1171.2126017400258
L88_115 V88 V115 1.5854196459962325e-10
C88_115 V88 V115 1.0562993640126657e-19

R88_116 V88 V116 -141.184734142269
L88_116 V88 V116 -7.913283588172024e-13
C88_116 V88 V116 -4.087853096560417e-19

R88_117 V88 V117 1558.4802443219435
L88_117 V88 V117 -2.637469812209996e-12
C88_117 V88 V117 -2.2744685857074173e-19

R88_118 V88 V118 -196.41596613048887
L88_118 V88 V118 -1.1937436050796434e-12
C88_118 V88 V118 -4.860591373594329e-19

R88_119 V88 V119 9948.94778755901
L88_119 V88 V119 -3.1463114837380106e-12
C88_119 V88 V119 -3.143788977023839e-19

R88_120 V88 V120 98.39844207673481
L88_120 V88 V120 -3.876564688240344e-12
C88_120 V88 V120 -7.446175264796347e-19

R88_121 V88 V121 -178.60737408230833
L88_121 V88 V121 -4.398078410438683e-12
C88_121 V88 V121 -5.732521979899135e-20

R88_122 V88 V122 452.0232382603218
L88_122 V88 V122 -5.368568818493161e-12
C88_122 V88 V122 -1.591922299280733e-19

R88_123 V88 V123 2266.7176737831533
L88_123 V88 V123 5.5067183538242406e-12
C88_123 V88 V123 5.876870815686612e-20

R88_124 V88 V124 -232.51725214343523
L88_124 V88 V124 4.1100838858042557e-13
C88_124 V88 V124 1.588048773688911e-18

R88_125 V88 V125 -18090.993191208003
L88_125 V88 V125 7.53275529058657e-12
C88_125 V88 V125 -2.9188867412723093e-21

R88_126 V88 V126 214.90220489102936
L88_126 V88 V126 1.007128830045879e-12
C88_126 V88 V126 3.1573849452689875e-19

R88_127 V88 V127 417.3811824811774
L88_127 V88 V127 1.1577314478941686e-12
C88_127 V88 V127 4.479558660017508e-19

R88_128 V88 V128 -667.4649028126066
L88_128 V88 V128 -7.600001061199951e-13
C88_128 V88 V128 -3.6469876843725323e-19

R88_129 V88 V129 157.05923944902534
L88_129 V88 V129 3.22644900570431e-12
C88_129 V88 V129 3.3204625241718604e-19

R88_130 V88 V130 -325.0991310918031
L88_130 V88 V130 -1.9283382945251178e-12
C88_130 V88 V130 -1.4178927518442712e-19

R88_131 V88 V131 -311.5768073979289
L88_131 V88 V131 -1.2545306651346525e-12
C88_131 V88 V131 -4.2772390728155516e-19

R88_132 V88 V132 1186.863774858643
L88_132 V88 V132 -2.097418592173926e-12
C88_132 V88 V132 -6.842718979083586e-19

R88_133 V88 V133 1643.195108159268
L88_133 V88 V133 -3.0262912660755653e-12
C88_133 V88 V133 -3.3305951280929026e-19

R88_134 V88 V134 1542.3634278043035
L88_134 V88 V134 -5.46492134282969e-12
C88_134 V88 V134 -3.1825478424686052e-19

R88_135 V88 V135 6315.016968240533
L88_135 V88 V135 -2.3850851343962397e-12
C88_135 V88 V135 -2.404364645093324e-19

R88_136 V88 V136 -144.77139701380975
L88_136 V88 V136 6.404932855126902e-13
C88_136 V88 V136 1.2177513909630877e-18

R88_137 V88 V137 -167.24669212152943
L88_137 V88 V137 6.120574147506385e-12
C88_137 V88 V137 9.582926103991748e-20

R88_138 V88 V138 1144.3460683702833
L88_138 V88 V138 1.6305676825252617e-12
C88_138 V88 V138 3.864569673737013e-19

R88_139 V88 V139 320.66454541902954
L88_139 V88 V139 1.5066083659605628e-12
C88_139 V88 V139 3.112431574808184e-19

R88_140 V88 V140 98.6017120337895
L88_140 V88 V140 -7.330860568829291e-13
C88_140 V88 V140 -1.2474852915881212e-18

R88_141 V88 V141 -392.2525882423697
L88_141 V88 V141 2.2703373958432182e-12
C88_141 V88 V141 2.851537869443523e-19

R88_142 V88 V142 4946.08258234991
L88_142 V88 V142 -1.6657788092470446e-11
C88_142 V88 V142 9.97587231638346e-21

R88_143 V88 V143 -606.8047269453256
L88_143 V88 V143 3.441073916852698e-12
C88_143 V88 V143 7.051911098330911e-20

R88_144 V88 V144 217.35115176335597
L88_144 V88 V144 3.725330934654045e-12
C88_144 V88 V144 1.636255411257673e-19

R88_145 V88 V145 119.96213641362988
L88_145 V88 V145 -9.143157254710941e-12
C88_145 V88 V145 -5.509900622934536e-20

R88_146 V88 V146 857.3998009518457
L88_146 V88 V146 -2.2872869390174635e-12
C88_146 V88 V146 -1.8385943899921956e-19

R88_147 V88 V147 1920.886961281507
L88_147 V88 V147 3.722972951030507e-10
C88_147 V88 V147 1.1303812855536164e-19

R88_148 V88 V148 -75.8160379869602
L88_148 V88 V148 6.794513320230263e-13
C88_148 V88 V148 8.189649206533254e-19

R88_149 V88 V149 814.0156922776774
L88_149 V88 V149 -1.2242314419117253e-12
C88_149 V88 V149 -4.470297242321293e-19

R88_150 V88 V150 -251.96094981788792
L88_150 V88 V150 3.111928501912798e-12
C88_150 V88 V150 2.3271464640962306e-19

R88_151 V88 V151 -3676.9335646901473
L88_151 V88 V151 -2.1333978482559423e-12
C88_151 V88 V151 -1.1271524265448268e-19

R88_152 V88 V152 -413.739622055723
L88_152 V88 V152 -7.013908894102927e-13
C88_152 V88 V152 -2.8355777370036774e-19

R88_153 V88 V153 -237.81655476523036
L88_153 V88 V153 -5.329160235955362e-12
C88_153 V88 V153 1.4194408956523752e-19

R88_154 V88 V154 -655.5111487567239
L88_154 V88 V154 -2.8779810701634003e-12
C88_154 V88 V154 9.869274744483989e-21

R88_155 V88 V155 -983.895098111309
L88_155 V88 V155 -3.1004473239866624e-12
C88_155 V88 V155 -6.041712246714415e-20

R88_156 V88 V156 553.6141930416676
L88_156 V88 V156 2.5673051819841706e-12
C88_156 V88 V156 -6.335729791682733e-19

R88_157 V88 V157 -142.50652677898896
L88_157 V88 V157 7.562912454736207e-13
C88_157 V88 V157 6.485441996926011e-19

R88_158 V88 V158 -1122.7812784439793
L88_158 V88 V158 -3.7642871650273965e-11
C88_158 V88 V158 -1.0738141640582109e-19

R88_159 V88 V159 -247.42181875028837
L88_159 V88 V159 8.048204515528757e-12
C88_159 V88 V159 -2.840490174918568e-20

R88_160 V88 V160 94.79993621164535
L88_160 V88 V160 1.4180663607263143e-12
C88_160 V88 V160 4.692572896786794e-19

R88_161 V88 V161 207.328199966923
L88_161 V88 V161 -1.1813222580653748e-12
C88_161 V88 V161 -3.790910974383734e-19

R88_162 V88 V162 324.70797000982907
L88_162 V88 V162 -2.819859758830041e-12
C88_162 V88 V162 -8.494362394977423e-20

R88_163 V88 V163 227.95505818759077
L88_163 V88 V163 2.9584698849059624e-12
C88_163 V88 V163 1.3030145350444111e-19

R88_164 V88 V164 -415.12067689020057
L88_164 V88 V164 -2.3323148644920853e-12
C88_164 V88 V164 -3.068596526770382e-19

R88_165 V88 V165 248.80172507005486
L88_165 V88 V165 2.1456617985345664e-11
C88_165 V88 V165 -4.810875499925383e-20

R88_166 V88 V166 -867.0223642838985
L88_166 V88 V166 5.092987897981184e-12
C88_166 V88 V166 1.7432352690470394e-19

R88_167 V88 V167 -634.0208935605623
L88_167 V88 V167 -2.3064238544981552e-12
C88_167 V88 V167 -1.5931069961371086e-19

R88_168 V88 V168 -267.8648436073095
L88_168 V88 V168 -1.932443623839166e-12
C88_168 V88 V168 -7.651276890484256e-20

R88_169 V88 V169 -214.63296895201293
L88_169 V88 V169 2.1901381539760928e-12
C88_169 V88 V169 4.61516097286541e-19

R88_170 V88 V170 -365.28979979550894
L88_170 V88 V170 -3.639228000918999e-12
C88_170 V88 V170 -1.2194669369570696e-19

R88_171 V88 V171 -389.0719044039312
L88_171 V88 V171 -1.5333303852781344e-12
C88_171 V88 V171 -9.662263159691092e-20

R88_172 V88 V172 -465.98934861431894
L88_172 V88 V172 1.0007279061829785e-12
C88_172 V88 V172 1.479231130138799e-19

R88_173 V88 V173 -713.1648660498287
L88_173 V88 V173 -2.426803584559379e-12
C88_173 V88 V173 -1.3858559593959092e-19

R88_174 V88 V174 670.4163704623703
L88_174 V88 V174 2.4225792194964502e-12
C88_174 V88 V174 2.1439993321598038e-19

R88_175 V88 V175 1307.698432836339
L88_175 V88 V175 1.4917408660978584e-12
C88_175 V88 V175 1.2409186980437685e-19

R88_176 V88 V176 221.9415872644666
L88_176 V88 V176 -9.561675907946258e-13
C88_176 V88 V176 -5.596644428122244e-19

R88_177 V88 V177 442.67837601809237
L88_177 V88 V177 2.424281769203754e-12
C88_177 V88 V177 -4.0718486235129195e-20

R88_178 V88 V178 978.3692107101591
L88_178 V88 V178 4.158663589741984e-12
C88_178 V88 V178 4.976296346407875e-20

R88_179 V88 V179 5452.4404425410685
L88_179 V88 V179 2.1533316332882183e-12
C88_179 V88 V179 1.785740299440318e-19

R88_180 V88 V180 143.6415880775055
L88_180 V88 V180 1.4245895430974278e-12
C88_180 V88 V180 5.688758292203912e-19

R88_181 V88 V181 -998.782275077421
L88_181 V88 V181 -5.985572635792803e-12
C88_181 V88 V181 -7.943505974867413e-20

R88_182 V88 V182 -479.3422633348778
L88_182 V88 V182 -1.9686549928920683e-12
C88_182 V88 V182 -1.2222199938351732e-19

R88_183 V88 V183 1024.058993835027
L88_183 V88 V183 2.6916883458366817e-12
C88_183 V88 V183 1.319317535187221e-19

R88_184 V88 V184 -134.96132146710946
L88_184 V88 V184 1.25142550452606e-12
C88_184 V88 V184 -6.064426878153676e-20

R88_185 V88 V185 -461.300610358117
L88_185 V88 V185 -1.6969534358492505e-12
C88_185 V88 V185 4.025043229732906e-20

R88_186 V88 V186 188876.32953043864
L88_186 V88 V186 2.268632313640571e-12
C88_186 V88 V186 -5.427623909708762e-20

R88_187 V88 V187 624.3216662203507
L88_187 V88 V187 -8.236570580987108e-12
C88_187 V88 V187 -2.209555647446988e-19

R88_188 V88 V188 -561.4953011368148
L88_188 V88 V188 -3.737789359358378e-13
C88_188 V88 V188 -5.209818396006475e-19

R88_189 V88 V189 862.1593320426841
L88_189 V88 V189 1.5487219628925824e-12
C88_189 V88 V189 1.1363431165695568e-19

R88_190 V88 V190 1979.1238232570354
L88_190 V88 V190 7.06247808689016e-12
C88_190 V88 V190 1.1756780903812007e-19

R88_191 V88 V191 -545.0354555222091
L88_191 V88 V191 -7.793306871315947e-13
C88_191 V88 V191 -2.0583162937256722e-19

R88_192 V88 V192 133.04914312490502
L88_192 V88 V192 7.994864983434689e-13
C88_192 V88 V192 5.868811112534386e-19

R88_193 V88 V193 369.6022471309556
L88_193 V88 V193 2.5717615296925985e-12
C88_193 V88 V193 1.4239252692637391e-19

R88_194 V88 V194 -765.2282524455787
L88_194 V88 V194 1.840915269055406e-12
C88_194 V88 V194 4.778006567500372e-19

R88_195 V88 V195 -8266.763631429456
L88_195 V88 V195 6.294523005119308e-13
C88_195 V88 V195 6.476498314383718e-19

R88_196 V88 V196 -182.3316316922655
L88_196 V88 V196 -1.3615796274245723e-12
C88_196 V88 V196 -8.519216056575769e-19

R88_197 V88 V197 -877.9995201280458
L88_197 V88 V197 -2.9934400299394895e-12
C88_197 V88 V197 -2.125267198140162e-19

R88_198 V88 V198 -457.20923585843593
L88_198 V88 V198 -1.1352119501699715e-10
C88_198 V88 V198 8.788447975703321e-20

R88_199 V88 V199 -365.25139817169253
L88_199 V88 V199 5.831224296901411e-12
C88_199 V88 V199 -2.2341125758318703e-20

R88_200 V88 V200 -629.5761868219705
L88_200 V88 V200 -4.164352058610411e-11
C88_200 V88 V200 7.650506777055223e-20

R89_89 V89 0 317.6328166739836
L89_89 V89 0 -9.266783248276995e-13
C89_89 V89 0 -1.677468730139108e-18

R89_90 V89 V90 332.8273674496935
L89_90 V89 V90 -7.752220748714793e-13
C89_90 V89 V90 -6.789240036468746e-19

R89_91 V89 V91 289.8112174904199
L89_91 V89 V91 1.8126914838887313e-12
C89_91 V89 V91 2.74462181311503e-19

R89_92 V89 V92 284.45732230575373
L89_92 V89 V92 1.3027439739359966e-12
C89_92 V89 V92 2.308199487970189e-19

R89_93 V89 V93 165.23271560303573
L89_93 V89 V93 2.1985035879053e-12
C89_93 V89 V93 1.6076389033823373e-19

R89_94 V89 V94 935.204281051269
L89_94 V89 V94 1.7142846293208956e-12
C89_94 V89 V94 3.1693900090190505e-19

R89_95 V89 V95 2974.116831553609
L89_95 V89 V95 2.634282384119572e-12
C89_95 V89 V95 2.5070634024450655e-19

R89_96 V89 V96 1090.398613396336
L89_96 V89 V96 2.5920666541401807e-12
C89_96 V89 V96 3.3202500782305234e-19

R89_97 V89 V97 -656.1371546093186
L89_97 V89 V97 6.232571421601728e-13
C89_97 V89 V97 9.018801586050224e-19

R89_98 V89 V98 -312.15712819047184
L89_98 V89 V98 1.62866774169797e-12
C89_98 V89 V98 3.9358190600760216e-19

R89_99 V89 V99 -270.7828515946549
L89_99 V89 V99 -9.651768367416086e-13
C89_99 V89 V99 -5.541662979514171e-19

R89_100 V89 V100 -270.6118316810459
L89_100 V89 V100 -1.6474327108012753e-12
C89_100 V89 V100 -4.53919842696179e-19

R89_101 V89 V101 -271.28920011509246
L89_101 V89 V101 -1.0731638629339645e-12
C89_101 V89 V101 -5.608332077186504e-19

R89_102 V89 V102 4223.199380542713
L89_102 V89 V102 -2.230492626933827e-12
C89_102 V89 V102 -3.0315419516529336e-19

R89_103 V89 V103 1460.9772448301444
L89_103 V89 V103 6.00302113432509e-12
C89_103 V89 V103 3.679344396359343e-20

R89_104 V89 V104 2450.0945496849786
L89_104 V89 V104 4.129793720273101e-12
C89_104 V89 V104 3.185587871036619e-20

R89_105 V89 V105 155.2302910659798
L89_105 V89 V105 -1.2190166435824758e-12
C89_105 V89 V105 -2.733724896934268e-19

R89_106 V89 V106 1496.9572827056386
L89_106 V89 V106 -1.8751365615107353e-12
C89_106 V89 V106 -3.2331787283202355e-19

R89_107 V89 V107 718.4498845593463
L89_107 V89 V107 1.4864937027051058e-12
C89_107 V89 V107 3.5384786183888273e-19

R89_108 V89 V108 583.3982904755368
L89_108 V89 V108 -5.105706353198098e-12
C89_108 V89 V108 4.0288435762587266e-20

R89_109 V89 V109 -790.759313025198
L89_109 V89 V109 2.7791418995848285e-12
C89_109 V89 V109 4.0520679075848363e-19

R89_110 V89 V110 -3979.6658181373928
L89_110 V89 V110 2.596533535910745e-12
C89_110 V89 V110 2.8791893773518573e-19

R89_111 V89 V111 -1154.6498567523377
L89_111 V89 V111 -1.2309277638749496e-11
C89_111 V89 V111 -2.249593147218299e-20

R89_112 V89 V112 -963.0366269100253
L89_112 V89 V112 2.249026756171225e-12
C89_112 V89 V112 2.0260127128829226e-19

R89_113 V89 V113 -303.3419415401451
L89_113 V89 V113 1.9338456298018777e-12
C89_113 V89 V113 1.3697777033954898e-19

R89_114 V89 V114 -93615.9457172946
L89_114 V89 V114 1.5163608832294904e-12
C89_114 V89 V114 3.261476219200917e-19

R89_115 V89 V115 -2485.7392022216836
L89_115 V89 V115 -1.6663283900311718e-12
C89_115 V89 V115 -2.2491069191950553e-19

R89_116 V89 V116 -896.5596585899142
L89_116 V89 V116 -3.6278530767894218e-12
C89_116 V89 V116 -6.751653500320506e-20

R89_117 V89 V117 279.37567796238096
L89_117 V89 V117 -1.1304034791862498e-11
C89_117 V89 V117 -4.432796433179289e-20

R89_118 V89 V118 -2642.7216583772133
L89_118 V89 V118 -1.1525205242411023e-12
C89_118 V89 V118 -4.668657121952653e-19

R89_119 V89 V119 3623.8645574179777
L89_119 V89 V119 -1.2204568653604631e-11
C89_119 V89 V119 -1.4809512937661696e-19

R89_120 V89 V120 935.2339563810348
L89_120 V89 V120 -2.333276453956434e-12
C89_120 V89 V120 -3.7081787931860513e-19

R89_121 V89 V121 3245.125916261187
L89_121 V89 V121 -2.44749841097231e-12
C89_121 V89 V121 -1.5939687603030974e-19

R89_122 V89 V122 148419.64781235022
L89_122 V89 V122 3.644314705317089e-12
C89_122 V89 V122 1.0198278318677819e-19

R89_123 V89 V123 -27771.21731458264
L89_123 V89 V123 1.4188611297528331e-12
C89_123 V89 V123 3.26701975201425e-19

R89_124 V89 V124 -15933.376870101138
L89_124 V89 V124 8.853856466255688e-13
C89_124 V89 V124 5.534588426133537e-19

R89_125 V89 V125 -1728.079739602195
L89_125 V89 V125 -2.163787598992861e-12
C89_125 V89 V125 -1.8172778719541038e-19

R89_126 V89 V126 1476.5089898262347
L89_126 V89 V126 1.6280803410014701e-12
C89_126 V89 V126 1.8795942438311984e-19

R89_127 V89 V127 2983.807339478957
L89_127 V89 V127 2.5207210024403422e-11
C89_127 V89 V127 4.687061175522847e-20

R89_128 V89 V128 -3033.7596389102114
L89_128 V89 V128 -2.4968539571243455e-12
C89_128 V89 V128 -3.839638800499959e-20

R89_129 V89 V129 894.8783323065007
L89_129 V89 V129 1.2595742575853887e-12
C89_129 V89 V129 5.77614430641774e-19

R89_130 V89 V130 -2021.767365530667
L89_130 V89 V130 -1.7142982547432702e-12
C89_130 V89 V130 -2.0082616756882275e-19

R89_131 V89 V131 -1484.670656096421
L89_131 V89 V131 -2.0366292936487586e-12
C89_131 V89 V131 -2.2480906964681326e-19

R89_132 V89 V132 -1895.622350682826
L89_132 V89 V132 -1.6599428641787717e-12
C89_132 V89 V132 -3.6264181578997214e-19

R89_133 V89 V133 -914.7113401658617
L89_133 V89 V133 -2.8201441676395204e-12
C89_133 V89 V133 -4.2360830096354697e-19

R89_134 V89 V134 4578.112815527597
L89_134 V89 V134 3.0762984671136363e-12
C89_134 V89 V134 8.569652359252805e-20

R89_135 V89 V135 3894.520953679966
L89_135 V89 V135 6.339297203406015e-12
C89_135 V89 V135 1.0761228918438427e-19

R89_136 V89 V136 -131570.43679865883
L89_136 V89 V136 1.5395231630022738e-12
C89_136 V89 V136 3.989752041087975e-19

R89_137 V89 V137 1080.2674719833433
L89_137 V89 V137 -8.427406780596274e-12
C89_137 V89 V137 -7.573193544060739e-20

R89_138 V89 V138 1885.9245020393923
L89_138 V89 V138 5.175060945134142e-12
C89_138 V89 V138 6.751700865588106e-20

R89_139 V89 V139 15243.66802501483
L89_139 V89 V139 -3.912749750954155e-12
C89_139 V89 V139 -2.231368450335295e-19

R89_140 V89 V140 1492.8524314293045
L89_140 V89 V140 -5.337575306125063e-12
C89_140 V89 V140 -3.509361203722208e-19

R89_141 V89 V141 -5680.618979730411
L89_141 V89 V141 1.4186757232698695e-12
C89_141 V89 V141 4.843283631220815e-19

R89_142 V89 V142 -773.946393544508
L89_142 V89 V142 -2.975573552250724e-12
C89_142 V89 V142 -6.552934462877059e-20

R89_143 V89 V143 -2405.6255453613007
L89_143 V89 V143 1.6162928827782746e-12
C89_143 V89 V143 2.139894434068713e-19

R89_144 V89 V144 -2813.71005106719
L89_144 V89 V144 -1.9966090114922715e-11
C89_144 V89 V144 4.4034169910271305e-20

R89_145 V89 V145 921.3495671164133
L89_145 V89 V145 -4.313627640404402e-12
C89_145 V89 V145 -3.3090561147769896e-20

R89_146 V89 V146 9648.447200969918
L89_146 V89 V146 8.075884043591627e-12
C89_146 V89 V146 -4.269962043543671e-20

R89_147 V89 V147 2160.0834002181155
L89_147 V89 V147 -4.889183200965817e-11
C89_147 V89 V147 1.932754881200891e-19

R89_148 V89 V148 11487.804644060536
L89_148 V89 V148 1.7819386113255247e-12
C89_148 V89 V148 2.492447503269477e-19

R89_149 V89 V149 -378.3255674462749
L89_149 V89 V149 -6.291284210451066e-13
C89_149 V89 V149 -7.12673891372435e-19

R89_150 V89 V150 1092.3413392500913
L89_150 V89 V150 -1.1421406106699179e-11
C89_150 V89 V150 3.3991397636864113e-19

R89_151 V89 V151 -2680.656414350645
L89_151 V89 V151 -1.7467119519593817e-12
C89_151 V89 V151 -2.4390823660047764e-19

R89_152 V89 V152 -1085.4579346019932
L89_152 V89 V152 -2.272733637276941e-12
C89_152 V89 V152 -4.5830701880970795e-20

R89_153 V89 V153 502.20149130008775
L89_153 V89 V153 3.5287839125865374e-12
C89_153 V89 V153 1.737931501179165e-19

R89_154 V89 V154 -2309.115714472989
L89_154 V89 V154 3.055984652189853e-11
C89_154 V89 V154 -1.9267986111773176e-19

R89_155 V89 V155 6166.317204443375
L89_155 V89 V155 -1.7491694372520064e-12
C89_155 V89 V155 -2.0764014776854043e-19

R89_156 V89 V156 2377.9860268658454
L89_156 V89 V156 1.526523548002614e-11
C89_156 V89 V156 -2.3572303208572677e-19

R89_157 V89 V157 722.2840733256809
L89_157 V89 V157 5.722796100875073e-13
C89_157 V89 V157 7.399371283121684e-19

R89_158 V89 V158 -1391.4790834765754
L89_158 V89 V158 -1.0057557000886858e-11
C89_158 V89 V158 -5.632312747501391e-20

R89_159 V89 V159 -7402.5299226403795
L89_159 V89 V159 1.5087057559681539e-12
C89_159 V89 V159 1.6068918518616263e-19

R89_160 V89 V160 1569.5867906720032
L89_160 V89 V160 2.895763608658187e-12
C89_160 V89 V160 1.0369912341583348e-19

R89_161 V89 V161 1030.376015769118
L89_161 V89 V161 -1.9791197390226263e-12
C89_161 V89 V161 -1.6914170623190606e-19

R89_162 V89 V162 -2202.931958475615
L89_162 V89 V162 -2.1374290285038526e-12
C89_162 V89 V162 -5.684401253434752e-20

R89_163 V89 V163 -1307.8383794859346
L89_163 V89 V163 2.3641147621741486e-12
C89_163 V89 V163 1.399261587948633e-19

R89_164 V89 V164 -1721.4084691403555
L89_164 V89 V164 1.219369470820043e-11
C89_164 V89 V164 -8.666168581934624e-20

R89_165 V89 V165 -6963.426466113696
L89_165 V89 V165 -7.888486089421561e-13
C89_165 V89 V165 -4.0088401074926327e-19

R89_166 V89 V166 -2189.968335338118
L89_166 V89 V166 -1.0816497742095404e-11
C89_166 V89 V166 8.231906194734948e-20

R89_167 V89 V167 -4331.907089691795
L89_167 V89 V167 -3.3927550255969515e-12
C89_167 V89 V167 -1.0151868290463705e-19

R89_168 V89 V168 -977.9783637201186
L89_168 V89 V168 -1.6195129115739946e-12
C89_168 V89 V168 -2.0133818592459767e-20

R89_169 V89 V169 2221.890588824426
L89_169 V89 V169 1.1403068812023168e-12
C89_169 V89 V169 3.877644502675722e-19

R89_170 V89 V170 1313.2817917239222
L89_170 V89 V170 -3.93570983134283e-12
C89_170 V89 V170 -2.2884543642173245e-19

R89_171 V89 V171 1046.0766618026762
L89_171 V89 V171 -1.0698645213534955e-12
C89_171 V89 V171 -2.565902309031198e-19

R89_172 V89 V172 1965.1862305542872
L89_172 V89 V172 7.099208411635466e-12
C89_172 V89 V172 -7.09175751700122e-20

R89_173 V89 V173 718.9377987902434
L89_173 V89 V173 2.8797342535214104e-12
C89_173 V89 V173 9.882971999043889e-21

R89_174 V89 V174 -2665.1779948174276
L89_174 V89 V174 1.3656983943065437e-12
C89_174 V89 V174 3.225842869232918e-19

R89_175 V89 V175 -1669.3159063391122
L89_175 V89 V175 2.8334579176831e-12
C89_175 V89 V175 -4.888496934964135e-20

R89_176 V89 V176 5447.695575132381
L89_176 V89 V176 6.632100533063447e-12
C89_176 V89 V176 -1.2696579025203485e-19

R89_177 V89 V177 -1184.690141989487
L89_177 V89 V177 -1.7322406527442296e-11
C89_177 V89 V177 -5.62538789695527e-20

R89_178 V89 V178 2096.919983584379
L89_178 V89 V178 3.4928783996123684e-12
C89_178 V89 V178 1.055337199023782e-19

R89_179 V89 V179 -2916834.864284411
L89_179 V89 V179 1.470307985481486e-12
C89_179 V89 V179 4.068475872010979e-19

R89_180 V89 V180 1677.0474395282042
L89_180 V89 V180 2.1071536210532943e-12
C89_180 V89 V180 3.715284112586685e-19

R89_181 V89 V181 -5347.004266003057
L89_181 V89 V181 -1.589186344197234e-12
C89_181 V89 V181 -1.6194954925490362e-19

R89_182 V89 V182 -2568.6150753738925
L89_182 V89 V182 -8.75553237796608e-13
C89_182 V89 V182 -2.5395245265802996e-19

R89_183 V89 V183 9423.185217044704
L89_183 V89 V183 2.2700294635786107e-12
C89_183 V89 V183 8.180978120469765e-20

R89_184 V89 V184 -1743.2713849037675
L89_184 V89 V184 4.490226720773873e-12
C89_184 V89 V184 -4.81706928662391e-20

R89_185 V89 V185 715.7855031853128
L89_185 V89 V185 -1.856574704644203e-11
C89_185 V89 V185 1.2675914946611433e-19

R89_186 V89 V186 -718.5959299430275
L89_186 V89 V186 -7.226344631418263e-12
C89_186 V89 V186 -8.612664436158788e-21

R89_187 V89 V187 -2633.08053902168
L89_187 V89 V187 -1.1969659178050721e-12
C89_187 V89 V187 -3.645726859835506e-19

R89_188 V89 V188 -1497.8389425484447
L89_188 V89 V188 -6.580555190058835e-13
C89_188 V89 V188 -3.4023541443041327e-19

R89_189 V89 V189 -820.5125570340865
L89_189 V89 V189 1.0825545401131761e-12
C89_189 V89 V189 -8.306749744852538e-21

R89_190 V89 V190 1239.8383610698565
L89_190 V89 V190 2.085152711613524e-12
C89_190 V89 V190 1.95095978126993e-19

R89_191 V89 V191 982.3201741154244
L89_191 V89 V191 -1.1841627447185221e-12
C89_191 V89 V191 -1.1235323946328513e-19

R89_192 V89 V192 632.7841114379034
L89_192 V89 V192 2.431464048440444e-12
C89_192 V89 V192 1.4392816405895157e-19

R89_193 V89 V193 -827.4824566377259
L89_193 V89 V193 -4.906474699332922e-12
C89_193 V89 V193 9.714232858947099e-20

R89_194 V89 V194 543.753011425981
L89_194 V89 V194 1.0909936934299727e-12
C89_194 V89 V194 2.9490992001654054e-19

R89_195 V89 V195 3469.4963162875915
L89_195 V89 V195 7.069680594254366e-13
C89_195 V89 V195 3.56663611255733e-19

R89_196 V89 V196 4016.9729267147763
L89_196 V89 V196 1.0746044579156829e-12
C89_196 V89 V196 7.528693899377825e-20

R89_197 V89 V197 536.238794040965
L89_197 V89 V197 8.362587938128876e-12
C89_197 V89 V197 -7.239571667014089e-23

R89_198 V89 V198 -528.9432462046502
L89_198 V89 V198 -1.8225822808078938e-12
C89_198 V89 V198 -3.9926087986476484e-20

R89_199 V89 V199 -396.2550422838592
L89_199 V89 V199 5.394069415258463e-12
C89_199 V89 V199 1.2595500056528698e-19

R89_200 V89 V200 -442.57730444490954
L89_200 V89 V200 -3.817433725350245e-12
C89_200 V89 V200 -2.352502970587689e-20

R90_90 V90 0 -80.1337415984462
L90_90 V90 0 -1.8487207506540208e-13
C90_90 V90 0 -2.87197710965494e-18

R90_91 V90 V91 -331.93308530550325
L90_91 V90 V91 6.614429000102931e-13
C90_91 V90 V91 7.708367720890995e-19

R90_92 V90 V92 -772.2124825252715
L90_92 V90 V92 7.724370801075261e-13
C90_92 V90 V92 4.111553540723235e-19

R90_93 V90 V93 -191.11335663738294
L90_93 V90 V93 4.667866315303497e-12
C90_93 V90 V93 2.6450453586343486e-19

R90_94 V90 V94 -20583.37061937688
L90_94 V90 V94 8.690568362913014e-13
C90_94 V90 V94 8.881061253105791e-19

R90_95 V90 V95 964.3298413108408
L90_95 V90 V95 3.79994450170167e-12
C90_95 V90 V95 3.6223100662871106e-19

R90_96 V90 V96 16849.250668300483
L90_96 V90 V96 9.667924270159675e-12
C90_96 V90 V96 4.649587764412225e-19

R90_97 V90 V97 1460.9075014140374
L90_97 V90 V97 6.381484441317346e-13
C90_97 V90 V97 1.0941405219961325e-18

R90_98 V90 V98 117.24500214767974
L90_98 V90 V98 4.555838983396567e-13
C90_98 V90 V98 1.142080931717986e-18

R90_99 V90 V99 2437.110288067903
L90_99 V90 V99 -4.5311694378221324e-13
C90_99 V90 V99 -1.2387836782985029e-18

R90_100 V90 V100 -1119.1382969259357
L90_100 V90 V100 -9.428663423612121e-13
C90_100 V90 V100 -7.963207895701316e-19

R90_101 V90 V101 627.5094497180778
L90_101 V90 V101 -8.347756937313848e-13
C90_101 V90 V101 -8.528879932190105e-19

R90_102 V90 V102 -170.85603173309536
L90_102 V90 V102 -6.109755051977344e-13
C90_102 V90 V102 -1.0880193114520413e-18

R90_103 V90 V103 533.7265922999196
L90_103 V90 V103 1.242458626799732e-12
C90_103 V90 V103 2.674320594583911e-19

R90_104 V90 V104 313.0474597954351
L90_104 V90 V104 1.1256420010119345e-12
C90_104 V90 V104 2.2573549396156254e-19

R90_105 V90 V105 -479.1356488232244
L90_105 V90 V105 -2.144324041822295e-12
C90_105 V90 V105 -2.7110268053109653e-19

R90_106 V90 V106 144.19829477566017
L90_106 V90 V106 -1.085374090463383e-12
C90_106 V90 V106 -3.9571724682779703e-19

R90_107 V90 V107 -693.8067812782167
L90_107 V90 V107 9.842251464525596e-13
C90_107 V90 V107 6.822969224572902e-19

R90_108 V90 V108 -2032.1019696159824
L90_108 V90 V108 -2.3548303348490814e-12
C90_108 V90 V108 8.001890063567677e-21

R90_109 V90 V109 -717.1710906363793
L90_109 V90 V109 1.2740730403487831e-12
C90_109 V90 V109 7.9926977633744385e-19

R90_110 V90 V110 -173.72155957951077
L90_110 V90 V110 9.890036457066598e-13
C90_110 V90 V110 5.861011352959925e-19

R90_111 V90 V111 -689.7801683663245
L90_111 V90 V111 -6.50133318934619e-12
C90_111 V90 V111 -8.677877786476487e-20

R90_112 V90 V112 -446.43040119348825
L90_112 V90 V112 2.0982177856684313e-12
C90_112 V90 V112 2.1028627022479629e-19

R90_113 V90 V113 -479.5221807865637
L90_113 V90 V113 3.8923897489352566e-12
C90_113 V90 V113 7.428172747613431e-20

R90_114 V90 V114 -169.92825284115557
L90_114 V90 V114 1.0345142017712968e-12
C90_114 V90 V114 6.096763612036065e-19

R90_115 V90 V115 525.8048484499557
L90_115 V90 V115 -8.738228209363033e-13
C90_115 V90 V115 -4.649119379068783e-19

R90_116 V90 V116 891.3646076677702
L90_116 V90 V116 -2.5372995398492994e-12
C90_116 V90 V116 -7.040969571125597e-21

R90_117 V90 V117 712.8393357899239
L90_117 V90 V117 -1.6710637639972124e-12
C90_117 V90 V117 -3.656969366491496e-19

R90_118 V90 V118 54.58626423351456
L90_118 V90 V118 -6.796297646039185e-13
C90_118 V90 V118 -1.0990082552699511e-18

R90_119 V90 V119 380.0726906941185
L90_119 V90 V119 -2.760304850896168e-11
C90_119 V90 V119 -2.1147356622313022e-19

R90_120 V90 V120 452.94286210470966
L90_120 V90 V120 -1.4647910408118012e-12
C90_120 V90 V120 -6.507599825792661e-19

R90_121 V90 V121 1170.6233843784164
L90_121 V90 V121 -6.605145311546454e-11
C90_121 V90 V121 7.30212902262303e-20

R90_122 V90 V122 -163.6164761386148
L90_122 V90 V122 2.3270354919140918e-12
C90_122 V90 V122 2.991030683259609e-19

R90_123 V90 V123 -651.6012339368638
L90_123 V90 V123 8.367285888894576e-13
C90_123 V90 V123 6.321617915814471e-19

R90_124 V90 V124 -632.8546780379049
L90_124 V90 V124 6.117935290994763e-13
C90_124 V90 V124 8.600798768454419e-19

R90_125 V90 V125 -548.4408343537386
L90_125 V90 V125 -5.228431462578957e-11
C90_125 V90 V125 -1.4259738424642004e-19

R90_126 V90 V126 -59.61656524981727
L90_126 V90 V126 7.781033672582387e-13
C90_126 V90 V126 7.883098502717135e-19

R90_127 V90 V127 -180.9706221857905
L90_127 V90 V127 -6.417104521692288e-12
C90_127 V90 V127 -2.7317650426017594e-21

R90_128 V90 V128 -215.49088597740885
L90_128 V90 V128 -2.45724769036205e-12
C90_128 V90 V128 6.995573074518803e-20

R90_129 V90 V129 -331.35848320414897
L90_129 V90 V129 1.6390100008483203e-12
C90_129 V90 V129 7.033519016315821e-19

R90_130 V90 V130 72.0927126763651
L90_130 V90 V130 -9.530449220140676e-13
C90_130 V90 V130 -8.336805618329581e-19

R90_131 V90 V131 121.70089540677355
L90_131 V90 V131 -2.0195672754620758e-12
C90_131 V90 V131 -3.7991306101642624e-19

R90_132 V90 V132 96.35613186054033
L90_132 V90 V132 -1.0899316847109893e-12
C90_132 V90 V132 -7.509806171220169e-19

R90_133 V90 V133 312.71038843435497
L90_133 V90 V133 -1.962177841255509e-12
C90_133 V90 V133 -5.140857330315958e-19

R90_134 V90 V134 218.37228309654964
L90_134 V90 V134 8.81771211798313e-12
C90_134 V90 V134 2.2923868791803387e-19

R90_135 V90 V135 1135.150029250627
L90_135 V90 V135 2.4872381548971075e-12
C90_135 V90 V135 4.2040851839863774e-19

R90_136 V90 V136 326.1787430871825
L90_136 V90 V136 1.0668363397160252e-12
C90_136 V90 V136 6.995593481038883e-19

R90_137 V90 V137 -1210.0778942176742
L90_137 V90 V137 -1.7575458947233496e-12
C90_137 V90 V137 -3.782821669242517e-19

R90_138 V90 V138 -87.7509692763465
L90_138 V90 V138 1.1560962110133403e-12
C90_138 V90 V138 3.4801851664532296e-19

R90_139 V90 V139 -122.80430916576401
L90_139 V90 V139 -1.0275309641585687e-12
C90_139 V90 V139 -7.212907630651017e-19

R90_140 V90 V140 -72.49531257447664
L90_140 V90 V140 -1.2915895888659615e-12
C90_140 V90 V140 -6.996982851226148e-19

R90_141 V90 V141 342.2049387980257
L90_141 V90 V141 6.976759833783359e-13
C90_141 V90 V141 9.615637153004146e-19

R90_142 V90 V142 -680.1567130042955
L90_142 V90 V142 -5.580065462144015e-12
C90_142 V90 V142 -2.115053464587389e-19

R90_143 V90 V143 157.4619279806081
L90_143 V90 V143 8.855734958440073e-13
C90_143 V90 V143 4.539103170178337e-19

R90_144 V90 V144 132.49482247250634
L90_144 V90 V144 3.4150443217137637e-12
C90_144 V90 V144 1.9009739530117404e-19

R90_145 V90 V145 -2831.453317994964
L90_145 V90 V145 1.4255213255953577e-12
C90_145 V90 V145 3.5488073843277356e-19

R90_146 V90 V146 68.64708095718609
L90_146 V90 V146 -2.7679750914001163e-12
C90_146 V90 V146 -1.7150223732315184e-19

R90_147 V90 V147 945.8116253037243
L90_147 V90 V147 1.9698614892316888e-12
C90_147 V90 V147 6.102852781025293e-19

R90_148 V90 V148 884.1285388321454
L90_148 V90 V148 7.370437317600176e-13
C90_148 V90 V148 5.379001288903178e-19

R90_149 V90 V149 -385.5882802038583
L90_149 V90 V149 -3.1523724251922694e-13
C90_149 V90 V149 -1.619260920639679e-18

R90_150 V90 V150 418.64497333220964
L90_150 V90 V150 -2.83872521039065e-11
C90_150 V90 V150 7.973059016785784e-19

R90_151 V90 V151 -149.3005901255492
L90_151 V90 V151 -1.3500621463604734e-12
C90_151 V90 V151 -4.525213119969777e-19

R90_152 V90 V152 -113.3980913380414
L90_152 V90 V152 -1.206705887938452e-12
C90_152 V90 V152 -1.243145701060788e-19

R90_153 V90 V153 -398.9927010124389
L90_153 V90 V153 -2.6563388743268952e-12
C90_153 V90 V153 -2.3255012302782266e-20

R90_154 V90 V154 -89.33906720797873
L90_154 V90 V154 3.254896174154051e-12
C90_154 V90 V154 -4.122974837144496e-19

R90_155 V90 V155 362.3740392531419
L90_155 V90 V155 -6.690274717459128e-13
C90_155 V90 V155 -5.989143355490576e-19

R90_156 V90 V156 178.06883382632537
L90_156 V90 V156 -3.2063347320163746e-12
C90_156 V90 V156 -5.088401800792496e-19

R90_157 V90 V157 313.6890350806923
L90_157 V90 V157 3.22766732004292e-13
C90_157 V90 V157 1.5422917186734545e-18

R90_158 V90 V158 213.82633891216858
L90_158 V90 V158 -2.280539418829608e-12
C90_158 V90 V158 -2.151633129295035e-19

R90_159 V90 V159 137.01557883182264
L90_159 V90 V159 1.0049222942797888e-12
C90_159 V90 V159 2.9575002344565527e-19

R90_160 V90 V160 105.75624634149128
L90_160 V90 V160 3.6284870988636335e-12
C90_160 V90 V160 1.1645052973657695e-19

R90_161 V90 V161 -141.06111925166135
L90_161 V90 V161 -2.652032101053482e-12
C90_161 V90 V161 -1.0662833287955424e-19

R90_162 V90 V162 1607.6818698575241
L90_162 V90 V162 -8.700480264349426e-13
C90_162 V90 V162 -1.158004033722341e-19

R90_163 V90 V163 -122.71529833104096
L90_163 V90 V163 2.115782966190658e-12
C90_163 V90 V163 1.7011621177119878e-19

R90_164 V90 V164 -78.75831706904881
L90_164 V90 V164 2.327871887766069e-12
C90_164 V90 V164 -1.0287801006689023e-19

R90_165 V90 V165 -25430.28563515631
L90_165 V90 V165 -6.906005433174427e-13
C90_165 V90 V165 -7.135948415658676e-19

R90_166 V90 V166 -364.0484327064992
L90_166 V90 V166 1.80405036433839e-12
C90_166 V90 V166 3.435773531155801e-19

R90_167 V90 V167 -4080.877585043291
L90_167 V90 V167 -2.752156508962936e-12
C90_167 V90 V167 -7.694098632577415e-20

R90_168 V90 V168 825.3876267432436
L90_168 V90 V168 -1.159528342653994e-12
C90_168 V90 V168 1.107397023402229e-19

R90_169 V90 V169 111.06064869298582
L90_169 V90 V169 1.5445194339487236e-12
C90_169 V90 V169 4.327758894542263e-19

R90_170 V90 V170 142.48982622917694
L90_170 V90 V170 5.796648107282514e-11
C90_170 V90 V170 -5.185793328166015e-19

R90_171 V90 V171 143.25172755684164
L90_171 V90 V171 -1.0563379032841897e-12
C90_171 V90 V171 -4.0112913566665703e-19

R90_172 V90 V172 131.1741346841227
L90_172 V90 V172 2.591451030130797e-12
C90_172 V90 V172 -1.894130536464526e-19

R90_173 V90 V173 -156.0124665209511
L90_173 V90 V173 4.047615995607799e-12
C90_173 V90 V173 4.569999199954346e-20

R90_174 V90 V174 5190.732796223534
L90_174 V90 V174 5.938967223087402e-12
C90_174 V90 V174 4.466088972173692e-19

R90_175 V90 V175 -603.9791531729193
L90_175 V90 V175 -8.693565838547314e-12
C90_175 V90 V175 -2.5830819873548515e-19

R90_176 V90 V176 -229.74464935076122
L90_176 V90 V176 -2.8704315985280406e-12
C90_176 V90 V176 -3.185443593954906e-19

R90_177 V90 V177 -251.86794965001218
L90_177 V90 V177 1.0674163351241803e-11
C90_177 V90 V177 -6.322209180226367e-20

R90_178 V90 V178 -111.18088813180013
L90_178 V90 V178 -1.8192691447500937e-11
C90_178 V90 V178 2.513848993747985e-19

R90_179 V90 V179 -529.557561184516
L90_179 V90 V179 9.53826121122896e-13
C90_179 V90 V179 7.554714190538391e-19

R90_180 V90 V180 -536.1473172911886
L90_180 V90 V180 1.2876793588100447e-12
C90_180 V90 V180 6.729740813153547e-19

R90_181 V90 V181 154.78481366108718
L90_181 V90 V181 -1.113367599900317e-11
C90_181 V90 V181 1.4240194277474854e-20

R90_182 V90 V182 105.85870588670406
L90_182 V90 V182 -1.1968046771957955e-12
C90_182 V90 V182 -4.236992435529593e-19

R90_183 V90 V183 788.1109785159596
L90_183 V90 V183 1.1392778245438924e-12
C90_183 V90 V183 1.062574300817026e-19

R90_184 V90 V184 481.23330801527317
L90_184 V90 V184 1.5977459615470795e-12
C90_184 V90 V184 -7.979401248924161e-20

R90_185 V90 V185 -1755.4721877440797
L90_185 V90 V185 -2.7279697909996017e-12
C90_185 V90 V185 -2.944001660362122e-20

R90_186 V90 V186 169.35655451992994
L90_186 V90 V186 1.3109463432996657e-12
C90_186 V90 V186 5.69919330507528e-20

R90_187 V90 V187 -1266.1548569569195
L90_187 V90 V187 -7.468816443972221e-13
C90_187 V90 V187 -6.7765151780575375e-19

R90_188 V90 V188 -310.3925295769016
L90_188 V90 V188 -4.601571814895541e-13
C90_188 V90 V188 -5.255639230610393e-19

R90_189 V90 V189 -452.0613140793566
L90_189 V90 V189 2.1159468619134693e-10
C90_189 V90 V189 -8.797880911687583e-20

R90_190 V90 V190 -157.85200147532467
L90_190 V90 V190 -2.1107062615029164e-12
C90_190 V90 V190 3.4747083823987794e-19

R90_191 V90 V191 -368.7101814250391
L90_191 V90 V191 -6.734513201430233e-13
C90_191 V90 V191 -6.464555516164722e-20

R90_192 V90 V192 -615.6807131971221
L90_192 V90 V192 7.833162105672965e-12
C90_192 V90 V192 1.8487453017832773e-19

R90_193 V90 V193 -2856.6695236947094
L90_193 V90 V193 2.2177081289103344e-12
C90_193 V90 V193 2.0779623548003726e-19

R90_194 V90 V194 351.95653134095545
L90_194 V90 V194 1.2392391677595298e-12
C90_194 V90 V194 4.107124181076052e-19

R90_195 V90 V195 427.6436046773238
L90_195 V90 V195 5.218506441259222e-13
C90_195 V90 V195 4.2342665574628577e-19

R90_196 V90 V196 740.6699797590292
L90_196 V90 V196 1.0656833853182135e-12
C90_196 V90 V196 1.0497311583475742e-19

R90_197 V90 V197 2440.5418841125384
L90_197 V90 V197 2.5344753560803398e-12
C90_197 V90 V197 8.314659556632794e-20

R90_198 V90 V198 211.62444216174654
L90_198 V90 V198 2.9712997445605063e-12
C90_198 V90 V198 -1.042821610690248e-19

R90_199 V90 V199 499.3037206994327
L90_199 V90 V199 1.743605768052827e-12
C90_199 V90 V199 1.165206750419472e-19

R90_200 V90 V200 2988.823077804585
L90_200 V90 V200 3.419960929453e-12
C90_200 V90 V200 -2.4075940947974088e-20

R91_91 V91 0 -202.9572361755966
L91_91 V91 0 3.3710757347825983e-13
C91_91 V91 0 1.6245833586586532e-18

R91_92 V91 V92 -450.7766862443444
L91_92 V91 V92 -3.1256632525534703e-12
C91_92 V91 V92 -9.437203925926359e-20

R91_93 V91 V93 -295.49721303167513
L91_93 V91 V93 1.8770004667691644e-12
C91_93 V91 V93 3.2218451352069946e-19

R91_94 V91 V94 -514.6996263669998
L91_94 V91 V94 -1.5415734776324757e-11
C91_94 V91 V94 -6.749735205466221e-20

R91_95 V91 V95 -257.59250575002295
L91_95 V91 V95 8.445210611752975e-12
C91_95 V91 V95 -1.0109248923218164e-19

R91_96 V91 V96 -1081.2252599906333
L91_96 V91 V96 1.243614889716265e-11
C91_96 V91 V96 -5.388773572768724e-20

R91_97 V91 V97 -1392.5394078312222
L91_97 V91 V97 -8.86243526323443e-13
C91_97 V91 V97 -7.263068909706484e-19

R91_98 V91 V98 307.8324405761729
L91_98 V91 V98 -7.705445760885279e-13
C91_98 V91 V98 -6.591364403347174e-19

R91_99 V91 V99 50.93867173420827
L91_99 V91 V99 2.3305856938784965e-13
C91_99 V91 V99 1.9501065214655574e-18

R91_100 V91 V100 591.9318782063777
L91_100 V91 V100 3.1812573702984187e-12
C91_100 V91 V100 2.3960784776464814e-19

R91_101 V91 V101 -4580.25307090777
L91_101 V91 V101 5.016691236022132e-12
C91_101 V91 V101 1.1053528700037188e-19

R91_102 V91 V102 1265.3950163081106
L91_102 V91 V102 1.7756189369496588e-12
C91_102 V91 V102 2.692720235161988e-19

R91_103 V91 V103 -151.22705329979817
L91_103 V91 V103 -4.2000783530896543e-13
C91_103 V91 V103 -9.732947542408254e-19

R91_104 V91 V104 760.7975139239858
L91_104 V91 V104 -2.3510131235459404e-12
C91_104 V91 V104 -2.1990377619066193e-19

R91_105 V91 V105 1500.5243668058824
L91_105 V91 V105 1.5188567554211513e-12
C91_105 V91 V105 3.7619897465390603e-19

R91_106 V91 V106 950.7994983965309
L91_106 V91 V106 7.343655339015857e-13
C91_106 V91 V106 7.385883052619611e-19

R91_107 V91 V107 -93.90122792154179
L91_107 V91 V107 -7.660076308761752e-13
C91_107 V91 V107 -5.432961496498542e-19

R91_108 V91 V108 -869.5840970121783
L91_108 V91 V108 9.025230493028861e-12
C91_108 V91 V108 4.4595680202566386e-20

R91_109 V91 V109 436.85438774014983
L91_109 V91 V109 -1.7520689723056012e-12
C91_109 V91 V109 -4.559989090382246e-19

R91_110 V91 V110 -663.8455656820978
L91_110 V91 V110 -1.2394778353062234e-12
C91_110 V91 V110 -4.603504955495669e-19

R91_111 V91 V111 98.63706649167597
L91_111 V91 V111 2.147241035225854e-12
C91_111 V91 V111 1.474788185476054e-20

R91_112 V91 V112 2658.5935258195223
L91_112 V91 V112 3.3621205036997924e-12
C91_112 V91 V112 2.0670137683512936e-19

R91_113 V91 V113 -134.37802727939854
L91_113 V91 V113 -2.3653566502162173e-12
C91_113 V91 V113 -7.085052983348259e-20

R91_114 V91 V114 -526.9917844816252
L91_114 V91 V114 -8.439669868286981e-13
C91_114 V91 V114 -6.3491395614355135e-19

R91_115 V91 V115 213.33703470746914
L91_115 V91 V115 4.683671048111629e-13
C91_115 V91 V115 6.86854890440505e-19

R91_116 V91 V116 681.6612121085759
L91_116 V91 V116 -2.6831324218597173e-11
C91_116 V91 V116 -1.8583851689217156e-19

R91_117 V91 V117 -1439.4387932523366
L91_117 V91 V117 1.4322075081023712e-12
C91_117 V91 V117 2.8918192816982475e-19

R91_118 V91 V118 242.36257151000532
L91_118 V91 V118 7.595523349493702e-13
C91_118 V91 V118 7.492090654691467e-19

R91_119 V91 V119 -123.27265844377463
L91_119 V91 V119 -1.2387683787598063e-12
C91_119 V91 V119 7.961446978283163e-20

R91_120 V91 V120 -489.2628853648748
L91_120 V91 V120 6.173734967201336e-12
C91_120 V91 V120 2.5128706458023297e-19

R91_121 V91 V121 170.34271042155297
L91_121 V91 V121 -2.147723180827668e-11
C91_121 V91 V121 -2.1551779905378647e-19

R91_122 V91 V122 -31795.28985424691
L91_122 V91 V122 1.2638518707363945e-11
C91_122 V91 V122 1.6154414619247437e-20

R91_123 V91 V123 225.95571504479128
L91_123 V91 V123 -5.049218836738012e-13
C91_123 V91 V123 -1.2129281310747538e-18

R91_124 V91 V124 767.798935851416
L91_124 V91 V124 -6.652370750478424e-12
C91_124 V91 V124 -9.243568156145308e-20

R91_125 V91 V125 -875.3278933263668
L91_125 V91 V125 -3.1701689125278913e-12
C91_125 V91 V125 3.3593427292247086e-20

R91_126 V91 V126 -213.9683589835126
L91_126 V91 V126 -6.824892155814791e-13
C91_126 V91 V126 -6.071668963185291e-19

R91_127 V91 V127 -518.0550988999019
L91_127 V91 V127 5.208606107451949e-13
C91_127 V91 V127 7.915801668592079e-19

R91_128 V91 V128 1109.6049031007103
L91_128 V91 V128 -2.319171846994694e-12
C91_128 V91 V128 -3.860626673713987e-19

R91_129 V91 V129 -195.41977425709487
L91_129 V91 V129 -2.6428072039953944e-12
C91_129 V91 V129 -2.7454456042836414e-19

R91_130 V91 V130 406.05426744076647
L91_130 V91 V130 1.270492174043918e-12
C91_130 V91 V130 3.161916826799302e-19

R91_131 V91 V131 362.2499078308184
L91_131 V91 V131 -5.80041001853931e-12
C91_131 V91 V131 1.784604622727301e-19

R91_132 V91 V132 -2671.395783295505
L91_132 V91 V132 1.067361620143943e-12
C91_132 V91 V132 7.865043544025338e-19

R91_133 V91 V133 11544.898789656967
L91_133 V91 V133 2.4376861119201965e-12
C91_133 V91 V133 2.5355141201569897e-19

R91_134 V91 V134 -937.8715837206009
L91_134 V91 V134 9.894165780941405e-12
C91_134 V91 V134 1.7813390919571934e-19

R91_135 V91 V135 120.28657734318591
L91_135 V91 V135 -5.003730198290632e-13
C91_135 V91 V135 -1.6248421427995528e-18

R91_136 V91 V136 1343.523104054243
L91_136 V91 V136 3.790132098941205e-12
C91_136 V91 V136 2.553524283921279e-20

R91_137 V91 V137 342.7482800367797
L91_137 V91 V137 1.8136725452033666e-12
C91_137 V91 V137 1.6853304834572435e-19

R91_138 V91 V138 -944.6789729709451
L91_138 V91 V138 -1.2363812582929787e-12
C91_138 V91 V138 -4.713048593103572e-19

R91_139 V91 V139 -63.84847337476453
L91_139 V91 V139 3.201406558820393e-13
C91_139 V91 V139 2.232537325071329e-18

R91_140 V91 V140 -187.43218390273367
L91_140 V91 V140 -1.6703098659757218e-12
C91_140 V91 V140 -2.1272158401493056e-19

R91_141 V91 V141 237.81546762363797
L91_141 V91 V141 -9.94715576531213e-13
C91_141 V91 V141 -5.399117422813204e-19

R91_142 V91 V142 420.2795287874687
L91_142 V91 V142 5.792173310018108e-12
C91_142 V91 V142 -1.591848944645693e-21

R91_143 V91 V143 879.8187404256386
L91_143 V91 V143 -9.19456271507128e-13
C91_143 V91 V143 -4.1129846761075356e-19

R91_144 V91 V144 261.88570592577105
L91_144 V91 V144 2.467547179584308e-10
C91_144 V91 V144 7.723931021054308e-20

R91_145 V91 V145 -191.95372456672746
L91_145 V91 V145 -1.3987335632741876e-12
C91_145 V91 V145 -1.9448837076218223e-19

R91_146 V91 V146 744.0133330557172
L91_146 V91 V146 2.8674537421474282e-12
C91_146 V91 V146 3.2797928058188885e-19

R91_147 V91 V147 86.0206641233676
L91_147 V91 V147 -8.158366066695986e-13
C91_147 V91 V147 -1.4958580626730471e-18

R91_148 V91 V148 -489.27429581475445
L91_148 V91 V148 8.749080160687877e-12
C91_148 V91 V148 -7.165275614261747e-20

R91_149 V91 V149 -458.2007559866724
L91_149 V91 V149 5.336902801555539e-13
C91_149 V91 V149 7.379767175257264e-19

R91_150 V91 V150 -853.1254349874235
L91_150 V91 V150 -3.3059635654534393e-12
C91_150 V91 V150 -1.768736718674908e-19

R91_151 V91 V151 464.6454115012116
L91_151 V91 V151 1.5032161161136733e-12
C91_151 V91 V151 6.484796732460061e-19

R91_152 V91 V152 -638.6505013538379
L91_152 V91 V152 -3.456265859090898e-12
C91_152 V91 V152 -7.524785006808307e-20

R91_153 V91 V153 -2766.4946284509674
L91_153 V91 V153 -8.404250010264066e-11
C91_153 V91 V153 -7.585474954600745e-20

R91_154 V91 V154 4608.184943198856
L91_154 V91 V154 -3.002837238461327e-11
C91_154 V91 V154 -1.052357683273277e-19

R91_155 V91 V155 -121.42594099656245
L91_155 V91 V155 4.658303301080692e-13
C91_155 V91 V155 8.775537571181813e-19

R91_156 V91 V156 620.6975263464271
L91_156 V91 V156 1.4534862479740566e-11
C91_156 V91 V156 -1.4999092910759742e-20

R91_157 V91 V157 169.01218893709634
L91_157 V91 V157 -9.64178359642945e-13
C91_157 V91 V157 -3.9968722917200986e-19

R91_158 V91 V158 442.8754795635246
L91_158 V91 V158 2.795641381879407e-12
C91_158 V91 V158 1.8013061967460796e-19

R91_159 V91 V159 -657.6105927525447
L91_159 V91 V159 -4.667329068575967e-13
C91_159 V91 V159 -8.718725498812604e-19

R91_160 V91 V160 200.85419865958931
L91_160 V91 V160 2.514456462547076e-12
C91_160 V91 V160 1.808367937374033e-19

R91_161 V91 V161 -218.87590301405433
L91_161 V91 V161 2.489229824333817e-12
C91_161 V91 V161 1.8472614492876112e-19

R91_162 V91 V162 -722.6007289577059
L91_162 V91 V162 1.3927960423900517e-12
C91_162 V91 V162 3.270079604864162e-19

R91_163 V91 V163 -373.85146350966806
L91_163 V91 V163 2.0842477567449095e-12
C91_163 V91 V163 5.349502393889082e-19

R91_164 V91 V164 -137.7575782535692
L91_164 V91 V164 -5.591774038537416e-12
C91_164 V91 V164 1.1480693517386927e-19

R91_165 V91 V165 -195.0404735090198
L91_165 V91 V165 -1.9432390974531872e-12
C91_165 V91 V165 -2.079429989233048e-19

R91_166 V91 V166 -492.0164951522268
L91_166 V91 V166 -1.795151828862001e-12
C91_166 V91 V166 -2.360139455803569e-19

R91_167 V91 V167 232.07914537224727
L91_167 V91 V167 3.0146984059305873e-12
C91_167 V91 V167 -3.372862301134992e-20

R91_168 V91 V168 2975.1917323096923
L91_168 V91 V168 1.572241458622997e-11
C91_168 V91 V168 -3.9598355376813235e-20

R91_169 V91 V169 224.18749788066316
L91_169 V91 V169 -2.8399313445435374e-12
C91_169 V91 V169 -3.0241647495198772e-19

R91_170 V91 V170 382.9732593491009
L91_170 V91 V170 -1.936938721155614e-11
C91_170 V91 V170 2.4651215456576048e-20

R91_171 V91 V171 212.54186345615395
L91_171 V91 V171 -3.4738471251312266e-12
C91_171 V91 V171 -3.1482645867463114e-19

R91_172 V91 V172 269.5605053148674
L91_172 V91 V172 -1.773057610467494e-11
C91_172 V91 V172 -9.888959800314257e-20

R91_173 V91 V173 837.2391231383488
L91_173 V91 V173 1.0113327776614596e-12
C91_173 V91 V173 4.2782022616909627e-19

R91_174 V91 V174 534.5487398619358
L91_174 V91 V174 1.7491511347584077e-12
C91_174 V91 V174 -1.7543260291903365e-20

R91_175 V91 V175 -193.81351878434128
L91_175 V91 V175 6.77317874804236e-13
C91_175 V91 V175 8.525974939639241e-19

R91_176 V91 V176 -501.75090226939807
L91_176 V91 V176 3.8624175248307234e-12
C91_176 V91 V176 6.948292830872158e-20

R91_177 V91 V177 -263.34882920600575
L91_177 V91 V177 -1.3805339549092736e-12
C91_177 V91 V177 -1.4192374393012708e-19

R91_178 V91 V178 -402.0252375576866
L91_178 V91 V178 -2.4642913681924382e-12
C91_178 V91 V178 -2.0854319375546036e-20

R91_179 V91 V179 -162.7298673003932
L91_179 V91 V179 -8.766039091505821e-13
C91_179 V91 V179 -5.853648504483284e-19

R91_180 V91 V180 -1494.03797490889
L91_180 V91 V180 -2.2976794013495294e-12
C91_180 V91 V180 -7.650733103862282e-20

R91_181 V91 V181 414.78975597874563
L91_181 V91 V181 3.356334148152093e-12
C91_181 V91 V181 -2.0089131951184765e-19

R91_182 V91 V182 621.42111804472
L91_182 V91 V182 2.0245258397491878e-12
C91_182 V91 V182 1.3960623278879392e-19

R91_183 V91 V183 128.53631509497953
L91_183 V91 V183 -1.7811853638039977e-12
C91_183 V91 V183 -9.060927761844882e-21

R91_184 V91 V184 1668.137910560539
L91_184 V91 V184 -1.6956382036462055e-12
C91_184 V91 V184 -1.3520032475288321e-19

R91_185 V91 V185 699.4128336586442
L91_185 V91 V185 6.5798504892900854e-12
C91_185 V91 V185 2.321962382272149e-19

R91_186 V91 V186 1079.409102912393
L91_186 V91 V186 -2.205238786080143e-12
C91_186 V91 V186 -2.7931369643981377e-19

R91_187 V91 V187 1000.157154208811
L91_187 V91 V187 5.709609770052988e-13
C91_187 V91 V187 6.323266397022347e-19

R91_188 V91 V188 -2104.56849964025
L91_188 V91 V188 1.2104712533224932e-12
C91_188 V91 V188 1.759016739395369e-19

R91_189 V91 V189 -663.2699015553975
L91_189 V91 V189 -3.0490408662865996e-12
C91_189 V91 V189 -9.628657561893164e-20

R91_190 V91 V190 -787.7391680047317
L91_190 V91 V190 -9.07593035804868e-11
C91_190 V91 V190 -1.8558841343418882e-20

R91_191 V91 V191 -156.89862693227278
L91_191 V91 V191 -2.147026940645162e-12
C91_191 V91 V191 -6.005360793748737e-19

R91_192 V91 V192 -1101.636401927764
L91_192 V91 V192 2.141363956320262e-12
C91_192 V91 V192 4.033364380887533e-20

R91_193 V91 V193 -1577.9892985507042
L91_193 V91 V193 3.4342052824287946e-12
C91_193 V91 V193 2.572983587823734e-20

R91_194 V91 V194 1256.2973750820388
L91_194 V91 V194 -3.5196741477196254e-11
C91_194 V91 V194 -1.931487310077695e-19

R91_195 V91 V195 249.51298740574816
L91_195 V91 V195 3.3842048252577928e-12
C91_195 V91 V195 8.380024072563445e-19

R91_196 V91 V196 2139.9611245461733
L91_196 V91 V196 -6.595033632721112e-13
C91_196 V91 V196 -4.540336678726273e-19

R91_197 V91 V197 747.9159342660079
L91_197 V91 V197 -4.5628915182532914e-11
C91_197 V91 V197 -6.862210653657103e-21

R91_198 V91 V198 696.7411184400787
L91_198 V91 V198 8.462069816493418e-12
C91_198 V91 V198 3.0112959294842733e-20

R91_199 V91 V199 279.100053543185
L91_199 V91 V199 2.7487994490433283e-12
C91_199 V91 V199 1.1945110437972923e-19

R91_200 V91 V200 471.27090101215737
L91_200 V91 V200 1.6240006068670247e-12
C91_200 V91 V200 3.237299340392458e-19

R92_92 V92 0 -72.56912153236877
L92_92 V92 0 2.086458448643579e-13
C92_92 V92 0 1.838152200240656e-18

R92_93 V92 V93 -607.865049954682
L92_93 V92 V93 2.211917624810227e-12
C92_93 V92 V93 2.0694208308900094e-19

R92_94 V92 V94 -1592.8087209407115
L92_94 V92 V94 7.118447209152355e-12
C92_94 V92 V94 3.975711098163071e-20

R92_95 V92 V95 -949.18256085128
L92_95 V92 V95 -4.40035712094166e-11
C92_95 V92 V95 -9.383987638030816e-21

R92_96 V92 V96 -200.25734515639292
L92_96 V92 V96 1.4968940042899975e-12
C92_96 V92 V96 5.51447395614786e-20

R92_97 V92 V97 -655.1647253474338
L92_97 V92 V97 -8.692390183745678e-13
C92_97 V92 V97 -6.221571378766538e-19

R92_98 V92 V98 1513.5118916544457
L92_98 V92 V98 -7.477018595830502e-13
C92_98 V92 V98 -4.695316108177112e-19

R92_99 V92 V99 298.0483531733993
L92_99 V92 V99 1.396640814155927e-12
C92_99 V92 V99 8.353264029060061e-20

R92_100 V92 V100 43.480578279783536
L92_100 V92 V100 3.1674552808576807e-13
C92_100 V92 V100 1.4046445947417888e-18

R92_101 V92 V101 -3198.686730488276
L92_101 V92 V101 3.699889746965244e-12
C92_101 V92 V101 8.566938945142794e-20

R92_102 V92 V102 1093.2058659269035
L92_102 V92 V102 2.6093764868108127e-12
C92_102 V92 V102 8.721270599926759e-20

R92_103 V92 V103 1103.7177422151483
L92_103 V92 V103 -6.035745203550473e-12
C92_103 V92 V103 -6.87970866813449e-20

R92_104 V92 V104 -173.61036097500178
L92_104 V92 V104 -4.086202099656772e-13
C92_104 V92 V104 -9.339513208515184e-19

R92_105 V92 V105 404.5137540433322
L92_105 V92 V105 1.4529230979143414e-12
C92_105 V92 V105 3.066871096484466e-19

R92_106 V92 V106 344.25980137105364
L92_106 V92 V106 9.409510497731588e-13
C92_106 V92 V106 5.098449266743992e-19

R92_107 V92 V107 -457.57051666427503
L92_107 V92 V107 -3.171032559019133e-12
C92_107 V92 V107 -3.954688909690629e-20

R92_108 V92 V108 -66.26832439416336
L92_108 V92 V108 8.234436612463737e-12
C92_108 V92 V108 8.861179112700357e-20

R92_109 V92 V109 1057.6210097882604
L92_109 V92 V109 -2.308049332754505e-12
C92_109 V92 V109 -3.3079926265040987e-19

R92_110 V92 V110 -280.57979014378935
L92_110 V92 V110 -3.179041821981373e-12
C92_110 V92 V110 -1.3046037420314433e-19

R92_111 V92 V111 1009.7020750894939
L92_111 V92 V111 5.100442962409131e-12
C92_111 V92 V111 1.4733159224984185e-19

R92_112 V92 V112 84.89190829323054
L92_112 V92 V112 -2.0755383476628486e-12
C92_112 V92 V112 -4.1797500279415523e-19

R92_113 V92 V113 -126.14001935726202
L92_113 V92 V113 -2.137352825422293e-12
C92_113 V92 V113 -6.203776422860195e-20

R92_114 V92 V114 -509.6663502574441
L92_114 V92 V114 -8.510023633659855e-13
C92_114 V92 V114 -4.861106061020146e-19

R92_115 V92 V115 71786.02370210936
L92_115 V92 V115 -1.219145415293712e-11
C92_115 V92 V115 -1.4684959991314166e-19

R92_116 V92 V116 110.97485944389827
L92_116 V92 V116 6.280102538755216e-13
C92_116 V92 V116 3.5632788026529342e-19

R92_117 V92 V117 1881.6918114428436
L92_117 V92 V117 1.6061787283812447e-12
C92_117 V92 V117 1.849023958895144e-19

R92_118 V92 V118 174.3930744611509
L92_118 V92 V118 1.176108006359188e-12
C92_118 V92 V118 3.9355729781250928e-19

R92_119 V92 V119 -1447.0873372575252
L92_119 V92 V119 2.044827427132418e-12
C92_119 V92 V119 3.4385366781091016e-19

R92_120 V92 V120 -62.71505533682536
L92_120 V92 V120 6.803955470581088e-12
C92_120 V92 V120 7.540250225061865e-19

R92_121 V92 V121 226.81255670950026
L92_121 V92 V121 -1.0616896900209133e-11
C92_121 V92 V121 -1.4594829556683493e-19

R92_122 V92 V122 -448.0561758912248
L92_122 V92 V122 3.7737241474951846e-12
C92_122 V92 V122 2.0353566915312527e-19

R92_123 V92 V123 1864.789704656591
L92_123 V92 V123 -3.999690875732009e-12
C92_123 V92 V123 -4.6045226924342064e-20

R92_124 V92 V124 129.56764540692154
L92_124 V92 V124 -3.2945726563554557e-13
C92_124 V92 V124 -1.6773543993363454e-18

R92_125 V92 V125 -538.5500203733893
L92_125 V92 V125 -2.721106967815269e-12
C92_125 V92 V125 3.288345019106649e-20

R92_126 V92 V126 -197.71159335759327
L92_126 V92 V126 -7.457430014223018e-13
C92_126 V92 V126 -3.7445096529121993e-19

R92_127 V92 V127 -409.0159037304493
L92_127 V92 V127 -7.895826113464757e-13
C92_127 V92 V127 -5.580252932636508e-19

R92_128 V92 V128 367.4367374371558
L92_128 V92 V128 5.760721894364376e-13
C92_128 V92 V128 4.523331028497977e-19

R92_129 V92 V129 -270.1067776421539
L92_129 V92 V129 7.383086066661756e-11
C92_129 V92 V129 -1.0293959926219167e-19

R92_130 V92 V130 303.9126649843481
L92_130 V92 V130 1.8183613001524069e-12
C92_130 V92 V130 1.0079227855144133e-19

R92_131 V92 V131 390.62078188705294
L92_131 V92 V131 8.399505769816396e-13
C92_131 V92 V131 5.755700919413743e-19

R92_132 V92 V132 -541.3309867792086
L92_132 V92 V132 1.8068965820619068e-12
C92_132 V92 V132 6.258770389442005e-19

R92_133 V92 V133 -1115.378550607565
L92_133 V92 V133 3.2400748387168694e-12
C92_133 V92 V133 2.0498682857533598e-19

R92_134 V92 V134 -424.63326442090107
L92_134 V92 V134 1.5945364585849366e-12
C92_134 V92 V134 6.018197769612205e-19

R92_135 V92 V135 -1394.4318915310275
L92_135 V92 V135 1.870570232366547e-12
C92_135 V92 V135 2.96587088192404e-19

R92_136 V92 V136 106.60488323436883
L92_136 V92 V136 -4.465337336537161e-13
C92_136 V92 V136 -1.370022090575552e-18

R92_137 V92 V137 266.7326714272041
L92_137 V92 V137 -4.2004489523804745e-12
C92_137 V92 V137 -1.9990975337562833e-19

R92_138 V92 V138 5203.7653148970785
L92_138 V92 V138 -9.328456193752133e-13
C92_138 V92 V138 -6.541796158231545e-19

R92_139 V92 V139 -328.5676618160029
L92_139 V92 V139 -7.979620756068991e-13
C92_139 V92 V139 -6.231826470656044e-19

R92_140 V92 V140 -60.40569756293364
L92_140 V92 V140 4.1789052554410667e-13
C92_140 V92 V140 1.615839056664981e-18

R92_141 V92 V141 307.6404815214898
L92_141 V92 V141 -1.865729394102766e-12
C92_141 V92 V141 -9.572697585958679e-20

R92_142 V92 V142 921.4461484876417
L92_142 V92 V142 -3.529631629416457e-12
C92_142 V92 V142 -9.816006380139673e-20

R92_143 V92 V143 351.535031550967
L92_143 V92 V143 -2.3159642239233387e-11
C92_143 V92 V143 1.4318745775208677e-19

R92_144 V92 V144 -1265.0593255100894
L92_144 V92 V144 -2.3371115194501193e-12
C92_144 V92 V144 -3.0918489579452217e-19

R92_145 V92 V145 -178.8359877506301
L92_145 V92 V145 9.628798826031718e-12
C92_145 V92 V145 1.1402466174974986e-19

R92_146 V92 V146 981.6572021978924
L92_146 V92 V146 1.0061923371173869e-12
C92_146 V92 V146 3.263351306731535e-19

R92_147 V92 V147 1080.2925384982198
L92_147 V92 V147 2.920911335590903e-11
C92_147 V92 V147 -8.979446860654996e-20

R92_148 V92 V148 64.71653180844237
L92_148 V92 V148 -4.156477589824265e-13
C92_148 V92 V148 -1.0400955944222007e-18

R92_149 V92 V149 -436.9086825557492
L92_149 V92 V149 1.8983674028233082e-12
C92_149 V92 V149 -3.0485863600510227e-20

R92_150 V92 V150 4154.833178982672
L92_150 V92 V150 -2.106189772848718e-12
C92_150 V92 V150 3.621019179446125e-20

R92_151 V92 V151 -543.6666298703301
L92_151 V92 V151 4.036997643255528e-12
C92_151 V92 V151 -3.9139308987869115e-20

R92_152 V92 V152 8886.51792618413
L92_152 V92 V152 5.629434191500275e-13
C92_152 V92 V152 4.275836680405413e-19

R92_153 V92 V153 949.1696064654388
L92_153 V92 V153 2.268425875266645e-12
C92_153 V92 V153 -5.537618902533279e-21

R92_154 V92 V154 -418875.12857629574
L92_154 V92 V154 2.608576145415627e-12
C92_154 V92 V154 -2.626560230672026e-19

R92_155 V92 V155 389.3904999807815
L92_155 V92 V155 3.582613563552195e-12
C92_155 V92 V155 -6.69487619084078e-20

R92_156 V92 V156 -170.41941427370153
L92_156 V92 V156 4.404552211410017e-12
C92_156 V92 V156 7.831233335387915e-19

R92_157 V92 V157 158.08649517314385
L92_157 V92 V157 -1.1236631758084217e-12
C92_157 V92 V157 -1.4398381598923383e-19

R92_158 V92 V158 312.09919994060033
L92_158 V92 V158 -9.57505154834276e-12
C92_158 V92 V158 1.365010471181251e-19

R92_159 V92 V159 255.76884806728512
L92_159 V92 V159 3.710009373073562e-12
C92_159 V92 V159 1.9413542134661504e-19

R92_160 V92 V160 -181.16222465496682
L92_160 V92 V160 -8.971692630962768e-13
C92_160 V92 V160 -6.784929597106605e-19

R92_161 V92 V161 -292.0208855635417
L92_161 V92 V161 1.0011388743465456e-12
C92_161 V92 V161 2.9989096644310466e-19

R92_162 V92 V162 -633.0856821571457
L92_162 V92 V162 1.7950397753324505e-12
C92_162 V92 V162 1.587245250484475e-19

R92_163 V92 V163 -204.58961717241584
L92_163 V92 V163 -7.808921759720175e-11
C92_163 V92 V163 2.4294988935906916e-20

R92_164 V92 V164 653.1241273196657
L92_164 V92 V164 7.980918439050796e-12
C92_164 V92 V164 4.291364442134195e-19

R92_165 V92 V165 -246.7643084261614
L92_165 V92 V165 -1.0964002806109162e-12
C92_165 V92 V165 -3.226592157695931e-19

R92_166 V92 V166 -526.1765836554822
L92_166 V92 V166 -1.7107318300319161e-12
C92_166 V92 V166 -2.0617385307022006e-19

R92_167 V92 V167 481.06070178287683
L92_167 V92 V167 9.493838813220802e-12
C92_167 V92 V167 1.1566468880338842e-19

R92_168 V92 V168 657.8215868779707
L92_168 V92 V168 8.644540668565113e-13
C92_168 V92 V168 5.517491226498123e-20

R92_169 V92 V169 247.14127079796216
L92_169 V92 V169 -2.5503489544445688e-12
C92_169 V92 V169 -3.3986146320318565e-19

R92_170 V92 V170 253.68586755451832
L92_170 V92 V170 2.5539451879734273e-12
C92_170 V92 V170 -3.8750117029531845e-20

R92_171 V92 V171 273.39732168624874
L92_171 V92 V171 2.574415776394e-12
C92_171 V92 V171 -1.5101201496387114e-19

R92_172 V92 V172 210.91920547616985
L92_172 V92 V172 -7.736755165408803e-13
C92_172 V92 V172 -3.5679391066136376e-19

R92_173 V92 V173 487.4815531216823
L92_173 V92 V173 8.928306496840049e-13
C92_173 V92 V173 3.9615940009734523e-19

R92_174 V92 V174 -2839.740509004044
L92_174 V92 V174 9.647875651870761e-12
C92_174 V92 V174 4.5011984062586924e-20

R92_175 V92 V175 -481.4876952142982
L92_175 V92 V175 -1.975577100923312e-12
C92_175 V92 V175 -9.502980859509358e-20

R92_176 V92 V176 -237.80836696998284
L92_176 V92 V176 7.035237615704248e-13
C92_176 V92 V176 7.98909201075213e-19

R92_177 V92 V177 -366.74521079894384
L92_177 V92 V177 -2.0836227571199853e-12
C92_177 V92 V177 -1.1191371143143964e-19

R92_178 V92 V178 -666.6750813294229
L92_178 V92 V178 -2.929073231117578e-12
C92_178 V92 V178 1.967764616944033e-20

R92_179 V92 V179 938.158272575523
L92_179 V92 V179 -5.3795299798426305e-12
C92_179 V92 V179 5.899928729861225e-20

R92_180 V92 V180 -93.9685538174975
L92_180 V92 V180 -8.793706465668941e-13
C92_180 V92 V180 -4.935060776117683e-19

R92_181 V92 V181 831.2894640139939
L92_181 V92 V181 4.204800016537196e-11
C92_181 V92 V181 -5.0288881537463444e-20

R92_182 V92 V182 519.9582611462022
L92_182 V92 V182 -5.257311738042328e-11
C92_182 V92 V182 -1.0960917756793989e-19

R92_183 V92 V183 -586.0747388178751
L92_183 V92 V183 -2.1099666358849434e-12
C92_183 V92 V183 -1.4251495555185992e-19

R92_184 V92 V184 109.44099199243874
L92_184 V92 V184 -2.214487519390005e-12
C92_184 V92 V184 1.402258343379629e-20

R92_185 V92 V185 414.47289061850125
L92_185 V92 V185 4.484860687815399e-12
C92_185 V92 V185 1.1301460197829603e-19

R92_186 V92 V186 -1551.8842605429052
L92_186 V92 V186 -1.6843677595629021e-12
C92_186 V92 V186 1.5681002799036922e-20

R92_187 V92 V187 -380.36931209652124
L92_187 V92 V187 -4.52723409910245e-12
C92_187 V92 V187 3.345274950134225e-20

R92_188 V92 V188 226.80196965381987
L92_188 V92 V188 3.802523125574045e-13
C92_188 V92 V188 3.3628561830204984e-19

R92_189 V92 V189 -676.9726966356532
L92_189 V92 V189 -1.7211977555256241e-12
C92_189 V92 V189 -2.199440195538017e-19

R92_190 V92 V190 -2998.2058190525263
L92_190 V92 V190 4.709500998622337e-12
C92_190 V92 V190 8.968466529323415e-20

R92_191 V92 V191 364.8973935421513
L92_191 V92 V191 7.842928829800218e-13
C92_191 V92 V191 1.6386048640772583e-19

R92_192 V92 V192 -104.33553906741614
L92_192 V92 V192 -4.4835125010330823e-13
C92_192 V92 V192 -6.770756899818489e-19

R92_193 V92 V193 -377.2196978761685
L92_193 V92 V193 1.0121112217592744e-11
C92_193 V92 V193 -4.135536750287368e-20

R92_194 V92 V194 861.2121771564994
L92_194 V92 V194 -1.348929145469131e-12
C92_194 V92 V194 -4.330518256026634e-19

R92_195 V92 V195 -3313.2875223809497
L92_195 V92 V195 -5.801259037982942e-13
C92_195 V92 V195 -5.540146695213102e-19

R92_196 V92 V196 171.63147075026833
L92_196 V92 V196 4.3421805989434087e-13
C92_196 V92 V196 1.3509645399337645e-18

R92_197 V92 V197 837.6244866835171
L92_197 V92 V197 2.595910626149685e-12
C92_197 V92 V197 2.2669643610544224e-19

R92_198 V92 V198 674.2502908948194
L92_198 V92 V198 7.676670612031981e-11
C92_198 V92 V198 -1.0738892969522842e-19

R92_199 V92 V199 412.7195746157188
L92_199 V92 V199 2.0229661080447426e-12
C92_199 V92 V199 2.771938402292653e-19

R92_200 V92 V200 354.50031908043377
L92_200 V92 V200 1.4886988297548365e-11
C92_200 V92 V200 -2.319560532329703e-19

R93_93 V93 0 98.37761325364606
L93_93 V93 0 -6.180732981465109e-13
C93_93 V93 0 -8.207863249727411e-20

R93_94 V93 V94 -1091.7725646217673
L93_94 V93 V94 -2.514476388082401e-12
C93_94 V93 V94 -3.4647157634858373e-19

R93_95 V93 V95 1009.3732705172283
L93_95 V93 V95 -4.38479211385714e-12
C93_95 V93 V95 -1.7147083885184058e-19

R93_96 V93 V96 1799.4409200054847
L93_96 V93 V96 -2.7150066577164338e-12
C93_96 V93 V96 -2.3436107300905405e-19

R93_97 V93 V97 378.3135703496902
L93_97 V93 V97 1.2039625072673296e-11
C93_97 V93 V97 -1.0714780564558069e-19

R93_98 V93 V98 184.23702184933452
L93_98 V93 V98 5.875040022137645e-12
C93_98 V93 V98 5.378115243898872e-20

R93_99 V93 V99 333.7285938938435
L93_99 V93 V99 -2.2579072786791665e-12
C93_99 V93 V99 -2.123674848198325e-19

R93_100 V93 V100 796.7805012656426
L93_100 V93 V100 -2.549504608479168e-12
C93_100 V93 V100 -1.294296082742483e-19

R93_101 V93 V101 131.46770317747126
L93_101 V93 V101 2.281425927849917e-12
C93_101 V93 V101 3.986478593186686e-19

R93_102 V93 V102 -588.8872019324776
L93_102 V93 V102 1.0611772688723515e-11
C93_102 V93 V102 1.60872666269752e-19

R93_103 V93 V103 -690.8575767477719
L93_103 V93 V103 2.8106313780520175e-12
C93_103 V93 V103 2.186064019083166e-19

R93_104 V93 V104 -1729.4984277804956
L93_104 V93 V104 2.5967999643627966e-12
C93_104 V93 V104 2.204693313269e-19

R93_105 V93 V105 -74.334921390474
L93_105 V93 V105 1.7195170290882618e-11
C93_105 V93 V105 1.932386417588319e-19

R93_106 V93 V106 -1257.542872663203
L93_106 V93 V106 -4.9805641765926615e-12
C93_106 V93 V106 -1.4486835488746056e-19

R93_107 V93 V107 1596.0944997771894
L93_107 V93 V107 1.3245725595209717e-11
C93_107 V93 V107 3.6273294289496757e-20

R93_108 V93 V108 705.6864809952733
L93_108 V93 V108 7.973297403803048e-12
C93_108 V93 V108 7.533951230873903e-20

R93_109 V93 V109 3905.2496179002233
L93_109 V93 V109 3.1734865614397646e-12
C93_109 V93 V109 -7.922604491086726e-20

R93_110 V93 V110 524.3608083154543
L93_110 V93 V110 -6.001755442367359e-11
C93_110 V93 V110 -4.9504679505902546e-21

R93_111 V93 V111 2563.6112185620823
L93_111 V93 V111 3.2893594903749706e-11
C93_111 V93 V111 -2.091984606701736e-20

R93_112 V93 V112 -4049.991783072943
L93_112 V93 V112 -3.928702117229437e-10
C93_112 V93 V112 -7.70829262826278e-20

R93_113 V93 V113 111.25322382716558
L93_113 V93 V113 -2.520506262025489e-12
C93_113 V93 V113 -4.1125771875792363e-19

R93_114 V93 V114 -14461.274169699273
L93_114 V93 V114 4.50063154792002e-12
C93_114 V93 V114 7.231524172607295e-20

R93_115 V93 V115 -1274.1357278715332
L93_115 V93 V115 -6.875583870998871e-12
C93_115 V93 V115 -6.483995139397976e-20

R93_116 V93 V116 -821.8637297330243
L93_116 V93 V116 -3.6665049979266555e-12
C93_116 V93 V116 -1.5456430570639296e-19

R93_117 V93 V117 -202.34592499385607
L93_117 V93 V117 -4.309245254601201e-12
C93_117 V93 V117 2.8683051690440373e-22

R93_118 V93 V118 -897.549394886125
L93_118 V93 V118 3.752784522084094e-11
C93_118 V93 V118 5.130987186404691e-20

R93_119 V93 V119 1272.9136076040525
L93_119 V93 V119 -3.856098054047598e-11
C93_119 V93 V119 2.548752518894364e-20

R93_120 V93 V120 519.9773369581894
L93_120 V93 V120 1.7129201854453225e-10
C93_120 V93 V120 7.272344553601117e-20

R93_121 V93 V121 -223.49334670667363
L93_121 V93 V121 3.211561563589427e-12
C93_121 V93 V121 3.214519742047354e-19

R93_122 V93 V122 1321.9830820648472
L93_122 V93 V122 -3.3242048727245343e-12
C93_122 V93 V122 -1.8392733893912038e-19

R93_123 V93 V123 -6027.033171246213
L93_123 V93 V123 5.7465257559438934e-12
C93_123 V93 V123 7.381704228014073e-20

R93_124 V93 V124 -960.643639125768
L93_124 V93 V124 3.281042410348001e-12
C93_124 V93 V124 1.2365055186007946e-19

R93_125 V93 V125 -850.16804282175
L93_125 V93 V125 4.912285067963512e-12
C93_125 V93 V125 1.0083169668082495e-19

R93_126 V93 V126 1086.4595965028866
L93_126 V93 V126 4.535019454978538e-12
C93_126 V93 V126 1.4421215320785812e-19

R93_127 V93 V127 1867.6674406055422
L93_127 V93 V127 -1.3399600358301375e-11
C93_127 V93 V127 -2.741795443990574e-20

R93_128 V93 V128 4032.852390796058
L93_128 V93 V128 -2.5894992571135533e-11
C93_128 V93 V128 1.1538217097773068e-20

R93_129 V93 V129 308.2777020538701
L93_129 V93 V129 -7.220079772285774e-12
C93_129 V93 V129 -1.4760437402373787e-19

R93_130 V93 V130 5029.954484229315
L93_130 V93 V130 7.183486750040305e-12
C93_130 V93 V130 9.646773043673741e-20

R93_131 V93 V131 744650.6395720784
L93_131 V93 V131 -3.160470179765672e-10
C93_131 V93 V131 -5.766593280924635e-20

R93_132 V93 V132 1081.2390160165437
L93_132 V93 V132 -7.333434553787365e-12
C93_132 V93 V132 -1.505574099412844e-19

R93_133 V93 V133 338.62385371511374
L93_133 V93 V133 9.452857287964112e-12
C93_133 V93 V133 -1.2404506642538593e-19

R93_134 V93 V134 -1163.52461383673
L93_134 V93 V134 -2.9542166563919134e-12
C93_134 V93 V134 -3.16523073245737e-19

R93_135 V93 V135 -422.2736504623187
L93_135 V93 V135 5.834408747694214e-12
C93_135 V93 V135 1.6584504545605037e-19

R93_136 V93 V136 -291.540403951789
L93_136 V93 V136 1.2925690503769967e-11
C93_136 V93 V136 -1.815498258890037e-21

R93_137 V93 V137 -128.1376502715567
L93_137 V93 V137 -3.774259395053356e-12
C93_137 V93 V137 -2.26170396935976e-20

R93_138 V93 V138 -1166.6359005023605
L93_138 V93 V138 7.722866558297734e-12
C93_138 V93 V138 2.0662867131639852e-19

R93_139 V93 V139 369.84801282590155
L93_139 V93 V139 -4.355120132799043e-12
C93_139 V93 V139 -1.6334599176749272e-19

R93_140 V93 V140 319.35940166781097
L93_140 V93 V140 -3.5619825835570877e-12
C93_140 V93 V140 -8.975370419916142e-20

R93_141 V93 V141 -2324.5880985245376
L93_141 V93 V141 3.5978942444325346e-12
C93_141 V93 V141 1.5552841373744746e-19

R93_142 V93 V142 233.6925185657202
L93_142 V93 V142 2.939462358738199e-12
C93_142 V93 V142 1.3466857436372362e-19

R93_143 V93 V143 419.53022649993403
L93_143 V93 V143 -1.0335876674398296e-10
C93_143 V93 V143 -1.0260664751024328e-19

R93_144 V93 V144 247.57891545083874
L93_144 V93 V144 4.384657040542251e-12
C93_144 V93 V144 1.1192094860958578e-19

R93_145 V93 V145 194.81765548684047
L93_145 V93 V145 8.02908050276988e-12
C93_145 V93 V145 -4.303125409131832e-20

R93_146 V93 V146 496.71724566762333
L93_146 V93 V146 -4.144294709803785e-12
C93_146 V93 V146 -1.3455033755481687e-19

R93_147 V93 V147 -723.2111655743122
L93_147 V93 V147 4.356941393123226e-12
C93_147 V93 V147 2.870903872684443e-19

R93_148 V93 V148 -215.77641641836607
L93_148 V93 V148 4.1381651969139196e-12
C93_148 V93 V148 1.157948283673501e-19

R93_149 V93 V149 259.0159798945135
L93_149 V93 V149 -5.704155482470122e-11
C93_149 V93 V149 3.042975704362472e-19

R93_150 V93 V150 -126.72928351944554
L93_150 V93 V150 7.000444217603553e-12
C93_150 V93 V150 -1.4650006509899565e-19

R93_151 V93 V151 -233.52682034163456
L93_151 V93 V151 9.19423800428665e-12
C93_151 V93 V151 3.2301555532613744e-20

R93_152 V93 V152 -1065.2311321842951
L93_152 V93 V152 -4.973300508390267e-12
C93_152 V93 V152 -9.628237498938761e-20

R93_153 V93 V153 -113.58022972240624
L93_153 V93 V153 -4.6072612230843366e-11
C93_153 V93 V153 -1.3066241935778923e-19

R93_154 V93 V154 -631.836624064669
L93_154 V93 V154 -4.634011160367222e-12
C93_154 V93 V154 1.5198376968827831e-19

R93_155 V93 V155 248.7131706810953
L93_155 V93 V155 -4.403677916071129e-12
C93_155 V93 V155 -1.844923908182462e-20

R93_156 V93 V156 -1279.7723547775738
L93_156 V93 V156 -1.022287022940878e-11
C93_156 V93 V156 -8.059946431680954e-20

R93_157 V93 V157 -153.5898744153326
L93_157 V93 V157 -3.635245748977803e-12
C93_157 V93 V157 -4.607417697309354e-19

R93_158 V93 V158 211.53453644488624
L93_158 V93 V158 4.9876326321048556e-11
C93_158 V93 V158 -6.938673609220153e-20

R93_159 V93 V159 2029.95924338202
L93_159 V93 V159 -6.660555373566631e-11
C93_159 V93 V159 -6.484665597510805e-20

R93_160 V93 V160 221.0522554691475
L93_160 V93 V160 -4.2621275444757195e-11
C93_160 V93 V160 3.3411975879769046e-20

R93_161 V93 V161 455.60488531189
L93_161 V93 V161 -4.003364796314117e-12
C93_161 V93 V161 1.1179002361905313e-19

R93_162 V93 V162 332.7964081856171
L93_162 V93 V162 1.0951887666589752e-10
C93_162 V93 V162 -1.1404398226378185e-19

R93_163 V93 V163 425.7970477436483
L93_163 V93 V163 -3.179484003441146e-12
C93_163 V93 V163 -2.293334763655211e-19

R93_164 V93 V164 2569.9273786407457
L93_164 V93 V164 -5.521352543786605e-11
C93_164 V93 V164 -4.282510681796373e-20

R93_165 V93 V165 1347.2451143220476
L93_165 V93 V165 8.922077440426932e-13
C93_165 V93 V165 4.677916860145819e-19

R93_166 V93 V166 -214.38169086862652
L93_166 V93 V166 2.6698093878902188e-12
C93_166 V93 V166 1.4006884450366957e-19

R93_167 V93 V167 -629.5047880272269
L93_167 V93 V167 6.7907318081451044e-12
C93_167 V93 V167 1.0344823585066043e-19

R93_168 V93 V168 708.9916713467495
L93_168 V93 V168 1.5586058711543836e-11
C93_168 V93 V168 1.3604668772166358e-19

R93_169 V93 V169 -266.82864071014615
L93_169 V93 V169 -3.354132077744099e-12
C93_169 V93 V169 -2.657182197183985e-19

R93_170 V93 V170 -1623.9435171920672
L93_170 V93 V170 -5.081630735056082e-12
C93_170 V93 V170 1.6047249859729353e-19

R93_171 V93 V171 -558.8076600193276
L93_171 V93 V171 2.3922099811734302e-12
C93_171 V93 V171 3.3718395110512997e-19

R93_172 V93 V172 -581.2952646970631
L93_172 V93 V172 3.999597066187127e-12
C93_172 V93 V172 1.3285611235225522e-19

R93_173 V93 V173 -472.30365485591335
L93_173 V93 V173 -1.1867593171660197e-12
C93_173 V93 V173 -2.66797500360347e-19

R93_174 V93 V174 198.42127387548666
L93_174 V93 V174 -2.5525097528170882e-12
C93_174 V93 V174 -3.434812041681746e-19

R93_175 V93 V175 561.2344806499473
L93_175 V93 V175 -3.272382640534493e-12
C93_175 V93 V175 -2.766882256351043e-19

R93_176 V93 V176 974.2366223081574
L93_176 V93 V176 -2.6054173909727935e-12
C93_176 V93 V176 -3.014031208163275e-19

R93_177 V93 V177 481.66049913637465
L93_177 V93 V177 1.4533086871545086e-12
C93_177 V93 V177 2.9495638409550796e-19

R93_178 V93 V178 -374.79412185032476
L93_178 V93 V178 4.932694506390032e-12
C93_178 V93 V178 -5.990232153017755e-20

R93_179 V93 V179 890.9977623651263
L93_179 V93 V179 -5.073996932890483e-12
C93_179 V93 V179 -1.3128519266561924e-19

R93_180 V93 V180 852.9617907371126
L93_180 V93 V180 -5.6456280340579225e-11
C93_180 V93 V180 -4.116382774289963e-20

R93_181 V93 V181 -41267.34886505619
L93_181 V93 V181 -5.563452883671261e-12
C93_181 V93 V181 2.1359815969672971e-19

R93_182 V93 V182 -530.8141491845377
L93_182 V93 V182 3.3549138884098996e-12
C93_182 V93 V182 1.7361434432117818e-19

R93_183 V93 V183 -807.2321050572466
L93_183 V93 V183 3.037755998807923e-10
C93_183 V93 V183 5.39887231938701e-21

R93_184 V93 V184 -852.1451812507305
L93_184 V93 V184 6.002727134429963e-12
C93_184 V93 V184 1.1990390258285415e-19

R93_185 V93 V185 -257.41113838776874
L93_185 V93 V185 -1.7644311702694283e-11
C93_185 V93 V185 -3.3635502752213947e-19

R93_186 V93 V186 297.315547146617
L93_186 V93 V186 2.8511799514617735e-12
C93_186 V93 V186 2.1149716866116888e-19

R93_187 V93 V187 1073.1104955292262
L93_187 V93 V187 3.8497989253440435e-12
C93_187 V93 V187 1.0652085819029355e-19

R93_188 V93 V188 -47636.79590152585
L93_188 V93 V188 3.382305714348834e-11
C93_188 V93 V188 1.1355785052134667e-19

R93_189 V93 V189 240.6434846735206
L93_189 V93 V189 3.87830495287796e-12
C93_189 V93 V189 9.958956925068881e-20

R93_190 V93 V190 -1412.9936933184854
L93_190 V93 V190 -5.0078049479176125e-12
C93_190 V93 V190 -1.8969026975006738e-19

R93_191 V93 V191 -522.2374541544958
L93_191 V93 V191 3.687634897045795e-12
C93_191 V93 V191 1.6919132821733758e-19

R93_192 V93 V192 -5024.255088761963
L93_192 V93 V192 4.661506843877344e-12
C93_192 V93 V192 -8.548056350112499e-22

R93_193 V93 V193 682.6143380543817
L93_193 V93 V193 -1.6957267761045945e-12
C93_193 V93 V193 -1.3813497100004603e-19

R93_194 V93 V194 -390.1542222350697
L93_194 V93 V194 -3.515534552155595e-12
C93_194 V93 V194 -1.5502501794548343e-19

R93_195 V93 V195 -9086.6151169678
L93_195 V93 V195 -2.8536295497736126e-12
C93_195 V93 V195 -2.80536071612003e-19

R93_196 V93 V196 -652.9323691962437
L93_196 V93 V196 -1.801257777088358e-12
C93_196 V93 V196 -3.084018115216318e-19

R93_197 V93 V197 -294.1379853082268
L93_197 V93 V197 3.4249655441053755e-11
C93_197 V93 V197 1.3616129699773708e-19

R93_198 V93 V198 2103.3238385515083
L93_198 V93 V198 6.176664176479367e-12
C93_198 V93 V198 8.881690465229194e-20

R93_199 V93 V199 579.6653104437025
L93_199 V93 V199 -2.9906200273284808e-12
C93_199 V93 V199 -2.253237055005369e-19

R93_200 V93 V200 355.0688078437393
L93_200 V93 V200 -9.690794839486445e-12
C93_200 V93 V200 9.45356078343443e-20

R94_94 V94 0 1287.6138887208972
L94_94 V94 0 5.893086956499229e-13
C94_94 V94 0 1.8208208694198314e-18

R94_95 V94 V95 -746.1302808803074
L94_95 V94 V95 -7.750058458994822e-12
C94_95 V94 V95 -1.2382572715275255e-19

R94_96 V94 V96 -661.9935840696093
L94_96 V94 V96 -4.121298689287258e-12
C94_96 V94 V96 -2.1060861972694088e-19

R94_97 V94 V97 -1430.8060789882193
L94_97 V94 V97 -1.661986048312092e-12
C94_97 V94 V97 -4.5122335875974655e-19

R94_98 V94 V98 299.74077359633543
L94_98 V94 V98 9.866747359168053e-12
C94_98 V94 V98 -1.2926578599665215e-19

R94_99 V94 V99 412.9302821455228
L94_99 V94 V99 3.6317235288872507e-12
C94_99 V94 V99 2.5823613002663824e-19

R94_100 V94 V100 1029.2252248322159
L94_100 V94 V100 -7.4385672301474e-12
C94_100 V94 V100 1.2043017399596018e-19

R94_101 V94 V101 -7356.647141504007
L94_101 V94 V101 2.0659549723968357e-12
C94_101 V94 V101 3.992325694437775e-19

R94_102 V94 V102 219.1079165688303
L94_102 V94 V102 8.33129999879339e-13
C94_102 V94 V102 8.82365274130266e-19

R94_103 V94 V103 942.9352356268502
L94_103 V94 V103 5.352608155840044e-12
C94_103 V94 V103 5.956925504959649e-20

R94_104 V94 V104 454.2247468596382
L94_104 V94 V104 5.941318267812348e-12
C94_104 V94 V104 6.0929061813969854e-21

R94_105 V94 V105 18272.08826054975
L94_105 V94 V105 2.790585314576614e-12
C94_105 V94 V105 2.971052773607033e-19

R94_106 V94 V106 -156.97823523684386
L94_106 V94 V106 -1.4762146219919735e-12
C94_106 V94 V106 -3.538328543355997e-19

R94_107 V94 V107 -533.7825288974743
L94_107 V94 V107 -2.480760858190112e-12
C94_107 V94 V107 -2.51327809386615e-19

R94_108 V94 V108 -662.9593093980285
L94_108 V94 V108 6.315374212790804e-12
C94_108 V94 V108 9.372750795197216e-20

R94_109 V94 V109 584.4360894999264
L94_109 V94 V109 -4.045356542213662e-12
C94_109 V94 V109 -3.1633147168005743e-19

R94_110 V94 V110 3005.573865961807
L94_110 V94 V110 -3.046461664684613e-12
C94_110 V94 V110 -3.7075987331527133e-19

R94_111 V94 V111 -821.1485616331914
L94_111 V94 V111 6.022103062464685e-11
C94_111 V94 V111 3.736764441731781e-20

R94_112 V94 V112 -591.3028506770294
L94_112 V94 V112 -9.39374980789625e-11
C94_112 V94 V112 -1.5636079372079774e-20

R94_113 V94 V113 -398.718146350242
L94_113 V94 V113 -2.126359392432618e-12
C94_113 V94 V113 -4.1758938121452785e-19

R94_114 V94 V114 225.25694451341778
L94_114 V94 V114 3.0847033484504765e-12
C94_114 V94 V114 1.5707412129171885e-19

R94_115 V94 V115 391.65490839218825
L94_115 V94 V115 2.4271747745520986e-12
C94_115 V94 V115 1.9828331126587538e-19

R94_116 V94 V116 430.5017600405481
L94_116 V94 V116 -8.84015817160079e-12
C94_116 V94 V116 -1.524319693169337e-19

R94_117 V94 V117 -313.0077034986677
L94_117 V94 V117 4.410031509165582e-12
C94_117 V94 V117 2.633434311202599e-19

R94_118 V94 V118 -334.7916733303791
L94_118 V94 V118 1.4031844363677315e-12
C94_118 V94 V118 5.691754703792584e-19

R94_119 V94 V119 6014.747812362905
L94_119 V94 V119 -5.996569679817734e-12
C94_119 V94 V119 1.3220008297842157e-20

R94_120 V94 V120 1217.4810043293683
L94_120 V94 V120 2.78397188962812e-11
C94_120 V94 V120 2.1607807855514007e-19

R94_121 V94 V121 207.62197049793704
L94_121 V94 V121 2.6477642167322575e-12
C94_121 V94 V121 2.654078202859249e-19

R94_122 V94 V122 -3102.1429487744717
L94_122 V94 V122 -1.0940670957677471e-12
C94_122 V94 V122 -5.816269509905337e-19

R94_123 V94 V123 -442.0399648527611
L94_123 V94 V123 1.7454686704242758e-11
C94_123 V94 V123 -4.1297200347301006e-20

R94_124 V94 V124 -372.72839050713986
L94_124 V94 V124 6.9674398683945686e-12
C94_124 V94 V124 -7.321065014231649e-20

R94_125 V94 V125 471.81641461082796
L94_125 V94 V125 -1.5471681904306743e-11
C94_125 V94 V125 -7.505703191791978e-20

R94_126 V94 V126 436.18904344827496
L94_126 V94 V126 -5.523106653709663e-12
C94_126 V94 V126 -2.1070450078168304e-19

R94_127 V94 V127 1184.4291745649882
L94_127 V94 V127 -8.884928524326951e-12
C94_127 V94 V127 -1.0991423608291082e-19

R94_128 V94 V128 1611.6528395365988
L94_128 V94 V128 -9.378209111012586e-12
C94_128 V94 V128 -1.1784843859578864e-19

R94_129 V94 V129 -139.99315088245956
L94_129 V94 V129 -1.2134777298918283e-12
C94_129 V94 V129 -5.43677874544553e-19

R94_130 V94 V130 -527.585279569737
L94_130 V94 V130 1.2044181360354052e-12
C94_130 V94 V130 6.407525910862719e-19

R94_131 V94 V131 1230.3377585946014
L94_131 V94 V131 -2.3599951763519987e-11
C94_131 V94 V131 5.419109242233337e-20

R94_132 V94 V132 790.467895725573
L94_132 V94 V132 2.2352909823945026e-11
C94_132 V94 V132 1.8460942629073536e-19

R94_133 V94 V133 958.487837882997
L94_133 V94 V133 1.227312749762303e-12
C94_133 V94 V133 4.913796574212183e-19

R94_134 V94 V134 1269.3135025982838
L94_134 V94 V134 -1.3583781657530258e-12
C94_134 V94 V134 -5.816342740771232e-19

R94_135 V94 V135 -1094.5942482169269
L94_135 V94 V135 2.279459465513776e-12
C94_135 V94 V135 1.8955544168682191e-19

R94_136 V94 V136 -535.9343735441632
L94_136 V94 V136 7.907931937730679e-12
C94_136 V94 V136 -1.0825992499031348e-19

R94_137 V94 V137 196.5825142885292
L94_137 V94 V137 1.8301671103046166e-12
C94_137 V94 V137 2.7357408581813467e-19

R94_138 V94 V138 478.62320444365935
L94_138 V94 V138 3.2511407227860376e-12
C94_138 V94 V138 2.070758540224567e-19

R94_139 V94 V139 769.6297681658215
L94_139 V94 V139 -6.552663226045296e-12
C94_139 V94 V139 -2.262417055391143e-20

R94_140 V94 V140 303.25989271140907
L94_140 V94 V140 -6.201433974612586e-12
C94_140 V94 V140 5.916688780975322e-20

R94_141 V94 V141 -1642.8703366369225
L94_141 V94 V141 -8.362502379498419e-13
C94_141 V94 V141 -7.370094014616114e-19

R94_142 V94 V142 -477.80707073805394
L94_142 V94 V142 1.6432667458492667e-12
C94_142 V94 V142 1.8570211195730782e-19

R94_143 V94 V143 -1289.3889402457582
L94_143 V94 V143 -2.183909959077593e-12
C94_143 V94 V143 -3.0834954537183386e-19

R94_144 V94 V144 -684.2789724410719
L94_144 V94 V144 -2.94523693397932e-11
C94_144 V94 V144 -5.308919385828051e-20

R94_145 V94 V145 -146.44058726337096
L94_145 V94 V145 -2.194568613918449e-12
C94_145 V94 V145 -2.060700272065403e-19

R94_146 V94 V146 -146.1839495063117
L94_146 V94 V146 -1.034677494605861e-12
C94_146 V94 V146 -1.1057531729795706e-19

R94_147 V94 V147 -316.01242800894477
L94_147 V94 V147 8.771548012700078e-12
C94_147 V94 V147 1.0589288097095468e-19

R94_148 V94 V148 -515.242806535229
L94_148 V94 V148 -5.9528367294159575e-12
C94_148 V94 V148 -6.075540518161757e-20

R94_149 V94 V149 2398.0404339027923
L94_149 V94 V149 4.798634094702967e-13
C94_149 V94 V149 1.2526723572147516e-18

R94_150 V94 V150 133.8434613969361
L94_150 V94 V150 2.9274884712894402e-12
C94_150 V94 V150 -6.302736460509683e-19

R94_151 V94 V151 616.2529547506624
L94_151 V94 V151 5.514002221196961e-12
C94_151 V94 V151 1.5883027227844213e-19

R94_152 V94 V152 -677.3499944683545
L94_152 V94 V152 -1.562170966200411e-11
C94_152 V94 V152 -5.150125956229075e-20

R94_153 V94 V153 167.0549112086997
L94_153 V94 V153 6.114255941776054e-12
C94_153 V94 V153 -3.182286614481533e-20

R94_154 V94 V154 112.7523122535405
L94_154 V94 V154 9.417124554665934e-12
C94_154 V94 V154 5.587313997195114e-19

R94_155 V94 V155 1413.7322798117086
L94_155 V94 V155 3.047402357392372e-12
C94_155 V94 V155 2.1917197760064074e-19

R94_156 V94 V156 158.09602232693666
L94_156 V94 V156 3.374062775886895e-12
C94_156 V94 V156 1.6138426113678232e-19

R94_157 V94 V157 197.44024137954227
L94_157 V94 V157 -5.610719872506125e-13
C94_157 V94 V157 -1.2061632751521605e-18

R94_158 V94 V158 -84.078177535581
L94_158 V94 V158 6.162018293464846e-12
C94_158 V94 V158 -8.060942900001166e-20

R94_159 V94 V159 636.7219071258368
L94_159 V94 V159 5.46792499056685e-11
C94_159 V94 V159 -1.9774661837065382e-20

R94_160 V94 V160 1860.53478471725
L94_160 V94 V160 7.933343821561106e-12
C94_160 V94 V160 9.895621902007273e-20

R94_161 V94 V161 -161.76099868592416
L94_161 V94 V161 -3.1528086387483466e-12
C94_161 V94 V161 -2.154461089356615e-21

R94_162 V94 V162 -100.37193114289936
L94_162 V94 V162 3.339068529615717e-12
C94_162 V94 V162 2.1927279599655472e-20

R94_163 V94 V163 -275.78117066985334
L94_163 V94 V163 -1.313984767611033e-12
C94_163 V94 V163 -3.5174879650113295e-19

R94_164 V94 V164 -209.4174007054161
L94_164 V94 V164 -1.91112170577117e-12
C94_164 V94 V164 -7.397005669213304e-20

R94_165 V94 V165 -179.99384885669028
L94_165 V94 V165 7.884678973065903e-13
C94_165 V94 V165 7.516307699021105e-19

R94_166 V94 V166 54.66324122135769
L94_166 V94 V166 5.7001434602249144e-12
C94_166 V94 V166 -2.3743585780925057e-20

R94_167 V94 V167 -402.9552930764185
L94_167 V94 V167 1.142588761180488e-11
C94_167 V94 V167 2.6901579971336784e-20

R94_168 V94 V168 -192.9196780382798
L94_168 V94 V168 2.4674585922539972e-11
C94_168 V94 V168 -1.0258256878375792e-19

R94_169 V94 V169 171.81067135784627
L94_169 V94 V169 -1.804374683673119e-11
C94_169 V94 V169 -2.7825250239423577e-19

R94_170 V94 V170 -1350.118122472086
L94_170 V94 V170 -5.260818357528161e-12
C94_170 V94 V170 3.1902439391761057e-19

R94_171 V94 V171 310.18504399041205
L94_171 V94 V171 8.85088812923759e-13
C94_171 V94 V171 5.661076637471846e-19

R94_172 V94 V172 182.82052074076532
L94_172 V94 V172 1.3477492359828013e-12
C94_172 V94 V172 3.3246757198718445e-19

R94_173 V94 V173 1561.6582005169362
L94_173 V94 V173 -1.6623949325827176e-12
C94_173 V94 V173 -1.9839659169213268e-19

R94_174 V94 V174 -58.53100082868283
L94_174 V94 V174 -4.727896601066814e-12
C94_174 V94 V174 -4.133184081942958e-19

R94_175 V94 V175 675.4028899091508
L94_175 V94 V175 -5.124553801796371e-12
C94_175 V94 V175 -6.341110383698129e-20

R94_176 V94 V176 347.5837474212255
L94_176 V94 V176 -4.6927689808663716e-12
C94_176 V94 V176 -3.364086953852129e-20

R94_177 V94 V177 -319.28247931390587
L94_177 V94 V177 7.243717815382757e-12
C94_177 V94 V177 2.6919570111417635e-19

R94_178 V94 V178 230.1526318222968
L94_178 V94 V178 7.555197528406658e-12
C94_178 V94 V178 -1.841201778913763e-19

R94_179 V94 V179 -394.3084683487224
L94_179 V94 V179 -1.279744703130202e-12
C94_179 V94 V179 -4.930028837835393e-19

R94_180 V94 V180 -247.72220545701373
L94_180 V94 V180 -1.3419090667690385e-12
C94_180 V94 V180 -3.6394967931638644e-19

R94_181 V94 V181 565.0436833066751
L94_181 V94 V181 -9.212538842941648e-12
C94_181 V94 V181 -1.3710693844615072e-19

R94_182 V94 V182 116.24235079287362
L94_182 V94 V182 1.1436639774550673e-12
C94_182 V94 V182 3.689463136759304e-19

R94_183 V94 V183 641.8896454076898
L94_183 V94 V183 -4.523244272682855e-12
C94_183 V94 V183 -1.111744556619097e-19

R94_184 V94 V184 917.1180246077544
L94_184 V94 V184 8.759218163533433e-12
C94_184 V94 V184 6.600636956639766e-20

R94_185 V94 V185 515.4940014151028
L94_185 V94 V185 6.341614882394503e-12
C94_185 V94 V185 -9.309504251063602e-20

R94_186 V94 V186 -512.3924120445658
L94_186 V94 V186 -8.356230042874625e-12
C94_186 V94 V186 5.591005912161552e-20

R94_187 V94 V187 -789.9051414647986
L94_187 V94 V187 1.666882070669922e-12
C94_187 V94 V187 4.071650119073849e-19

R94_188 V94 V188 -771.7445176951198
L94_188 V94 V188 1.9257841759433953e-12
C94_188 V94 V188 3.0540084205792297e-19

R94_189 V94 V189 -951.0866759359445
L94_189 V94 V189 1.9001309098629276e-12
C94_189 V94 V189 3.736462874326659e-19

R94_190 V94 V190 -146.42974011353584
L94_190 V94 V190 -1.1170977091783384e-11
C94_190 V94 V190 -3.6095978931271277e-19

R94_191 V94 V191 -485.15053557043194
L94_191 V94 V191 1.1421574752257353e-12
C94_191 V94 V191 3.8522613588334873e-19

R94_192 V94 V192 -4121.807983707693
L94_192 V94 V192 1.9293362593083694e-12
C94_192 V94 V192 2.2560258184657588e-19

R94_193 V94 V193 -569.092609464251
L94_193 V94 V193 -1.751730775861502e-12
C94_193 V94 V193 -2.47156926369323e-19

R94_194 V94 V194 384.33017769603015
L94_194 V94 V194 -8.45999642338741e-12
C94_194 V94 V194 -1.5586995014123597e-19

R94_195 V94 V195 375.9551841184695
L94_195 V94 V195 -8.902988089634642e-13
C94_195 V94 V195 -7.012379873326401e-19

R94_196 V94 V196 675.3244739221502
L94_196 V94 V196 -8.473913644300141e-13
C94_196 V94 V196 -6.269112679080191e-19

R94_197 V94 V197 456.1774413700265
L94_197 V94 V197 -1.5984520269577144e-12
C94_197 V94 V197 -1.9610748379332076e-19

R94_198 V94 V198 171.4522922851536
L94_198 V94 V198 1.724411951097336e-11
C94_198 V94 V198 1.1464352915437873e-19

R94_199 V94 V199 771.2994615954449
L94_199 V94 V199 -1.4472773651485485e-12
C94_199 V94 V199 -3.4228428562089938e-19

R94_200 V94 V200 -4701.876014601496
L94_200 V94 V200 -2.2836281975240006e-12
C94_200 V94 V200 -3.850195850066039e-20

R95_95 V95 0 -239.86712522310185
L95_95 V95 0 -1.0430949455076732e-12
C95_95 V95 0 3.317814078397769e-19

R95_96 V95 V96 -544.736234573175
L95_96 V95 V96 -6.536133693794451e-12
C95_96 V95 V96 -1.2030876648563726e-19

R95_97 V95 V97 -692.9913768352811
L95_97 V95 V97 -2.594899438850186e-12
C95_97 V95 V97 -4.005858426698056e-19

R95_98 V95 V98 5381.329206316946
L95_98 V95 V98 -1.5412657659315068e-11
C95_98 V95 V98 -2.0229861789018672e-19

R95_99 V95 V99 126.98590096445922
L95_99 V95 V99 2.6734136942250585e-12
C95_99 V95 V99 4.612192614367738e-19

R95_100 V95 V100 493.50836792982153
L95_100 V95 V100 4.337244100101746e-11
C95_100 V95 V100 8.568828288002025e-20

R95_101 V95 V101 -618.3331925088038
L95_101 V95 V101 3.3233679098291734e-12
C95_101 V95 V101 3.9812009049634217e-19

R95_102 V95 V102 635.7398347077516
L95_102 V95 V102 -1.756774488172653e-11
C95_102 V95 V102 3.2282352592573945e-20

R95_103 V95 V103 991.3129833071744
L95_103 V95 V103 1.970353992294435e-12
C95_103 V95 V103 2.508964979194362e-19

R95_104 V95 V104 964.3639734901202
L95_104 V95 V104 -2.8853246468742453e-11
C95_104 V95 V104 -4.4907795905239187e-20

R95_105 V95 V105 317.38912898235503
L95_105 V95 V105 4.7781052591153504e-12
C95_105 V95 V105 1.0352528345885923e-19

R95_106 V95 V106 -2867.9886238363247
L95_106 V95 V106 5.507250376004635e-12
C95_106 V95 V106 2.3996104252540995e-19

R95_107 V95 V107 -148.39084779307763
L95_107 V95 V107 -1.90171943681335e-12
C95_107 V95 V107 -3.938604657356262e-19

R95_108 V95 V108 -687.5142074914993
L95_108 V95 V108 5.5312832297357125e-12
C95_108 V95 V108 1.2475016657701354e-19

R95_109 V95 V109 552.2609137491896
L95_109 V95 V109 1.6184083573905424e-10
C95_109 V95 V109 -1.9807766518671959e-19

R95_110 V95 V110 -810.139782476149
L95_110 V95 V110 -4.5105855447204915e-10
C95_110 V95 V110 -5.231347415246442e-20

R95_111 V95 V111 229.38509498601485
L95_111 V95 V111 -6.870651796233981e-12
C95_111 V95 V111 -1.9448374789415237e-19

R95_112 V95 V112 1531.2995708173466
L95_112 V95 V112 1.0495133939448416e-11
C95_112 V95 V112 5.518571046395338e-20

R95_113 V95 V113 -181.8192120758322
L95_113 V95 V113 -4.587922169162471e-12
C95_113 V95 V113 -1.1844241934415173e-19

R95_114 V95 V114 -238216.8208721632
L95_114 V95 V114 -4.915149393085585e-12
C95_114 V95 V114 -2.8647773414307224e-19

R95_115 V95 V115 468.9851891510002
L95_115 V95 V115 3.6181004121568238e-12
C95_115 V95 V115 3.357094263296925e-19

R95_116 V95 V116 1946.7663881659676
L95_116 V95 V116 -4.432472897898872e-12
C95_116 V95 V116 -2.3115318361243174e-19

R95_117 V95 V117 -493.35232218617386
L95_117 V95 V117 -5.600036263025817e-12
C95_117 V95 V117 1.7141993639927345e-22

R95_118 V95 V118 1065.5667262442946
L95_118 V95 V118 1.1830029246720394e-11
C95_118 V95 V118 1.6959368021916995e-19

R95_119 V95 V119 -224.7140358367212
L95_119 V95 V119 1.1910440626733772e-10
C95_119 V95 V119 1.4349779696063425e-19

R95_120 V95 V120 -4845.315775308867
L95_120 V95 V120 7.555990187791322e-11
C95_120 V95 V120 1.5244369133141023e-19

R95_121 V95 V121 168.359092621788
L95_121 V95 V121 3.748134967831366e-12
C95_121 V95 V121 1.550715189471114e-19

R95_122 V95 V122 7315.881847617275
L95_122 V95 V122 4.945761865570847e-11
C95_122 V95 V122 4.570822321984346e-20

R95_123 V95 V123 277.521339896451
L95_123 V95 V123 -4.8719588364536055e-12
C95_123 V95 V123 -4.894894452814592e-19

R95_124 V95 V124 2983.7226392428497
L95_124 V95 V124 7.68793316231745e-12
C95_124 V95 V124 4.620303804769291e-20

R95_125 V95 V125 379.24085592657093
L95_125 V95 V125 4.124810257613321e-12
C95_125 V95 V125 1.1171034813658065e-19

R95_126 V95 V126 -2404.146172265525
L95_126 V95 V126 5.407784016140113e-11
C95_126 V95 V126 -6.12426304878945e-20

R95_127 V95 V127 1504.734053567047
L95_127 V95 V127 -1.3605835310046275e-11
C95_127 V95 V127 1.1805268619030262e-19

R95_128 V95 V128 -6825.927355873119
L95_128 V95 V128 2.1299226206914884e-11
C95_128 V95 V128 -5.1494196267424196e-20

R95_129 V95 V129 -135.09417040449102
L95_129 V95 V129 -4.416873669158807e-12
C95_129 V95 V129 -2.2478608106510196e-19

R95_130 V95 V130 -937.057102678811
L95_130 V95 V130 1.13894430587555e-10
C95_130 V95 V130 2.908629698616412e-20

R95_131 V95 V131 -357.7820648984019
L95_131 V95 V131 1.2857235507962116e-11
C95_131 V95 V131 1.6122110368345365e-19

R95_132 V95 V132 -1771.613465372057
L95_132 V95 V132 -1.2198608996699768e-11
C95_132 V95 V132 6.536512378926996e-20

R95_133 V95 V133 -680.7310854643854
L95_133 V95 V133 -1.0540198167587149e-11
C95_133 V95 V133 3.6701791551477413e-20

R95_134 V95 V134 -3196.7983588869083
L95_134 V95 V134 -4.6786669639882475e-12
C95_134 V95 V134 -8.354479904732138e-20

R95_135 V95 V135 186.41189662562502
L95_135 V95 V135 3.426920644555347e-12
C95_135 V95 V135 -2.4777477623822634e-19

R95_136 V95 V136 2718.157832326737
L95_136 V95 V136 -3.403364064317657e-11
C95_136 V95 V136 -4.6915650177115935e-20

R95_137 V95 V137 137.60681250137517
L95_137 V95 V137 4.576356877449775e-11
C95_137 V95 V137 1.0044801375753414e-20

R95_138 V95 V138 896.6523117696445
L95_138 V95 V138 6.825999828202488e-12
C95_138 V95 V138 2.5082274921614094e-21

R95_139 V95 V139 -234.87659568637065
L95_139 V95 V139 -4.276413944834853e-12
C95_139 V95 V139 3.10270912365388e-19

R95_140 V95 V140 -3088.420930771192
L95_140 V95 V140 -3.1391805813419916e-11
C95_140 V95 V140 1.118812642602799e-21

R95_141 V95 V141 443.2427780762889
L95_141 V95 V141 1.0783044411477672e-11
C95_141 V95 V141 -7.376461418586329e-20

R95_142 V95 V142 -28567.14448129368
L95_142 V95 V142 4.620130243091956e-12
C95_142 V95 V142 8.44259217528803e-20

R95_143 V95 V143 -225.11084378505404
L95_143 V95 V143 -2.519026763797273e-12
C95_143 V95 V143 -1.424134444872447e-19

R95_144 V95 V144 -2413.610932840496
L95_144 V95 V144 4.523600310345457e-11
C95_144 V95 V144 4.7848513685929757e-20

R95_145 V95 V145 -107.61671492863705
L95_145 V95 V145 2.4480181903011423e-11
C95_145 V95 V145 2.1133283603345924e-20

R95_146 V95 V146 -221.27218572782064
L95_146 V95 V146 -3.444566280274616e-12
C95_146 V95 V146 -3.3346828119335234e-20

R95_147 V95 V147 540.2012447423162
L95_147 V95 V147 1.4676627139759335e-12
C95_147 V95 V147 -1.2135987973890856e-19

R95_148 V95 V148 -368.14030936182485
L95_148 V95 V148 -5.413448939987078e-11
C95_148 V95 V148 -1.3576483293250882e-20

R95_149 V95 V149 -195255.0059849525
L95_149 V95 V149 8.650358009350277e-12
C95_149 V95 V149 3.409420777885132e-19

R95_150 V95 V150 240.75511962502114
L95_150 V95 V150 1.1354431257933758e-11
C95_150 V95 V150 -1.2396467381898516e-19

R95_151 V95 V151 63.052276047402
L95_151 V95 V151 3.5985845365512364e-12
C95_151 V95 V151 1.4882857797669361e-19

R95_152 V95 V152 511.3946186791942
L95_152 V95 V152 -8.542620682385712e-11
C95_152 V95 V152 -2.1426543828075963e-20

R95_153 V95 V153 189.20744295825781
L95_153 V95 V153 -1.1678214176248645e-11
C95_153 V95 V153 -1.839526997371168e-19

R95_154 V95 V154 196.68953332558988
L95_154 V95 V154 -2.0250162996987284e-11
C95_154 V95 V154 5.2239565503451365e-20

R95_155 V95 V155 -55.845987643187826
L95_155 V95 V155 -2.3455913177168357e-12
C95_155 V95 V155 1.5801420844219567e-19

R95_156 V95 V156 509.064737225811
L95_156 V95 V156 8.775361954535926e-12
C95_156 V95 V156 -3.917043975186064e-21

R95_157 V95 V157 179.7770024743876
L95_157 V95 V157 -4.018658053712081e-12
C95_157 V95 V157 -3.6808874847694315e-19

R95_158 V95 V158 -591.5337745686613
L95_158 V95 V158 6.227599349232016e-12
C95_158 V95 V158 5.1433160462649305e-20

R95_159 V95 V159 -173.94309452344936
L95_159 V95 V159 -3.347537679766344e-12
C95_159 V95 V159 -1.7865956730667715e-19

R95_160 V95 V160 -37281.30980646091
L95_160 V95 V160 -6.567750894287865e-12
C95_160 V95 V160 -1.458161775196856e-20

R95_161 V95 V161 -277.947193897712
L95_161 V95 V161 1.0503397492677674e-11
C95_161 V95 V161 1.7415763167266754e-19

R95_162 V95 V162 -299.15001700469065
L95_162 V95 V162 -1.5505640462746836e-11
C95_162 V95 V162 -1.9973361777468125e-20

R95_163 V95 V163 363.0653721739844
L95_163 V95 V163 2.0876939661546643e-12
C95_163 V95 V163 -5.3282270285558513e-20

R95_164 V95 V164 -1255.9722472312012
L95_164 V95 V164 -3.6848249830054637e-11
C95_164 V95 V164 1.56427279355661e-20

R95_165 V95 V165 -229.86229350392532
L95_165 V95 V165 2.013295653507159e-12
C95_165 V95 V165 2.4392309317494905e-19

R95_166 V95 V166 465.6336303033273
L95_166 V95 V166 5.562194968533976e-12
C95_166 V95 V166 1.8830722748289763e-20

R95_167 V95 V167 97.31500516634188
L95_167 V95 V167 -4.533076644252647e-12
C95_167 V95 V167 6.815596768804821e-20

R95_168 V95 V168 -279.2258151493122
L95_168 V95 V168 3.38847101337994e-12
C95_168 V95 V168 1.186892791855769e-19

R95_169 V95 V169 366.00388738849665
L95_169 V95 V169 -5.044522059415989e-12
C95_169 V95 V169 -2.4916893376032278e-19

R95_170 V95 V170 -3833.19414810147
L95_170 V95 V170 5.7665430703050686e-12
C95_170 V95 V170 1.315947945881424e-19

R95_171 V95 V171 -153.1817101145647
L95_171 V95 V171 9.770019582585135e-12
C95_171 V95 V171 1.2946377034675233e-19

R95_172 V95 V172 1563.7096245802795
L95_172 V95 V172 1.6268374664192878e-11
C95_172 V95 V172 1.7681622148609266e-20

R95_173 V95 V173 497.3777795769488
L95_173 V95 V173 -3.667850793424514e-12
C95_173 V95 V173 -9.736198219036816e-20

R95_174 V95 V174 -1201.5025803377068
L95_174 V95 V174 -2.051356125634669e-12
C95_174 V95 V174 -2.620406664455629e-19

R95_175 V95 V175 -331.5145974040152
L95_175 V95 V175 2.9681158105440684e-11
C95_175 V95 V175 6.412026695869783e-20

R95_176 V95 V176 1460.0625276691903
L95_176 V95 V176 -3.508092148975308e-12
C95_176 V95 V176 -1.3743759092072165e-19

R95_177 V95 V177 -2352.5835520340083
L95_177 V95 V177 1.575634646962113e-11
C95_177 V95 V177 1.2321858228082448e-19

R95_178 V95 V178 514.0145837276306
L95_178 V95 V178 5.7301316631058e-11
C95_178 V95 V178 -2.6945290455162048e-20

R95_179 V95 V179 -322.6644393081154
L95_179 V95 V179 2.124118609858072e-10
C95_179 V95 V179 -2.703225241690272e-19

R95_180 V95 V180 1912.8585176662716
L95_180 V95 V180 -1.6236133275402968e-11
C95_180 V95 V180 -6.911563661047034e-20

R95_181 V95 V181 -1468.8959304065954
L95_181 V95 V181 6.926760075631152e-12
C95_181 V95 V181 1.7944767817283412e-19

R95_182 V95 V182 -507.0319368746978
L95_182 V95 V182 2.598766684215497e-12
C95_182 V95 V182 1.6357511171337394e-19

R95_183 V95 V183 127.5727761251004
L95_183 V95 V183 -2.7954126460149936e-12
C95_183 V95 V183 -1.9021418779773336e-20

R95_184 V95 V184 15086.216565924691
L95_184 V95 V184 7.515847843026015e-12
C95_184 V95 V184 4.112723667062908e-20

R95_185 V95 V185 1180.6599357208274
L95_185 V95 V185 5.014823129610267e-12
C95_185 V95 V185 -1.7090765336135985e-19

R95_186 V95 V186 -963.9124866741938
L95_186 V95 V186 1.7284992326393605e-11
C95_186 V95 V186 3.0700786708754855e-20

R95_187 V95 V187 -911.23728008975
L95_187 V95 V187 2.910454443754933e-12
C95_187 V95 V187 2.9964319974617224e-19

R95_188 V95 V188 -499.3785808675231
L95_188 V95 V188 6.996046462034123e-12
C95_188 V95 V188 1.1976299287869948e-19

R95_189 V95 V189 4116.114822277213
L95_189 V95 V189 -4.486345857113208e-12
C95_189 V95 V189 -4.062068307744722e-20

R95_190 V95 V190 657.0977562579319
L95_190 V95 V190 -6.56992374756554e-12
C95_190 V95 V190 -1.0247058251549811e-19

R95_191 V95 V191 -188.79742007503685
L95_191 V95 V191 3.09147673320947e-12
C95_191 V95 V191 -6.363051995196871e-20

R95_192 V95 V192 8200.597138923174
L95_192 V95 V192 -8.849866775001431e-11
C95_192 V95 V192 -5.0888033071759756e-20

R95_193 V95 V193 -969.2416464034524
L95_193 V95 V193 -3.419240839909418e-12
C95_193 V95 V193 -6.177082866510518e-20

R95_194 V95 V194 6268.5607382659755
L95_194 V95 V194 -6.809394351305182e-12
C95_194 V95 V194 -1.8039031180362594e-19

R95_195 V95 V195 240.07847691115853
L95_195 V95 V195 -2.125382931945917e-12
C95_195 V95 V195 4.031091377239286e-20

R95_196 V95 V196 304.1911013263491
L95_196 V95 V196 -3.5288475326854127e-12
C95_196 V95 V196 -1.9422045788532454e-19

R95_197 V95 V197 683.0548481282343
L95_197 V95 V197 7.368830719447317e-12
C95_197 V95 V197 1.1395375160890486e-19

R95_198 V95 V198 2522.786256279914
L95_198 V95 V198 1.154917348289034e-11
C95_198 V95 V198 5.934067394878527e-20

R95_199 V95 V199 414.34480989280297
L95_199 V95 V199 -1.3719109850741603e-10
C95_199 V95 V199 -1.1062545451969054e-19

R95_200 V95 V200 -2568.766608423424
L95_200 V95 V200 -8.299960676293177e-11
C95_200 V95 V200 1.0362287213493452e-19

R96_96 V96 0 -57.51262666067581
L96_96 V96 0 -1.5371296970053174e-12
C96_96 V96 0 1.1390484516639257e-18

R96_97 V96 V97 -608.7036066025884
L96_97 V96 V97 -2.706871202270171e-12
C96_97 V96 V97 -5.048746708191949e-19

R96_98 V96 V98 882.8412518721497
L96_98 V96 V98 7.015008541466545e-12
C96_98 V96 V98 -2.480805434716396e-19

R96_99 V96 V99 410.4936554159196
L96_99 V96 V99 -1.8985278041981218e-11
C96_99 V96 V99 2.038979950594547e-19

R96_100 V96 V100 99.42551664918759
L96_100 V96 V100 -3.653897550311986e-11
C96_100 V96 V100 2.785451052569346e-19

R96_101 V96 V101 -749.2197471899829
L96_101 V96 V101 3.338575543461422e-12
C96_101 V96 V101 4.619336641503311e-19

R96_102 V96 V102 643.6780897875907
L96_102 V96 V102 -3.213323998568962e-11
C96_102 V96 V102 1.3905909631627944e-19

R96_103 V96 V103 790.3934522200137
L96_103 V96 V103 6.104961137874877e-11
C96_103 V96 V103 -6.195818399377415e-20

R96_104 V96 V104 599.6697194600326
L96_104 V96 V104 1.0958076479249304e-12
C96_104 V96 V104 3.543810138371652e-19

R96_105 V96 V105 336.6611529135476
L96_105 V96 V105 4.413833921074005e-12
C96_105 V96 V105 1.4313603124179685e-19

R96_106 V96 V106 -3892.460705850642
L96_106 V96 V106 7.798859852857903e-11
C96_106 V96 V106 1.802855553336487e-19

R96_107 V96 V107 -520.6856709463754
L96_107 V96 V107 -2.814411648903034e-11
C96_107 V96 V107 -1.034920177743537e-19

R96_108 V96 V108 -114.87701238951166
L96_108 V96 V108 -2.5010323049930153e-12
C96_108 V96 V108 -1.783725544187269e-19

R96_109 V96 V109 880.5192524066686
L96_109 V96 V109 5.643578807024802e-10
C96_109 V96 V109 -2.6342843059997186e-19

R96_110 V96 V110 -473.8198433833176
L96_110 V96 V110 4.670434521288981e-11
C96_110 V96 V110 -4.046816650560004e-20

R96_111 V96 V111 4205.481788304805
L96_111 V96 V111 5.271633004370696e-12
C96_111 V96 V111 1.1047354121487025e-19

R96_112 V96 V112 234.19772958875973
L96_112 V96 V112 -5.444317647232463e-12
C96_112 V96 V112 -3.919563140264487e-19

R96_113 V96 V113 -183.0244725978174
L96_113 V96 V113 -3.834267653353377e-12
C96_113 V96 V113 -1.817211381614063e-19

R96_114 V96 V114 5514.020062995687
L96_114 V96 V114 1.252688595691738e-09
C96_114 V96 V114 -2.67138105347064e-19

R96_115 V96 V115 15243.73746032041
L96_115 V96 V115 -2.4155777402596432e-11
C96_115 V96 V115 -3.875447033283065e-20

R96_116 V96 V116 269.53140083206154
L96_116 V96 V116 3.6845329185921624e-11
C96_116 V96 V116 1.9851402932303076e-19

R96_117 V96 V117 -461.767584804066
L96_117 V96 V117 -4.235914927793969e-12
C96_117 V96 V117 4.6264452552931765e-20

R96_118 V96 V118 356.21304610941115
L96_118 V96 V118 1.1013952248776425e-11
C96_118 V96 V118 2.1554525298790318e-19

R96_119 V96 V119 1212.2787594175225
L96_119 V96 V119 -9.115766844362787e-12
C96_119 V96 V119 8.119794203756287e-20

R96_120 V96 V120 -244.75940565456577
L96_120 V96 V120 1.7090257424974207e-11
C96_120 V96 V120 2.8983363369149583e-19

R96_121 V96 V121 182.44988928351805
L96_121 V96 V121 2.564653707407824e-12
C96_121 V96 V121 2.1129813494275052e-19

R96_122 V96 V122 -715.6062494535968
L96_122 V96 V122 -8.831233180549015e-12
C96_122 V96 V122 -7.854338949644512e-21

R96_123 V96 V123 -1654.222330919793
L96_123 V96 V123 8.13355244931769e-12
C96_123 V96 V123 -3.3484122373850356e-20

R96_124 V96 V124 562.0527052998168
L96_124 V96 V124 4.692728416932701e-12
C96_124 V96 V124 -4.753892959534966e-19

R96_125 V96 V125 391.6729269638033
L96_125 V96 V125 3.3282162065144673e-12
C96_125 V96 V125 6.224315782041258e-20

R96_126 V96 V126 -547.3948823878713
L96_126 V96 V126 6.480222411395939e-12
C96_126 V96 V126 -6.089962900975828e-20

R96_127 V96 V127 -464.2591820954833
L96_127 V96 V127 6.080884495207893e-12
C96_127 V96 V127 -3.70299453926264e-20

R96_128 V96 V128 3266.189199303088
L96_128 V96 V128 -3.0182332325733337e-12
C96_128 V96 V128 3.08746820406148e-20

R96_129 V96 V129 -120.82190444697639
L96_129 V96 V129 -2.307412090578661e-12
C96_129 V96 V129 -3.1629952013182665e-19

R96_130 V96 V130 1879.2379153557551
L96_130 V96 V130 1.1479119994472811e-11
C96_130 V96 V130 1.33405892836394e-19

R96_131 V96 V131 322.98819861943014
L96_131 V96 V131 -5.93203196306235e-12
C96_131 V96 V131 2.4222297256741156e-20

R96_132 V96 V132 -1039.550539771875
L96_132 V96 V132 -9.087398838613904e-12
C96_132 V96 V132 2.0720452891438592e-19

R96_133 V96 V133 -1583.7304645027987
L96_133 V96 V133 4.0581186567457045e-11
C96_133 V96 V133 1.7330085610895262e-19

R96_134 V96 V134 1951.2790686003245
L96_134 V96 V134 -2.6717323232632177e-12
C96_134 V96 V134 -1.741319048533143e-19

R96_135 V96 V135 -2917.7239909964815
L96_135 V96 V135 2.438329503623068e-11
C96_135 V96 V135 3.5879715533771e-20

R96_136 V96 V136 276.53272657191405
L96_136 V96 V136 1.4748979613722309e-12
C96_136 V96 V136 -2.131903271545999e-19

R96_137 V96 V137 137.97716325578781
L96_137 V96 V137 7.61663221314364e-12
C96_137 V96 V137 3.7945725310491666e-20

R96_138 V96 V138 -1923.5919468883458
L96_138 V96 V138 3.30814527781296e-12
C96_138 V96 V138 7.546292010005976e-20

R96_139 V96 V139 -466.8249017742071
L96_139 V96 V139 6.564495084235893e-12
C96_139 V96 V139 9.446231932978342e-20

R96_140 V96 V140 -969.9143627606791
L96_140 V96 V140 -1.537567359175746e-12
C96_140 V96 V140 1.2689720168043493e-19

R96_141 V96 V141 545.2600587443231
L96_141 V96 V141 1.0353955353440846e-11
C96_141 V96 V141 -2.192801433388506e-19

R96_142 V96 V142 -1400.1980257872237
L96_142 V96 V142 2.7714566473397355e-12
C96_142 V96 V142 1.0975425345581532e-19

R96_143 V96 V143 991.662373324513
L96_143 V96 V143 -7.233687118339426e-12
C96_143 V96 V143 -1.780796158155018e-19

R96_144 V96 V144 -100.1317541996777
L96_144 V96 V144 -8.12764515083382e-12
C96_144 V96 V144 2.7806856031545406e-20

R96_145 V96 V145 -99.34628640668745
L96_145 V96 V145 -1.6313231994268085e-11
C96_145 V96 V145 -8.120818170229285e-22

R96_146 V96 V146 -206.91065444503099
L96_146 V96 V146 -1.8504458978224572e-12
C96_146 V96 V146 -7.249732230393575e-20

R96_147 V96 V147 -306.9787618685584
L96_147 V96 V147 2.449259327159168e-11
C96_147 V96 V147 -6.54548789422662e-21

R96_148 V96 V148 75.57934469291743
L96_148 V96 V148 9.776167162803438e-13
C96_148 V96 V148 -5.865828016954396e-20

R96_149 V96 V149 9802.189469241906
L96_149 V96 V149 3.852171134868175e-12
C96_149 V96 V149 5.313251585674201e-19

R96_150 V96 V150 159.06764968341074
L96_150 V96 V150 5.7434963940916305e-12
C96_150 V96 V150 -2.8714849103200208e-19

R96_151 V96 V151 359.544074703164
L96_151 V96 V151 4.8642325806632214e-12
C96_151 V96 V151 1.533096215449253e-19

R96_152 V96 V152 255.3948469159894
L96_152 V96 V152 -4.466574832411926e-11
C96_152 V96 V152 -5.1571525870538346e-20

R96_153 V96 V153 178.56661071066821
L96_153 V96 V153 -6.596180329359599e-12
C96_153 V96 V153 -1.6294454951860336e-19

R96_154 V96 V154 290.62178067571506
L96_154 V96 V154 -2.0744565773715583e-11
C96_154 V96 V154 1.864947100316456e-19

R96_155 V96 V155 -531.0639201354797
L96_155 V96 V155 -7.33189989474242e-11
C96_155 V96 V155 1.0524829734876232e-19

R96_156 V96 V156 445.1180129191135
L96_156 V96 V156 -1.109431956897663e-12
C96_156 V96 V156 9.009637063584089e-20

R96_157 V96 V157 133.94316174222828
L96_157 V96 V157 -2.476224105907257e-12
C96_157 V96 V157 -6.401336605560694e-19

R96_158 V96 V158 -5081.995029114685
L96_158 V96 V158 6.9786424811214084e-12
C96_158 V96 V158 1.3035211977978227e-20

R96_159 V96 V159 201.62220901607614
L96_159 V96 V159 -4.017143480168855e-12
C96_159 V96 V159 -1.2399016188378797e-19

R96_160 V96 V160 -59.25285273452453
L96_160 V96 V160 -2.7985371687813105e-11
C96_160 V96 V160 2.904023762425341e-20

R96_161 V96 V161 -198.46803874383616
L96_161 V96 V161 -6.484762801330228e-12
C96_161 V96 V161 1.6598612097152854e-19

R96_162 V96 V162 -227.2473539189789
L96_162 V96 V162 -4.387906709341499e-12
C96_162 V96 V162 -3.73486623635261e-20

R96_163 V96 V163 -422.8420178079177
L96_163 V96 V163 -2.3314797359805087e-12
C96_163 V96 V163 -1.8990567211993425e-19

R96_164 V96 V164 120.64280754919652
L96_164 V96 V164 2.183397465723e-12
C96_164 V96 V164 -7.177235402387259e-21

R96_165 V96 V165 -343.3046088855737
L96_165 V96 V165 1.2061883564518448e-12
C96_165 V96 V165 3.8948823680757544e-19

R96_166 V96 V166 248.58025496176177
L96_166 V96 V166 3.068740366465113e-12
C96_166 V96 V166 -7.831077858287183e-21

R96_167 V96 V167 520.4890273001893
L96_167 V96 V167 2.9246252700079435e-12
C96_167 V96 V167 1.158297591790614e-19

R96_168 V96 V168 599.7612379090344
L96_168 V96 V168 -3.4931804152139858e-12
C96_168 V96 V168 5.442273888002534e-20

R96_169 V96 V169 301.1621179063449
L96_169 V96 V169 -5.0323018062442985e-12
C96_169 V96 V169 -2.8506512601759976e-19

R96_170 V96 V170 1302.9271304491879
L96_170 V96 V170 1.542789779742671e-11
C96_170 V96 V170 1.9694960423787143e-19

R96_171 V96 V171 -1243.4573299761807
L96_171 V96 V171 2.7262946584393186e-12
C96_171 V96 V171 2.5740368461951745e-19

R96_172 V96 V172 -1424.6870806954644
L96_172 V96 V172 3.406036146668451e-12
C96_172 V96 V172 1.1509363338569773e-19

R96_173 V96 V173 669.0368437208414
L96_173 V96 V173 -1.979844491163606e-12
C96_173 V96 V173 -1.587030414853123e-19

R96_174 V96 V174 -343.46094248826427
L96_174 V96 V174 -2.0715865522768967e-12
C96_174 V96 V174 -3.2567313226336404e-19

R96_175 V96 V175 903.6582476207004
L96_175 V96 V175 -3.917843615467897e-12
C96_175 V96 V175 -9.812342813485541e-20

R96_176 V96 V176 -356.7800093002738
L96_176 V96 V176 -2.430563873653675e-12
C96_176 V96 V176 -3.1546178739857666e-20

R96_177 V96 V177 -25279.275300223293
L96_177 V96 V177 7.632141928935364e-12
C96_177 V96 V177 1.5894305101229e-19

R96_178 V96 V178 891.528826404969
L96_178 V96 V178 1.693532203554899e-11
C96_178 V96 V178 -6.898651043950626e-20

R96_179 V96 V179 -1619.1890346609653
L96_179 V96 V179 -4.3315936961252164e-12
C96_179 V96 V179 -2.424207653231034e-19

R96_180 V96 V180 -245.6011532310549
L96_180 V96 V180 4.098137275090375e-12
C96_180 V96 V180 -2.3778312382553586e-19

R96_181 V96 V181 -1466.3267981250876
L96_181 V96 V181 6.771380211350826e-12
C96_181 V96 V181 1.6708765110752758e-19

R96_182 V96 V182 -5113.714741079024
L96_182 V96 V182 1.9524361946112603e-12
C96_182 V96 V182 2.1924468775096466e-19

R96_183 V96 V183 69270.55153738588
L96_183 V96 V183 8.391715803235507e-12
C96_183 V96 V183 -4.14944553210611e-20

R96_184 V96 V184 153.110422692334
L96_184 V96 V184 -6.738922475483205e-12
C96_184 V96 V184 5.369648490257143e-20

R96_185 V96 V185 845.1885501534691
L96_185 V96 V185 5.253251985228863e-12
C96_185 V96 V185 -1.917128032310831e-19

R96_186 V96 V186 2795.842907272441
L96_186 V96 V186 1.0699141477414726e-11
C96_186 V96 V186 5.642559197276369e-20

R96_187 V96 V187 -1104.806855655255
L96_187 V96 V187 4.74860906783548e-12
C96_187 V96 V187 2.061505924987109e-19

R96_188 V96 V188 -362.73214849551397
L96_188 V96 V188 1.1316552554071533e-11
C96_188 V96 V188 3.2034898901367573e-19

R96_189 V96 V189 2794.7335549028676
L96_189 V96 V189 -7.248476067964569e-12
C96_189 V96 V189 4.061075960349695e-20

R96_190 V96 V190 1321.994180863888
L96_190 V96 V190 -3.5482554025396035e-12
C96_190 V96 V190 -1.8737652054104114e-19

R96_191 V96 V191 9145.907228111955
L96_191 V96 V191 6.7727493111022625e-12
C96_191 V96 V191 1.3576932494519152e-19

R96_192 V96 V192 -195.11475070934176
L96_192 V96 V192 2.7973652499099338e-12
C96_192 V96 V192 -1.3701033032463236e-19

R96_193 V96 V193 -365.5866666530086
L96_193 V96 V193 -2.9102898203795707e-12
C96_193 V96 V193 -1.233332887126514e-19

R96_194 V96 V194 1566.2540728512033
L96_194 V96 V194 -1.8525698075455765e-11
C96_194 V96 V194 -2.2904780470598945e-19

R96_195 V96 V195 674.6447268421792
L96_195 V96 V195 -9.262615757915551e-12
C96_195 V96 V195 -3.1306742409531997e-19

R96_196 V96 V196 154.1719617091459
L96_196 V96 V196 -8.672718166225594e-13
C96_196 V96 V196 -1.1137714059729126e-19

R96_197 V96 V197 1733.498651847698
L96_197 V96 V197 3.393929534292742e-11
C96_197 V96 V197 7.708516399024721e-20

R96_198 V96 V198 403.78243412014945
L96_198 V96 V198 3.4247965431099936e-11
C96_198 V96 V198 2.994799921990581e-20

R96_199 V96 V199 221.65548012996527
L96_199 V96 V199 -1.9395731151924052e-12
C96_199 V96 V199 -1.9195092108516917e-19

R96_200 V96 V200 -1135.5729089777099
L96_200 V96 V200 2.9327017212591936e-12
C96_200 V96 V200 9.697564492853893e-20

R97_97 V97 0 -349.2986716341752
L97_97 V97 0 5.115738130770007e-13
C97_97 V97 0 2.6515429675002784e-18

R97_98 V97 V98 -5703.921079201165
L97_98 V97 V98 -1.047125122049778e-12
C97_98 V97 V98 -7.933617768624719e-19

R97_99 V97 V99 505.10117885388485
L97_99 V97 V99 5.817743892876556e-13
C97_99 V97 V99 1.1103486066270527e-18

R97_100 V97 V100 325.650346427998
L97_100 V97 V100 9.505679396769791e-13
C97_100 V97 V100 1.0065717741331017e-18

R97_101 V97 V101 -653.2469197747758
L97_101 V97 V101 7.602333670641724e-13
C97_101 V97 V101 1.061120627405857e-18

R97_102 V97 V102 1924.519304933283
L97_102 V97 V102 1.404991236032626e-12
C97_102 V97 V102 4.903808695630664e-19

R97_103 V97 V103 5546.2434074543735
L97_103 V97 V103 -2.1653454630856197e-12
C97_103 V97 V103 -2.910423990993347e-19

R97_104 V97 V104 7091.391491293395
L97_104 V97 V104 -1.7907762540616043e-12
C97_104 V97 V104 -3.4038925752468387e-19

R97_105 V97 V105 219.31771209294772
L97_105 V97 V105 7.790713518093984e-13
C97_105 V97 V105 5.758232766829011e-19

R97_106 V97 V106 652.1417971118124
L97_106 V97 V106 1.2449093353348004e-12
C97_106 V97 V106 7.140133424189312e-19

R97_107 V97 V107 -687.0584759444791
L97_107 V97 V107 -1.0941370828537141e-12
C97_107 V97 V107 -5.399995474540574e-19

R97_108 V97 V108 -439.4145345422248
L97_108 V97 V108 4.9185643067785085e-12
C97_108 V97 V108 3.9969012036961716e-20

R97_109 V97 V109 -1060.2835946028194
L97_109 V97 V109 -1.0319889656956517e-12
C97_109 V97 V109 -8.149854227679593e-19

R97_110 V97 V110 -583.0297149008662
L97_110 V97 V110 -1.8450211103859953e-12
C97_110 V97 V110 -4.801046357923801e-19

R97_111 V97 V111 645.780119639374
L97_111 V97 V111 4.348421647623983e-12
C97_111 V97 V111 1.5151860474483223e-19

R97_112 V97 V112 593.0163272162488
L97_112 V97 V112 -2.5030990417219807e-12
C97_112 V97 V112 -3.275986539647447e-19

R97_113 V97 V113 -197.81554471104397
L97_113 V97 V113 -2.4420882693190697e-12
C97_113 V97 V113 -1.5207290645722138e-19

R97_114 V97 V114 -790.7914815376148
L97_114 V97 V114 -9.653591321263835e-13
C97_114 V97 V114 -7.444907127036018e-19

R97_115 V97 V115 -3538.9945532038655
L97_115 V97 V115 1.1851638465087927e-12
C97_115 V97 V115 2.745596389082608e-19

R97_116 V97 V116 1908.6006667012632
L97_116 V97 V116 2.146361322340467e-12
C97_116 V97 V116 1.948001073499235e-20

R97_117 V97 V117 495.41791879798797
L97_117 V97 V117 4.13505305100234e-11
C97_117 V97 V117 -9.580177291141311e-20

R97_118 V97 V118 317.06891744092815
L97_118 V97 V118 7.827899856035003e-13
C97_118 V97 V118 9.093503498825893e-19

R97_119 V97 V119 -10174.388946561643
L97_119 V97 V119 1.258017040061572e-11
C97_119 V97 V119 3.2953945843661443e-19

R97_120 V97 V120 -1006.4376736892633
L97_120 V97 V120 1.969970750731995e-12
C97_120 V97 V120 7.71753670337326e-19

R97_121 V97 V121 585.3427944697906
L97_121 V97 V121 3.231211475963416e-12
C97_121 V97 V121 4.906114654788126e-19

R97_122 V97 V122 -1400.3590898486134
L97_122 V97 V122 -5.426309419318867e-12
C97_122 V97 V122 -4.370493620164478e-20

R97_123 V97 V123 1166.232941830603
L97_123 V97 V123 -9.765602767472254e-13
C97_123 V97 V123 -6.861560180184326e-19

R97_124 V97 V124 905.6754703557501
L97_124 V97 V124 -6.722514159034827e-13
C97_124 V97 V124 -1.1192842219906714e-18

R97_125 V97 V125 -2973.2179790542577
L97_125 V97 V125 2.298525206369116e-12
C97_125 V97 V125 1.4915320772238724e-19

R97_126 V97 V126 -525.3991583290232
L97_126 V97 V126 -9.4621108809556e-13
C97_126 V97 V126 -4.472398618103682e-19

R97_127 V97 V127 -641.2054365271509
L97_127 V97 V127 1.8088420039440858e-11
C97_127 V97 V127 -8.347747907901756e-21

R97_128 V97 V128 -1273.3928241389358
L97_128 V97 V128 2.2214902615174926e-12
C97_128 V97 V128 8.276521105618216e-20

R97_129 V97 V129 -526.4983122186218
L97_129 V97 V129 -1.0525530004858976e-12
C97_129 V97 V129 -8.470674515613431e-19

R97_130 V97 V130 1379.3960174054978
L97_130 V97 V130 1.222507332613608e-12
C97_130 V97 V130 3.466589746089281e-19

R97_131 V97 V131 707.5671409702409
L97_131 V97 V131 1.6063189871596816e-12
C97_131 V97 V131 4.633763104290807e-19

R97_132 V97 V132 1139.2748916252262
L97_132 V97 V132 1.2086624179286288e-12
C97_132 V97 V132 7.722690973955097e-19

R97_133 V97 V133 -1074.1176092091814
L97_133 V97 V133 1.4357748040977168e-12
C97_133 V97 V133 6.230868523163018e-19

R97_134 V97 V134 2708.529143831753
L97_134 V97 V134 -3.753022212212044e-12
C97_134 V97 V134 4.881543145905433e-20

R97_135 V97 V135 812.9538125169544
L97_135 V97 V135 -2.9164116310028156e-12
C97_135 V97 V135 -4.408178071338545e-19

R97_136 V97 V136 555.0101366871817
L97_136 V97 V136 -1.2889907940590333e-12
C97_136 V97 V136 -9.142341305577778e-19

R97_137 V97 V137 354.9784643981625
L97_137 V97 V137 4.4694772893776056e-12
C97_137 V97 V137 -3.439680413149204e-21

R97_138 V97 V138 -1947.673377526433
L97_138 V97 V138 -2.7644868842811344e-12
C97_138 V97 V138 -3.0104653260894203e-19

R97_139 V97 V139 -320.6644424455088
L97_139 V97 V139 1.7381504754822573e-12
C97_139 V97 V139 6.688937296042278e-19

R97_140 V97 V140 -297.87176888157904
L97_140 V97 V140 2.36766630135414e-12
C97_140 V97 V140 8.496737167981141e-19

R97_141 V97 V141 845.9720097652475
L97_141 V97 V141 -8.270606444379373e-13
C97_141 V97 V141 -7.250081806589057e-19

R97_142 V97 V142 -1049.5179668835126
L97_142 V97 V142 4.103114482446705e-12
C97_142 V97 V142 6.3629452628964e-20

R97_143 V97 V143 995.0014299655109
L97_143 V97 V143 -1.3054656610317058e-12
C97_143 V97 V143 -3.7793332122958036e-19

R97_144 V97 V144 -2039.7291971702737
L97_144 V97 V144 -1.121829032599095e-11
C97_144 V97 V144 -7.270366908793653e-20

R97_145 V97 V145 -274.6024995796697
L97_145 V97 V145 -1.1602640776601588e-10
C97_145 V97 V145 1.2257984189156865e-19

R97_146 V97 V146 1124.5423272486537
L97_146 V97 V146 1.782742312343432e-11
C97_146 V97 V146 1.6715988158398493e-19

R97_147 V97 V147 8405.75156223129
L97_147 V97 V147 -9.855533704755216e-12
C97_147 V97 V147 -5.204776975604857e-19

R97_148 V97 V148 310.61454244343867
L97_148 V97 V148 -1.3816257237567926e-12
C97_148 V97 V148 -5.588729809926306e-19

R97_149 V97 V149 2761.8803064401786
L97_149 V97 V149 4.708450228263243e-13
C97_149 V97 V149 1.075915288943397e-18

R97_150 V97 V150 507.65320594526577
L97_150 V97 V150 1.3596072806441292e-11
C97_150 V97 V150 -4.391504259690922e-19

R97_151 V97 V151 546.4196947411025
L97_151 V97 V151 1.9829652397400197e-12
C97_151 V97 V151 4.465640474882506e-19

R97_152 V97 V152 -1051.1738971352327
L97_152 V97 V152 1.8014302820542375e-12
C97_152 V97 V152 1.125782509770159e-19

R97_153 V97 V153 1249.6595727804065
L97_153 V97 V153 -3.2674028073633065e-12
C97_153 V97 V153 -3.544283121600751e-19

R97_154 V97 V154 -3862.8592191912517
L97_154 V97 V154 -9.370095962110728e-12
C97_154 V97 V154 1.1644183225930944e-19

R97_155 V97 V155 -226.85198692315342
L97_155 V97 V155 1.1429292365452193e-12
C97_155 V97 V155 4.396948845761308e-19

R97_156 V97 V156 955.6479360424368
L97_156 V97 V156 -7.882289087672824e-12
C97_156 V97 V156 4.243332758154326e-19

R97_157 V97 V157 518.7701443197155
L97_157 V97 V157 -4.625122001391744e-13
C97_157 V97 V157 -1.2187274232880145e-18

R97_158 V97 V158 8580.05435973348
L97_158 V97 V158 4.76559041420898e-12
C97_158 V97 V158 1.3093383507449953e-19

R97_159 V97 V159 375.40461344562016
L97_159 V97 V159 -1.291513843498301e-12
C97_159 V97 V159 -4.330718074107742e-19

R97_160 V97 V160 -874.6761298084672
L97_160 V97 V160 -3.5713784925566448e-12
C97_160 V97 V160 -2.487354446059539e-19

R97_161 V97 V161 -842.160297806265
L97_161 V97 V161 8.394624823193241e-13
C97_161 V97 V161 5.897028091089407e-19

R97_162 V97 V162 -928.1457224335496
L97_162 V97 V162 1.4603554094356317e-12
C97_162 V97 V162 1.127494204060293e-19

R97_163 V97 V163 -1151.8751477362862
L97_163 V97 V163 -4.786457744565186e-12
C97_163 V97 V163 -9.699199372750292e-20

R97_164 V97 V164 1759.45668511546
L97_164 V97 V164 -3.8146585511849216e-11
C97_164 V97 V164 2.55738766331341e-19

R97_165 V97 V165 -792.1581132470468
L97_165 V97 V165 2.7384433746686662e-12
C97_165 V97 V165 2.069915111975475e-19

R97_166 V97 V166 1044.6948239157289
L97_166 V97 V166 -5.952103331375946e-12
C97_166 V97 V166 -1.550252198052378e-19

R97_167 V97 V167 840.0653700038413
L97_167 V97 V167 2.7154121521534622e-12
C97_167 V97 V167 2.5632803050172193e-19

R97_168 V97 V168 -628.2435784707565
L97_168 V97 V168 1.257635357527143e-12
C97_168 V97 V168 1.7090583757806468e-19

R97_169 V97 V169 576.2103201951777
L97_169 V97 V169 -1.3346352410734026e-12
C97_169 V97 V169 -5.739398468740075e-19

R97_170 V97 V170 676.8815380229535
L97_170 V97 V170 2.7264253263004615e-12
C97_170 V97 V170 3.3398627795510905e-19

R97_171 V97 V171 -33740.669388061666
L97_171 V97 V171 1.2147473715043607e-12
C97_171 V97 V171 2.6351916340605186e-19

R97_172 V97 V172 669.4780836301228
L97_172 V97 V172 -3.432191385998956e-12
C97_172 V97 V172 -1.2425364482985508e-20

R97_173 V97 V173 2684.3544029169348
L97_173 V97 V173 2.3076090081069374e-12
C97_173 V97 V173 -1.536989182516031e-22

R97_174 V97 V174 -467.7820893162638
L97_174 V97 V174 -1.3056655648765819e-12
C97_174 V97 V174 -5.699076579226438e-19

R97_175 V97 V175 -3764.1007377318906
L97_175 V97 V175 -3.056987678874728e-12
C97_175 V97 V175 9.83922291517744e-20

R97_176 V97 V176 -2916.4098976933806
L97_176 V97 V176 -6.92526933268886e-12
C97_176 V97 V176 1.7921258561709588e-19

R97_177 V97 V177 -3049.54599745706
L97_177 V97 V177 -1.5568422715102532e-12
C97_177 V97 V177 1.8923109429592813e-19

R97_178 V97 V178 10109.791861962914
L97_178 V97 V178 -4.076213074623893e-12
C97_178 V97 V178 -9.669319210309796e-20

R97_179 V97 V179 -690.1124748316531
L97_179 V97 V179 -1.4799993848355553e-12
C97_179 V97 V179 -6.333763116530721e-19

R97_180 V97 V180 -532.6622427732051
L97_180 V97 V180 -2.1184569282604678e-12
C97_180 V97 V180 -5.5249410070469605e-19

R97_181 V97 V181 514.1598902889418
L97_181 V97 V181 8.851303721946204e-13
C97_181 V97 V181 2.490201042412086e-19

R97_182 V97 V182 1349.526258987037
L97_182 V97 V182 8.592928346748195e-13
C97_182 V97 V182 3.404608251996192e-19

R97_183 V97 V183 500.9769302108911
L97_183 V97 V183 -1.5253886821413968e-12
C97_183 V97 V183 -1.271417366548376e-19

R97_184 V97 V184 530.8982640886097
L97_184 V97 V184 -2.0094026587735762e-12
C97_184 V97 V184 8.451065324442407e-20

R97_185 V97 V185 -597.6219565431328
L97_185 V97 V185 4.160806971161694e-12
C97_185 V97 V185 -2.879185640856753e-19

R97_186 V97 V186 -4037.0757213851152
L97_186 V97 V186 -2.728059865012792e-12
C97_186 V97 V186 4.9155811605107344e-20

R97_187 V97 V187 -1049.951735662035
L97_187 V97 V187 1.0628669878417227e-12
C97_187 V97 V187 6.85509262731328e-19

R97_188 V97 V188 -705.0417144756648
L97_188 V97 V188 5.380081944379521e-13
C97_188 V97 V188 6.20316194211211e-19

R97_189 V97 V189 -2134.6469539572513
L97_189 V97 V189 -8.973651870749961e-13
C97_189 V97 V189 -6.037952739700282e-20

R97_190 V97 V190 7263.887005267208
L97_190 V97 V190 -3.832717297328181e-12
C97_190 V97 V190 -2.7251828471802044e-19

R97_191 V97 V191 -665.7019765678448
L97_191 V97 V191 9.215378149861471e-13
C97_191 V97 V191 5.50759868927739e-20

R97_192 V97 V192 -636.3468889194954
L97_192 V97 V192 -2.377110883712445e-12
C97_192 V97 V192 -4.04502830097937e-19

R97_193 V97 V193 904.7776161469994
L97_193 V97 V193 4.658038839628601e-12
C97_193 V97 V193 -1.588037294564069e-19

R97_194 V97 V194 -4661.82375722686
L97_194 V97 V194 -1.2922409497654795e-12
C97_194 V97 V194 -6.399461131659717e-19

R97_195 V97 V195 669.0918286113159
L97_195 V97 V195 -6.752494168244137e-13
C97_195 V97 V195 -4.272506885294636e-19

R97_196 V97 V196 381.1573944316804
L97_196 V97 V196 -1.1472360779044412e-12
C97_196 V97 V196 8.875353628567411e-20

R97_197 V97 V197 2190.5528372928275
L97_197 V97 V197 9.513633583794744e-12
C97_197 V97 V197 2.6036890552949766e-19

R97_198 V97 V198 962.5318772592461
L97_198 V97 V198 3.577606091294613e-12
C97_198 V97 V198 4.584277072564955e-20

R97_199 V97 V199 533.4399935092928
L97_199 V97 V199 -4.182711936656716e-12
C97_199 V97 V199 -1.7495602815298623e-19

R97_200 V97 V200 19298.898593178434
L97_200 V97 V200 3.407244847997773e-12
C97_200 V97 V200 1.7705208563529042e-19

R98_98 V98 0 209.21268012199823
L98_98 V98 0 3.05028574806482e-13
C98_98 V98 0 1.8638642126003832e-18

R98_99 V98 V99 -491.17740497928656
L98_99 V98 V99 5.732795789584607e-13
C98_99 V98 V99 9.126451370419761e-19

R98_100 V98 V100 4581.65710150657
L98_100 V98 V100 8.482856281623719e-13
C98_100 V98 V100 7.407132980654657e-19

R98_101 V98 V101 -441.8903186894313
L98_101 V98 V101 1.5506184949083146e-12
C98_101 V98 V101 4.9513640621687e-19

R98_102 V98 V102 1141.2467800322288
L98_102 V98 V102 1.1952217947903216e-12
C98_102 V98 V102 5.071469839217453e-19

R98_103 V98 V103 -560.5099624591171
L98_103 V98 V103 -1.0975523563889702e-12
C98_103 V98 V103 -3.096619587863899e-19

R98_104 V98 V104 -262.18666891476164
L98_104 V98 V104 -9.128530427282765e-13
C98_104 V98 V104 -3.4525047041943254e-19

R98_105 V98 V105 256.7913924079849
L98_105 V98 V105 5.914936531294546e-12
C98_105 V98 V105 8.519587540625292e-20

R98_106 V98 V106 1138.7120558708957
L98_106 V98 V106 6.914655451260603e-13
C98_106 V98 V106 6.302438739431243e-19

R98_107 V98 V107 620.713967226992
L98_107 V98 V107 -1.7446230311889983e-12
C98_107 V98 V107 -4.1262846078073213e-19

R98_108 V98 V108 1374.6179668483544
L98_108 V98 V108 3.76836362290292e-12
C98_108 V98 V108 -1.858573555136191e-20

R98_109 V98 V109 -10590.966636670375
L98_109 V98 V109 -2.177890174489425e-12
C98_109 V98 V109 -5.388158100431198e-19

R98_110 V98 V110 446.2558292519376
L98_110 V98 V110 -1.0492035503707987e-12
C98_110 V98 V110 -4.672640533134897e-19

R98_111 V98 V111 507.17545430124983
L98_111 V98 V111 3.797847731306714e-12
C98_111 V98 V111 9.512843743632419e-20

R98_112 V98 V112 340.36374322962473
L98_112 V98 V112 -4.122665004272657e-12
C98_112 V98 V112 -1.723543387691031e-19

R98_113 V98 V113 1107.9569818611449
L98_113 V98 V113 4.931866709560863e-12
C98_113 V98 V113 2.55988435620511e-19

R98_114 V98 V114 3320.8057907331604
L98_114 V98 V114 -9.977256543378583e-13
C98_114 V98 V114 -5.343453146300595e-19

R98_115 V98 V115 -412.45489410749224
L98_115 V98 V115 1.6305217482158221e-12
C98_115 V98 V115 2.5051438329492475e-19

R98_116 V98 V116 -636.3452068313219
L98_116 V98 V116 2.1345475800737096e-12
C98_116 V98 V116 1.0254950800617465e-19

R98_117 V98 V117 446.993708955447
L98_117 V98 V117 3.481689052046531e-12
C98_117 V98 V117 8.900089609406068e-20

R98_118 V98 V118 -126.72200556706393
L98_118 V98 V118 1.2767631778995761e-12
C98_118 V98 V118 6.131286828052823e-19

R98_119 V98 V119 -399.5438634156329
L98_119 V98 V119 1.0888613811377548e-11
C98_119 V98 V119 1.8951851963717995e-19

R98_120 V98 V120 -306.3109117987253
L98_120 V98 V120 2.4310569898003043e-12
C98_120 V98 V120 4.778559530839533e-19

R98_121 V98 V121 -409.67512271699724
L98_121 V98 V121 -3.2461351860397986e-12
C98_121 V98 V121 -2.0593094646237515e-19

R98_122 V98 V122 291.95069114473256
L98_122 V98 V122 2.8073761819016213e-12
C98_122 V98 V122 1.0721080502070348e-19

R98_123 V98 V123 351.4219680878535
L98_123 V98 V123 -1.0192014334708529e-12
C98_123 V98 V123 -4.987121825769841e-19

R98_124 V98 V124 288.54045777664027
L98_124 V98 V124 -6.537558063188002e-13
C98_124 V98 V124 -8.281726134362373e-19

R98_125 V98 V125 -9989.90988147195
L98_125 V98 V125 1.3489960548777589e-11
C98_125 V98 V125 1.525247195138237e-19

R98_126 V98 V126 138.61762159725694
L98_126 V98 V126 -8.492529887592369e-13
C98_126 V98 V126 -5.223287595432216e-19

R98_127 V98 V127 366.338771859072
L98_127 V98 V127 7.224583497313277e-12
C98_127 V98 V127 2.662895972908793e-20

R98_128 V98 V128 376.53212986675294
L98_128 V98 V128 2.0975206776553145e-12
C98_128 V98 V128 6.676590843765415e-20

R98_129 V98 V129 173.12955953164305
L98_129 V98 V129 6.085555541184791e-12
C98_129 V98 V129 -2.6542889831638678e-19

R98_130 V98 V130 -157.32526095355743
L98_130 V98 V130 2.603151143460632e-12
C98_130 V98 V130 2.5838064595989725e-19

R98_131 V98 V131 -174.52231288220372
L98_131 V98 V131 2.1516377229227376e-12
C98_131 V98 V131 3.323779023973822e-19

R98_132 V98 V132 -129.8295324990585
L98_132 V98 V132 1.5126706530692125e-12
C98_132 V98 V132 5.552805095594703e-19

R98_133 V98 V133 -311.8854011770016
L98_133 V98 V133 -3.406872959440303e-12
C98_133 V98 V133 1.8212150261617342e-19

R98_134 V98 V134 -379.77088607284855
L98_134 V98 V134 1.4418931744029093e-12
C98_134 V98 V134 2.2493048418853803e-19

R98_135 V98 V135 940.5074408598153
L98_135 V98 V135 -1.6638645316510725e-12
C98_135 V98 V135 -4.546126731423875e-19

R98_136 V98 V136 1337.6946882990471
L98_136 V98 V136 -1.1038761230124723e-12
C98_136 V98 V136 -6.468492093857e-19

R98_137 V98 V137 -981.3056907070797
L98_137 V98 V137 7.975402803750689e-12
C98_137 V98 V137 1.0041426271073769e-19

R98_138 V98 V138 196.33082870355287
L98_138 V98 V138 -8.572235382248062e-13
C98_138 V98 V138 -3.871080617097022e-19

R98_139 V98 V139 352.53037578515796
L98_139 V98 V139 1.2040241911571488e-12
C98_139 V98 V139 6.061245408757607e-19

R98_140 V98 V140 247.1813963433248
L98_140 V98 V140 1.2229261463953241e-12
C98_140 V98 V140 7.224236304661525e-19

R98_141 V98 V141 -829.8334436188952
L98_141 V98 V141 -3.722031543137184e-12
C98_141 V98 V141 -3.9005926987863793e-19

R98_142 V98 V142 1197.5923560120361
L98_142 V98 V142 -2.3385754969534915e-12
C98_142 V98 V142 -2.6433044867614462e-20

R98_143 V98 V143 -264.96414531047134
L98_143 V98 V143 -1.5994518928089672e-12
C98_143 V98 V143 -1.8787612590789328e-19

R98_144 V98 V144 -281.51631230072036
L98_144 V98 V144 -3.4609157835267996e-12
C98_144 V98 V144 -1.6424769977115093e-19

R98_145 V98 V145 287.41705727202907
L98_145 V98 V145 -2.298907387785274e-12
C98_145 V98 V145 -1.4774799853616985e-19

R98_146 V98 V146 -214.16800571388768
L98_146 V98 V146 8.629373043396479e-13
C98_146 V98 V146 2.4013499923782067e-19

R98_147 V98 V147 393.7707482171281
L98_147 V98 V147 -2.1643202295771756e-12
C98_147 V98 V147 -6.132994218000522e-19

R98_148 V98 V148 755.1253681851856
L98_148 V98 V148 -1.0495123430853042e-12
C98_148 V98 V148 -4.8181362476076185e-19

R98_149 V98 V149 1824.0827968406613
L98_149 V98 V149 8.185537553709718e-13
C98_149 V98 V149 5.882567719225037e-19

R98_150 V98 V150 -414.3543901232306
L98_150 V98 V150 -6.943338915585124e-12
C98_150 V98 V150 -2.7380975689552966e-19

R98_151 V98 V151 334.3888520858102
L98_151 V98 V151 2.471121272710085e-12
C98_151 V98 V151 2.9628334612827586e-19

R98_152 V98 V152 171.74401529739285
L98_152 V98 V152 1.38633843430822e-12
C98_152 V98 V152 1.6378800794996415e-19

R98_153 V98 V153 -4713.080561903487
L98_153 V98 V153 3.997520195985864e-12
C98_153 V98 V153 4.5899579731046326e-20

R98_154 V98 V154 2175.5439501938704
L98_154 V98 V154 -4.391907976711556e-12
C98_154 V98 V154 4.3232790846672934e-21

R98_155 V98 V155 -367.8858545977367
L98_155 V98 V155 9.858354590781499e-13
C98_155 V98 V155 3.4907829112890737e-19

R98_156 V98 V156 -123.3619985075225
L98_156 V98 V156 -2.415495580743746e-11
C98_156 V98 V156 3.631382319310267e-19

R98_157 V98 V157 -240.92470428560662
L98_157 V98 V157 -7.636745451367553e-13
C98_157 V98 V157 -5.910476273819494e-19

R98_158 V98 V158 487.3107999580553
L98_158 V98 V158 -1.2038252018429029e-11
C98_158 V98 V158 1.9495703464376915e-19

R98_159 V98 V159 -196.67098965040304
L98_159 V98 V159 -1.2995175501760262e-12
C98_159 V98 V159 -2.3082733269110856e-19

R98_160 V98 V160 -202.95664150422772
L98_160 V98 V160 -3.3300116179865052e-12
C98_160 V98 V160 -1.859878394573414e-19

R98_161 V98 V161 138.161306013811
L98_161 V98 V161 1.8070064392450277e-12
C98_161 V98 V161 1.2016154109671591e-19

R98_162 V98 V162 190.5298715257787
L98_162 V98 V162 1.0462950548236317e-12
C98_162 V98 V162 1.4583497055685639e-19

R98_163 V98 V163 158.75028902421542
L98_163 V98 V163 6.591270011266422e-12
C98_163 V98 V163 8.30644537157828e-20

R98_164 V98 V164 106.06232888524414
L98_164 V98 V164 1.2464263921111472e-10
C98_164 V98 V164 1.7040912076169423e-19

R98_165 V98 V165 248.453858576783
L98_165 V98 V165 4.484827373118329e-12
C98_165 V98 V165 7.57619344806986e-20

R98_166 V98 V166 -160.54102642726838
L98_166 V98 V166 -2.117359449835137e-12
C98_166 V98 V166 -3.4671011877020358e-19

R98_167 V98 V167 1662.3957905195714
L98_167 V98 V167 4.757598428956883e-12
C98_167 V98 V167 6.413537000229743e-20

R98_168 V98 V168 1225.099828232304
L98_168 V98 V168 1.3595463446090353e-12
C98_168 V98 V168 -1.9320734432510222e-20

R98_169 V98 V169 -132.81192513376817
L98_169 V98 V169 -2.5904533976820154e-12
C98_169 V98 V169 -1.5474293735085636e-19

R98_170 V98 V170 -211.79204199844588
L98_170 V98 V170 -1.1818391247439956e-11
C98_170 V98 V170 2.6886284179266296e-19

R98_171 V98 V171 -231.44081895735786
L98_171 V98 V171 2.1931438714771858e-11
C98_171 V98 V171 -3.4700358954950576e-20

R98_172 V98 V172 -155.4960845273183
L98_172 V98 V172 -1.2820194573482789e-12
C98_172 V98 V172 -5.585835096301794e-20

R98_173 V98 V173 349.77082026299075
L98_173 V98 V173 4.376893263524116e-12
C98_173 V98 V173 7.369784947442148e-20

R98_174 V98 V174 134.59304038161474
L98_174 V98 V174 4.425295414312012e-12
C98_174 V98 V174 -9.343250932143376e-20

R98_175 V98 V175 33109.347319236134
L98_175 V98 V175 3.44438553798839e-12
C98_175 V98 V175 2.6906311378284746e-19

R98_176 V98 V176 706.52781774614
L98_176 V98 V176 1.9211858059151017e-12
C98_176 V98 V176 3.3074564404336444e-19

R98_177 V98 V177 280.2946576327361
L98_177 V98 V177 -2.791766719145245e-12
C98_177 V98 V177 -1.3801724225227322e-19

R98_178 V98 V178 215.99352970238357
L98_178 V98 V178 -1.6837472219754105e-11
C98_178 V98 V178 -1.214327119915128e-19

R98_179 V98 V179 574.4736858863017
L98_179 V98 V179 -2.444495945583729e-12
C98_179 V98 V179 -3.4835763412193207e-19

R98_180 V98 V180 487.82293093984345
L98_180 V98 V180 -3.822555973092941e-12
C98_180 V98 V180 -3.7897171378717744e-19

R98_181 V98 V181 -217.65618691758587
L98_181 V98 V181 2.936257656232937e-12
C98_181 V98 V181 9.649121608011697e-20

R98_182 V98 V182 -111.1185867206112
L98_182 V98 V182 8.126717942357944e-11
C98_182 V98 V182 9.997147931590456e-20

R98_183 V98 V183 -532.8186199966963
L98_183 V98 V183 -1.8118129087708608e-12
C98_183 V98 V183 -2.2097064885314937e-20

R98_184 V98 V184 -514.390078413301
L98_184 V98 V184 -1.6328648725521403e-12
C98_184 V98 V184 3.0892015017890886e-20

R98_185 V98 V185 4633.012475866189
L98_185 V98 V185 4.9385565863996345e-12
C98_185 V98 V185 7.834646889552644e-20

R98_186 V98 V186 -255.93701864926072
L98_186 V98 V186 -1.5099679779963165e-12
C98_186 V98 V186 -7.141541844042085e-20

R98_187 V98 V187 686.8900248564132
L98_187 V98 V187 1.420163168663226e-12
C98_187 V98 V187 3.4264032034742706e-19

R98_188 V98 V188 243.02106659650107
L98_188 V98 V188 6.279728122495335e-13
C98_188 V98 V188 2.9277026090525945e-19

R98_189 V98 V189 1358.1587447326838
L98_189 V98 V189 -1.964210237594364e-12
C98_189 V98 V189 -1.858445324419484e-19

R98_190 V98 V190 130.99551958590345
L98_190 V98 V190 2.6576196648659897e-12
C98_190 V98 V190 -7.902636682572583e-20

R98_191 V98 V191 254.60810065749845
L98_191 V98 V191 1.5525077520676544e-12
C98_191 V98 V191 -1.8805100621753713e-19

R98_192 V98 V192 875.6331857228816
L98_192 V98 V192 -1.6988012769654945e-12
C98_192 V98 V192 -3.574590972498583e-19

R98_193 V98 V193 983.145334467408
L98_193 V98 V193 1.1241719001515219e-11
C98_193 V98 V193 -6.615444859735215e-21

R98_194 V98 V194 -377.2899009638497
L98_194 V98 V194 -1.4023518110925595e-12
C98_194 V98 V194 -2.670328073231025e-19

R98_195 V98 V195 -277.9644957784848
L98_195 V98 V195 -1.279988691476627e-12
C98_195 V98 V195 3.1717308994857675e-20

R98_196 V98 V196 -461.87480995863666
L98_196 V98 V196 5.13356341899063e-12
C98_196 V98 V196 4.011051006611277e-19

R98_197 V98 V197 -1303.408444089135
L98_197 V98 V197 4.672961136815561e-12
C98_197 V98 V197 7.56806557704912e-20

R98_198 V98 V198 -172.47000537884566
L98_198 V98 V198 -1.0770250864437234e-11
C98_198 V98 V198 -7.203035435003801e-21

R98_199 V98 V199 -365.37593233489235
L98_199 V98 V199 9.2831297330179e-12
C98_199 V98 V199 1.1605452219641954e-19

R98_200 V98 V200 -1361.9212793236568
L98_200 V98 V200 7.440858411774915e-12
C98_200 V98 V200 6.163861241100395e-20

R99_99 V99 0 425.2206887184873
L99_99 V99 0 -2.6529144188081764e-13
C99_99 V99 0 -2.1241208551017326e-18

R99_100 V99 V100 -215.20901706496724
L99_100 V99 V100 -1.691066736005669e-12
C99_100 V99 V100 -2.767718298164533e-19

R99_101 V99 V101 1117.653143488928
L99_101 V99 V101 -1.7523944430978538e-12
C99_101 V99 V101 -4.911839931014865e-19

R99_102 V99 V102 -420.38533955174165
L99_102 V99 V102 -1.2053014593526403e-12
C99_102 V99 V102 -4.56536474482293e-19

R99_103 V99 V103 124.90879215832317
L99_103 V99 V103 4.0205713065878216e-13
C99_103 V99 V103 9.731640924965186e-19

R99_104 V99 V104 -1242.0809580406717
L99_104 V99 V104 1.5499018093521762e-12
C99_104 V99 V104 1.3238301756985772e-19

R99_105 V99 V105 -658.756566186774
L99_105 V99 V105 -1.1602360011736061e-12
C99_105 V99 V105 -4.2991675939285223e-19

R99_106 V99 V106 -1402.0939503468305
L99_106 V99 V106 -5.89043265983171e-13
C99_106 V99 V106 -8.87254818530564e-19

R99_107 V99 V107 63.490611163339246
L99_107 V99 V107 5.468833435107461e-13
C99_107 V99 V107 8.997650573954733e-19

R99_108 V99 V108 436.1490213966654
L99_108 V99 V108 -3.2988639765667393e-12
C99_108 V99 V108 -6.420390777025101e-20

R99_109 V99 V109 -263.55500330642707
L99_109 V99 V109 1.2017382661574468e-12
C99_109 V99 V109 6.57028820284649e-19

R99_110 V99 V110 718.657889232729
L99_110 V99 V110 9.733118059220888e-13
C99_110 V99 V110 5.718428967186309e-19

R99_111 V99 V111 -62.73470140685968
L99_111 V99 V111 -1.433782411644532e-12
C99_111 V99 V111 1.21898575192071e-21

R99_112 V99 V112 -423.3563115849314
L99_112 V99 V112 -9.793653467093107e-12
C99_112 V99 V112 -2.178374313491407e-19

R99_113 V99 V113 93.21057212580521
L99_113 V99 V113 1.78088546194976e-12
C99_113 V99 V113 1.1717243830622135e-19

R99_114 V99 V114 595.0182249866449
L99_114 V99 V114 6.569565270488626e-13
C99_114 V99 V114 8.584821377006256e-19

R99_115 V99 V115 -194.10539065819063
L99_115 V99 V115 -4.2772629940702204e-13
C99_115 V99 V115 -9.017009280998337e-19

R99_116 V99 V116 -881.5375847669316
L99_116 V99 V116 -1.2293355270555675e-10
C99_116 V99 V116 2.9148358464265797e-19

R99_117 V99 V117 440.24640755126717
L99_117 V99 V117 -1.430313660792806e-12
C99_117 V99 V117 -3.1560450066735394e-19

R99_118 V99 V118 -494.22080408314787
L99_118 V99 V118 -6.169106444473248e-13
C99_118 V99 V118 -9.745101719394277e-19

R99_119 V99 V119 75.03948843744088
L99_119 V99 V119 1.0777252328508794e-12
C99_119 V99 V119 -1.9706306561215129e-19

R99_120 V99 V120 336.0443653979237
L99_120 V99 V120 -2.5263537144951085e-12
C99_120 V99 V120 -3.607956273451777e-19

R99_121 V99 V121 -112.246130985686
L99_121 V99 V121 -6.782278674919853e-12
C99_121 V99 V121 1.156205934002968e-19

R99_122 V99 V122 -698.0586247315949
L99_122 V99 V122 -8.541094713985164e-12
C99_122 V99 V122 2.3577450949471166e-20

R99_123 V99 V123 -110.02428638867656
L99_123 V99 V123 4.667766248037767e-13
C99_123 V99 V123 1.6447878218716069e-18

R99_124 V99 V124 -371.03077256899917
L99_124 V99 V124 1.7393345381814817e-12
C99_124 V99 V124 7.502260166321983e-20

R99_125 V99 V125 1762.6895583436958
L99_125 V99 V125 3.636704948410436e-12
C99_125 V99 V125 -1.0352322658366215e-19

R99_126 V99 V126 430.9420415045505
L99_126 V99 V126 5.676181790163105e-13
C99_126 V99 V126 7.502918456496712e-19

R99_127 V99 V127 -3251.1028247289264
L99_127 V99 V127 -5.124778264297113e-13
C99_127 V99 V127 -9.210505242083182e-19

R99_128 V99 V128 -560.6303128722373
L99_128 V99 V128 4.047713706078124e-12
C99_128 V99 V128 4.583468510962602e-19

R99_129 V99 V129 127.23832329631058
L99_129 V99 V129 1.7227713141757577e-12
C99_129 V99 V129 5.438873378803607e-19

R99_130 V99 V130 1659.44517422365
L99_130 V99 V130 -1.0375233132582238e-12
C99_130 V99 V130 -4.585434424096874e-19

R99_131 V99 V131 500.35983700613576
L99_131 V99 V131 4.425436762467493e-12
C99_131 V99 V131 -2.609727286462255e-19

R99_132 V99 V132 282.6515720888261
L99_132 V99 V132 -9.16003330198569e-13
C99_132 V99 V132 -9.0362127161384e-19

R99_133 V99 V133 934.2654635205558
L99_133 V99 V133 -2.4249163855771153e-12
C99_133 V99 V133 -3.8908341802208903e-19

R99_134 V99 V134 352.79137995326226
L99_134 V99 V134 -3.0110388148386215e-11
C99_134 V99 V134 -8.762319142869329e-23

R99_135 V99 V135 -81.52786512960677
L99_135 V99 V135 5.750345018990433e-13
C99_135 V99 V135 1.826750958454248e-18

R99_136 V99 V136 -2775.6712340875324
L99_136 V99 V136 7.1087376049104245e-12
C99_136 V99 V136 -2.2687910404420776e-20

R99_137 V99 V137 -189.62431833437893
L99_137 V99 V137 -1.6749764287469851e-12
C99_137 V99 V137 -2.9687622021699446e-19

R99_138 V99 V138 -632.5846678877813
L99_138 V99 V138 1.1014356069533946e-12
C99_138 V99 V138 4.33243919915517e-19

R99_139 V99 V139 54.40018406209235
L99_139 V99 V139 -3.509526323747271e-13
C99_139 V99 V139 -2.5271081947807235e-18

R99_140 V99 V140 323.25145224103466
L99_140 V99 V140 4.093282041022267e-12
C99_140 V99 V140 2.558613157145162e-19

R99_141 V99 V141 -157.54229905461972
L99_141 V99 V141 8.835704128290459e-13
C99_141 V99 V141 8.299318569621247e-19

R99_142 V99 V142 -202.36655617828634
L99_142 V99 V142 -3.074168379059939e-12
C99_142 V99 V142 -8.708011298173297e-20

R99_143 V99 V143 883.7035107197669
L99_143 V99 V143 6.84926155002502e-13
C99_143 V99 V143 5.911957735990132e-19

R99_144 V99 V144 -348.05290002125275
L99_144 V99 V144 -1.2969568766741536e-10
C99_144 V99 V144 -6.259605520043318e-20

R99_145 V99 V145 99.81465280272873
L99_145 V99 V145 1.3914899313336655e-12
C99_145 V99 V145 2.6977028985877244e-19

R99_146 V99 V146 227.3239701592669
L99_146 V99 V146 -3.435955391217576e-12
C99_146 V99 V146 -2.8713897576249547e-19

R99_147 V99 V147 -73.57196546026536
L99_147 V99 V147 1.7225400258121303e-12
C99_147 V99 V147 1.5793397017814033e-18

R99_148 V99 V148 251.32424663469772
L99_148 V99 V148 2.2031543679638996e-12
C99_148 V99 V148 7.235118725090853e-20

R99_149 V99 V149 876.1146613041452
L99_149 V99 V149 -4.199522000707521e-13
C99_149 V99 V149 -1.3068671023096063e-18

R99_150 V99 V150 685.1846005829664
L99_150 V99 V150 3.152397374884902e-12
C99_150 V99 V150 3.930275559410732e-19

R99_151 V99 V151 -82.52430680025402
L99_151 V99 V151 -1.3032853381019669e-12
C99_151 V99 V151 -7.69178982919269e-19

R99_152 V99 V152 -399.59510210226364
L99_152 V99 V152 2.0434059196324667e-11
C99_152 V99 V152 8.437445205713729e-20

R99_153 V99 V153 -16477.331281742674
L99_153 V99 V153 1.6776842730778385e-11
C99_153 V99 V153 1.6598195526423227e-19

R99_154 V99 V154 -206.5975020901366
L99_154 V99 V154 2.7286470834183635e-11
C99_154 V99 V154 -6.240647307412432e-20

R99_155 V99 V155 44.53638652421951
L99_155 V99 V155 -5.404321916453869e-13
C99_155 V99 V155 -1.0509458056044663e-18

R99_156 V99 V156 -5991.9304948867375
L99_156 V99 V156 -3.3811452527751547e-12
C99_156 V99 V156 -2.445739098085097e-20

R99_157 V99 V157 -126.50362964310199
L99_157 V99 V157 5.693187279457361e-13
C99_157 V99 V157 8.862431145127232e-19

R99_158 V99 V158 -362.11870697148834
L99_158 V99 V158 -2.4121484553296886e-12
C99_158 V99 V158 -2.287400082357662e-19

R99_159 V99 V159 270.6179650483242
L99_159 V99 V159 4.662078545621993e-13
C99_159 V99 V159 9.390816865882856e-19

R99_160 V99 V160 -421.92122085166494
L99_160 V99 V160 -3.2837107489783318e-12
C99_160 V99 V160 -1.8716425223713483e-19

R99_161 V99 V161 218.5267602811881
L99_161 V99 V161 -1.5077051782858085e-12
C99_161 V99 V161 -2.337046689069837e-19

R99_162 V99 V162 382.094472209549
L99_162 V99 V162 -1.125499175418521e-12
C99_162 V99 V162 -3.3665569709506953e-19

R99_163 V99 V163 -434.2253316318767
L99_163 V99 V163 -1.3901114501747258e-12
C99_163 V99 V163 -4.295755441160657e-19

R99_164 V99 V164 283.72660557772105
L99_164 V99 V164 3.000650793058099e-12
C99_164 V99 V164 -1.0017823875708687e-19

R99_165 V99 V165 126.92039762380206
L99_165 V99 V165 3.823053708909922e-12
C99_165 V99 V165 -9.564009518547719e-20

R99_166 V99 V166 438.2918125285354
L99_166 V99 V166 1.8873535774835715e-12
C99_166 V99 V166 2.8288591450228486e-19

R99_167 V99 V167 -125.75806879718944
L99_167 V99 V167 -1.9433119558447505e-11
C99_167 V99 V167 -6.176919434582708e-20

R99_168 V99 V168 1228.410451175575
L99_168 V99 V168 -2.5836067920377354e-12
C99_168 V99 V168 3.616771430523195e-20

R99_169 V99 V169 -281.99994690411745
L99_169 V99 V169 2.17194734898669e-12
C99_169 V99 V169 4.0201146802413125e-19

R99_170 V99 V170 -735.5200860153857
L99_170 V99 V170 -1.203637269126588e-11
C99_170 V99 V170 -2.368243067974323e-19

R99_171 V99 V171 2274.75613391352
L99_171 V99 V171 -2.3236593396028893e-11
C99_171 V99 V171 1.8665997968126926e-19

R99_172 V99 V172 -791.6562428696616
L99_172 V99 V172 4.981116077992517e-12
C99_172 V99 V172 3.425786072794864e-20

R99_173 V99 V173 -326.62805703780816
L99_173 V99 V173 -1.108591421084374e-12
C99_173 V99 V173 -3.1118739433409614e-19

R99_174 V99 V174 -303.95715782425845
L99_174 V99 V174 -4.763877008995631e-12
C99_174 V99 V174 2.440501424618144e-19

R99_175 V99 V175 210.66277846367083
L99_175 V99 V175 -6.996268306317832e-13
C99_175 V99 V175 -9.517656345364887e-19

R99_176 V99 V176 1315.860728735254
L99_176 V99 V176 -4.199624372169136e-12
C99_176 V99 V176 -4.3476196721403114e-20

R99_177 V99 V177 384.6735119882217
L99_177 V99 V177 1.2126085639420906e-12
C99_177 V99 V177 7.109625387334519e-20

R99_178 V99 V178 3021.5151828292896
L99_178 V99 V178 2.4132784675650877e-12
C99_178 V99 V178 1.105507783998446e-19

R99_179 V99 V179 99.73466872405123
L99_179 V99 V179 7.327559224356076e-13
C99_179 V99 V179 8.89370697920657e-19

R99_180 V99 V180 -16785.30785904923
L99_180 V99 V180 1.760047132267653e-12
C99_180 V99 V180 2.4197011189370785e-19

R99_181 V99 V181 -1199.7494001568557
L99_181 V99 V181 -2.1339301535686624e-12
C99_181 V99 V181 1.1767981142046939e-19

R99_182 V99 V182 378.6578315685429
L99_182 V99 V182 -1.2395914086872897e-12
C99_182 V99 V182 -3.1401527419676347e-19

R99_183 V99 V183 -76.37352314840814
L99_183 V99 V183 1.1087273103251723e-12
C99_183 V99 V183 1.3349932598832517e-20

R99_184 V99 V184 -4738.780764456767
L99_184 V99 V184 1.4077312290622737e-12
C99_184 V99 V184 1.2896883657104463e-19

R99_185 V99 V185 -2143.9001420847744
L99_185 V99 V185 -3.2041190283219e-12
C99_185 V99 V185 -1.5199596848032104e-19

R99_186 V99 V186 -4509.586767562697
L99_186 V99 V186 1.5306788632582997e-12
C99_186 V99 V186 3.1045629238436605e-19

R99_187 V99 V187 -639.4087320385597
L99_187 V99 V187 -4.4331251105902244e-13
C99_187 V99 V187 -9.252027634994879e-19

R99_188 V99 V188 1360.8535526975563
L99_188 V99 V188 -7.219356606483079e-13
C99_188 V99 V188 -3.441128175504753e-19

R99_189 V99 V189 -1488.8057018095035
L99_189 V99 V189 1.9917330798518988e-12
C99_189 V99 V189 6.781558421786098e-20

R99_190 V99 V190 -822.0799493364447
L99_190 V99 V190 -1.4643232444792453e-10
C99_190 V99 V190 1.1312182870973649e-19

R99_191 V99 V191 97.67505549743947
L99_191 V99 V191 2.9166878655858514e-11
C99_191 V99 V191 6.390639661330903e-19

R99_192 V99 V192 761.4004243201375
L99_192 V99 V192 -3.0429139875983088e-12
C99_192 V99 V192 -5.061009390330067e-20

R99_193 V99 V193 1163.2168387825375
L99_193 V99 V193 -8.583101013089335e-12
C99_193 V99 V193 4.684081496470254e-20

R99_194 V99 V194 1311.1632301753098
L99_194 V99 V194 3.4530310017021475e-12
C99_194 V99 V194 3.1792167841950505e-19

R99_195 V99 V195 -158.39174475115746
L99_195 V99 V195 3.4720377567439087e-12
C99_195 V99 V195 -8.459564184573223e-19

R99_196 V99 V196 -414.8323244267398
L99_196 V99 V196 6.067143231533217e-13
C99_196 V99 V196 6.953201262040391e-19

R99_197 V99 V197 -897.4737851920888
L99_197 V99 V197 -4.3149814727609926e-11
C99_197 V99 V197 2.747809558125123e-20

R99_198 V99 V198 -760.0227012661549
L99_198 V99 V198 -7.456489990690527e-12
C99_198 V99 V198 -1.2806089443903236e-19

R99_199 V99 V199 -174.4879478614603
L99_199 V99 V199 -3.4890932202326123e-12
C99_199 V99 V199 -2.8512043588196955e-20

R99_200 V99 V200 -345.3402720334895
L99_200 V99 V200 -1.869533813261972e-12
C99_200 V99 V200 -3.260218108664526e-19

R100_100 V100 0 56.649576675380736
L100_100 V100 0 -1.9344789666073068e-13
C100_100 V100 0 -3.3843507274280194e-18

R100_101 V100 V101 1588.4629728292512
L100_101 V100 V101 -6.346508288172116e-12
C100_101 V100 V101 -3.323097117855855e-19

R100_102 V100 V102 -428.2766130792125
L100_102 V100 V102 -2.775680450483285e-12
C100_102 V100 V102 -2.838543001144166e-19

R100_103 V100 V103 -811.4071836206177
L100_103 V100 V103 8.466342054802225e-12
C100_103 V100 V103 9.320729704312284e-20

R100_104 V100 V104 137.16146372397316
L100_104 V100 V104 4.794658841788189e-13
C100_104 V100 V104 1.029047625872998e-18

R100_105 V100 V105 -334.7282397170636
L100_105 V100 V105 -1.8832324690596744e-12
C100_105 V100 V105 -3.413772635905025e-19

R100_106 V100 V106 -346.4320682502027
L100_106 V100 V106 -9.720369354766526e-13
C100_106 V100 V106 -6.496424593189917e-19

R100_107 V100 V107 425.2217366318826
L100_107 V100 V107 3.4709818907832056e-12
C100_107 V100 V107 2.2482088139871515e-19

R100_108 V100 V108 45.02789896856367
L100_108 V100 V108 2.1428581072557704e-12
C100_108 V100 V108 3.8668508845689505e-20

R100_109 V100 V109 -743.5862124366442
L100_109 V100 V109 2.1970935498899974e-12
C100_109 V100 V109 5.449954558397027e-19

R100_110 V100 V110 242.71012956025064
L100_110 V100 V110 2.310281179280252e-12
C100_110 V100 V110 1.923907623836717e-19

R100_111 V100 V111 -621.0494671738207
L100_111 V100 V111 -5.946815440467016e-12
C100_111 V100 V111 -2.110741949246407e-19

R100_112 V100 V112 -55.13142727205617
L100_112 V100 V112 1.847157040387054e-11
C100_112 V100 V112 5.549061774437841e-19

R100_113 V100 V113 96.65963853274762
L100_113 V100 V113 2.821482500738441e-12
C100_113 V100 V113 4.966255414782766e-20

R100_114 V100 V114 640.4889460036516
L100_114 V100 V114 1.0584935782801743e-12
C100_114 V100 V114 6.721736350280983e-19

R100_115 V100 V115 682.7809441488716
L100_115 V100 V115 1.0381062210871228e-11
C100_115 V100 V115 5.110262276059758e-20

R100_116 V100 V116 -94.4602228835574
L100_116 V100 V116 -7.497714982456814e-13
C100_116 V100 V116 -4.503569907091976e-19

R100_117 V100 V117 1208.3546905395553
L100_117 V100 V117 -2.71668368470538e-12
C100_117 V100 V117 -2.188669861275885e-19

R100_118 V100 V118 -210.56408157731983
L100_118 V100 V118 -1.28730978207387e-12
C100_118 V100 V118 -5.956143024025519e-19

R100_119 V100 V119 4359.211655441932
L100_119 V100 V119 -2.4129836335720482e-12
C100_119 V100 V119 -4.0802954466547934e-19

R100_120 V100 V120 48.78224209909709
L100_120 V100 V120 1.0817388526914658e-11
C100_120 V100 V120 -1.0282400635127904e-18

R100_121 V100 V121 -167.89335996503695
L100_121 V100 V121 1.1625028920873538e-11
C100_121 V100 V121 1.4189899153230876e-19

R100_122 V100 V122 520.1859936404401
L100_122 V100 V122 -3.807930244380256e-12
C100_122 V100 V122 -2.2837094736148003e-19

R100_123 V100 V123 -1023.7932793635813
L100_123 V100 V123 8.945028954356536e-12
C100_123 V100 V123 1.3375451847604635e-19

R100_124 V100 V124 -92.61260160893143
L100_124 V100 V124 4.564881593430871e-13
C100_124 V100 V124 2.1520459107744976e-18

R100_125 V100 V125 615.6430375640884
L100_125 V100 V125 3.5535173493764303e-12
C100_125 V100 V125 -6.438200236361026e-20

R100_126 V100 V126 311.18776081150367
L100_126 V100 V126 8.907339078894683e-13
C100_126 V100 V126 5.044390675310144e-19

R100_127 V100 V127 309.99963445442967
L100_127 V100 V127 9.186127667598728e-13
C100_127 V100 V127 5.950427735016823e-19

R100_128 V100 V128 -228.3815792744312
L100_128 V100 V128 -6.94581325994544e-13
C100_128 V100 V128 -4.946669204341166e-19

R100_129 V100 V129 166.11582221588685
L100_129 V100 V129 2.1394826461366532e-10
C100_129 V100 V129 2.8827696185767804e-19

R100_130 V100 V130 -886.4296351734495
L100_130 V100 V130 -2.0987904060236015e-12
C100_130 V100 V130 -2.8534178832234746e-19

R100_131 V100 V131 -336.88309849076614
L100_131 V100 V131 -9.669167315975009e-13
C100_131 V100 V131 -6.662751685179101e-19

R100_132 V100 V132 179.2402920405122
L100_132 V100 V132 -1.458675680110178e-10
C100_132 V100 V132 -8.090568680139072e-19

R100_133 V100 V133 739.2611919407638
L100_133 V100 V133 -8.575684328990428e-12
C100_133 V100 V133 -3.8216287332419443e-19

R100_134 V100 V134 298.5725690280647
L100_134 V100 V134 -1.675479450406939e-12
C100_134 V100 V134 -5.729704507748148e-19

R100_135 V100 V135 577.9583009841547
L100_135 V100 V135 -2.5754377906539025e-12
C100_135 V100 V135 -3.0717329243502336e-19

R100_136 V100 V136 -88.61776991241251
L100_136 V100 V136 7.48224288467283e-13
C100_136 V100 V136 1.630654050715471e-18

R100_137 V100 V137 -191.42757647287084
L100_137 V100 V137 1.497180731341432e-11
C100_137 V100 V137 1.4325989972601484e-19

R100_138 V100 V138 -606.5296445537292
L100_138 V100 V138 1.0984710778021307e-12
C100_138 V100 V138 6.755921733451526e-19

R100_139 V100 V139 409.69093898053336
L100_139 V100 V139 1.0265484428160963e-12
C100_139 V100 V139 5.323171947541086e-19

R100_140 V100 V140 65.53461250399323
L100_140 V100 V140 -6.59008310514105e-13
C100_140 V100 V140 -1.8823715740556696e-18

R100_141 V100 V141 -209.5070881719205
L100_141 V100 V141 4.171157524945701e-12
C100_141 V100 V141 3.7270705130989276e-19

R100_142 V100 V142 -341.45823030834464
L100_142 V100 V142 4.017944646472114e-12
C100_142 V100 V142 6.828759997518204e-20

R100_143 V100 V143 -298.95344719887584
L100_143 V100 V143 -1.314440045981422e-11
C100_143 V100 V143 -3.0255325871871853e-20

R100_144 V100 V144 128.86443655120712
L100_144 V100 V144 1.496162520560144e-12
C100_144 V100 V144 3.3833251492112673e-19

R100_145 V100 V145 98.50871349548933
L100_145 V100 V145 4.469223661403395e-12
C100_145 V100 V145 -1.0079866631879398e-19

R100_146 V100 V146 223.43639940065694
L100_146 V100 V146 -1.3997863793947764e-12
C100_146 V100 V146 -3.2735022686847527e-19

R100_147 V100 V147 873.1732231251914
L100_147 V100 V147 1.2137998186892812e-11
C100_147 V100 V147 1.407412002318776e-19

R100_148 V100 V148 -38.485703695358566
L100_148 V100 V148 1.0982823013840407e-12
C100_148 V100 V148 1.1279988123686042e-18

R100_149 V100 V149 1445.4802469509175
L100_149 V100 V149 -2.5730483816662474e-12
C100_149 V100 V149 -2.9352487307435746e-19

R100_150 V100 V150 -878.8642630453306
L100_150 V100 V150 3.988309893439266e-12
C100_150 V100 V150 2.2642869287674734e-19

R100_151 V100 V151 1529.5985830209388
L100_151 V100 V151 -5.5135318315454225e-12
C100_151 V100 V151 -1.0776704358736448e-20

R100_152 V100 V152 -328.33097372373834
L100_152 V100 V152 -6.715743462379319e-13
C100_152 V100 V152 -3.8266131886091626e-19

R100_153 V100 V153 -1352.9151321292518
L100_153 V100 V153 -2.6519090008394453e-12
C100_153 V100 V153 1.2732100847601221e-21

R100_154 V100 V154 -380.3306722585709
L100_154 V100 V154 -3.740200246985475e-12
C100_154 V100 V154 1.3048640054522038e-19

R100_155 V100 V155 -397.5443629002211
L100_155 V100 V155 -3.89542767545271e-12
C100_155 V100 V155 -6.635217643249605e-20

R100_156 V100 V156 117.59630170086359
L100_156 V100 V156 1.4954013239870897e-12
C100_156 V100 V156 -8.97581808385497e-19

R100_157 V100 V157 -114.10578088654134
L100_157 V100 V157 1.4141160734715263e-12
C100_157 V100 V157 6.118117853008196e-19

R100_158 V100 V158 -193.9964453530939
L100_158 V100 V158 1.1905464600817836e-11
C100_158 V100 V158 -1.4200285176490449e-19

R100_159 V100 V159 -193.7484612583093
L100_159 V100 V159 -8.157210927739515e-12
C100_159 V100 V159 -8.925745220522423e-20

R100_160 V100 V160 62.49977568495193
L100_160 V100 V160 1.2666006249528659e-12
C100_160 V100 V160 6.008627636131529e-19

R100_161 V100 V161 250.54771071744594
L100_161 V100 V161 -1.3184248315367e-12
C100_161 V100 V161 -3.4030478810628085e-19

R100_162 V100 V162 303.4352453440745
L100_162 V100 V162 -2.5245741634487737e-12
C100_162 V100 V162 -1.4717884456046522e-19

R100_163 V100 V163 284.0325029409764
L100_163 V100 V163 -1.541446541360962e-11
C100_163 V100 V163 7.306640347230143e-20

R100_164 V100 V164 -75.35006054606238
L100_164 V100 V164 -1.647417768669827e-12
C100_164 V100 V164 -3.989225713669045e-19

R100_165 V100 V165 195.6068620915484
L100_165 V100 V165 1.0869673098776624e-12
C100_165 V100 V165 1.7490895890484472e-19

R100_166 V100 V166 1253.7239542424243
L100_166 V100 V166 2.7371407280376457e-12
C100_166 V100 V166 3.271289591718158e-19

R100_167 V100 V167 -230.0975300593789
L100_167 V100 V167 -5.807839703115081e-12
C100_167 V100 V167 -1.2111382639564882e-19

R100_168 V100 V168 453.52878466218766
L100_168 V100 V168 -2.4900984632003925e-12
C100_168 V100 V168 -7.395196414283856e-20

R100_169 V100 V169 -349.1190763688498
L100_169 V100 V169 3.99828372877299e-12
C100_169 V100 V169 4.696547804585364e-19

R100_170 V100 V170 -364.83848720379103
L100_170 V100 V170 -5.726135671577445e-12
C100_170 V100 V170 -1.1322493173743725e-19

R100_171 V100 V171 -4482.461387976446
L100_171 V100 V171 -1.5747928291376545e-11
C100_171 V100 V171 3.4380329475480587e-20

R100_172 V100 V172 -320.3620337109566
L100_172 V100 V172 1.0510939521402535e-12
C100_172 V100 V172 2.586156554237788e-19

R100_173 V100 V173 -300.18257316810184
L100_173 V100 V173 -1.0201069189118081e-12
C100_173 V100 V173 -3.8327685908497e-19

R100_174 V100 V174 2456.2326739089217
L100_174 V100 V174 4.691220611283323e-10
C100_174 V100 V174 1.0763346261166613e-19

R100_175 V100 V175 1473.7914675074926
L100_175 V100 V175 3.813021044476373e-12
C100_175 V100 V175 4.910920771206336e-20

R100_176 V100 V176 416.6028086854477
L100_176 V100 V176 -9.92634445383943e-13
C100_176 V100 V176 -8.423806977297763e-19

R100_177 V100 V177 1334.7355463642634
L100_177 V100 V177 2.1103629647501183e-12
C100_177 V100 V177 1.0785359375459206e-19

R100_178 V100 V178 -1446.5500590167494
L100_178 V100 V178 1.254335131510667e-11
C100_178 V100 V178 1.248821955376373e-20

R100_179 V100 V179 -391.1730977063587
L100_179 V100 V179 2.556421408260277e-11
C100_179 V100 V179 1.0398430474357265e-19

R100_180 V100 V180 64.6494925772111
L100_180 V100 V180 1.2027858597711584e-12
C100_180 V100 V180 6.557225226623274e-19

R100_181 V100 V181 2202.6704319837777
L100_181 V100 V181 -2.3093717100217188e-11
C100_181 V100 V181 2.6635690818258064e-20

R100_182 V100 V182 653.5953780890064
L100_182 V100 V182 1.0614204830764419e-11
C100_182 V100 V182 2.033890201942414e-20

R100_183 V100 V183 304.05557947068513
L100_183 V100 V183 2.4166939510346767e-12
C100_183 V100 V183 1.782052371647843e-19

R100_184 V100 V184 -73.80866576244858
L100_184 V100 V184 2.6154147496719174e-12
C100_184 V100 V184 -9.507081748094283e-20

R100_185 V100 V185 -829.9893607262167
L100_185 V100 V185 -4.8769634205075645e-12
C100_185 V100 V185 -7.7399018247646e-20

R100_186 V100 V186 2870.96491888056
L100_186 V100 V186 1.3630711403069536e-12
C100_186 V100 V186 1.425381081666556e-20

R100_187 V100 V187 336.97467634465164
L100_187 V100 V187 2.8930474496479876e-12
C100_187 V100 V187 -2.0854847273330084e-19

R100_188 V100 V188 -266.1971446281221
L100_188 V100 V188 -4.589411625894199e-13
C100_188 V100 V188 -4.924361156926087e-19

R100_189 V100 V189 -883.4543263958537
L100_189 V100 V189 2.517614332345672e-12
C100_189 V100 V189 1.7557927151662353e-19

R100_190 V100 V190 -567.2626624379416
L100_190 V100 V190 -3.0316584431738818e-12
C100_190 V100 V190 2.193011262010298e-20

R100_191 V100 V191 -314.6991447948191
L100_191 V100 V191 -9.37345444227993e-13
C100_191 V100 V191 -1.7806742256481777e-19

R100_192 V100 V192 74.66078588069134
L100_192 V100 V192 5.803442507675565e-13
C100_192 V100 V192 8.0477539273662045e-19

R100_193 V100 V193 246.00206039315484
L100_193 V100 V193 -1.722993525048347e-11
C100_193 V100 V193 8.542980428487902e-20

R100_194 V100 V194 -23969.61722408227
L100_194 V100 V194 1.923576686697172e-12
C100_194 V100 V194 6.026048979388426e-19

R100_195 V100 V195 13212.552960794495
L100_195 V100 V195 7.929895506382627e-13
C100_195 V100 V195 7.393834150217395e-19

R100_196 V100 V196 -99.12852571088307
L100_196 V100 V196 -5.882227054905125e-13
C100_196 V100 V196 -1.3839874411186818e-18

R100_197 V100 V197 -8995.670604926614
L100_197 V100 V197 -3.889736389838946e-12
C100_197 V100 V197 -2.2782463845237936e-19

R100_198 V100 V198 -393.0255681477241
L100_198 V100 V198 5.354849557259382e-12
C100_198 V100 V198 1.276094893391493e-19

R100_199 V100 V199 -151.73434354106894
L100_199 V100 V199 -4.827780365423208e-12
C100_199 V100 V199 -1.2815167775745675e-19

R100_200 V100 V200 -446.01912670163085
L100_200 V100 V200 -6.219590737803636e-12
C100_200 V100 V200 1.088051347373562e-19

R101_101 V101 0 -94.73657077751628
L101_101 V101 0 2.1607679827090458e-11
C101_101 V101 0 -6.965424858141082e-19

R101_102 V101 V102 488.8180127851332
L101_102 V101 V102 -1.8596227373754843e-12
C101_102 V101 V102 -3.60117012005285e-19

R101_103 V101 V103 549.8820064834672
L101_103 V101 V103 3.6417298305602704e-11
C101_103 V101 V103 -1.0023749157319901e-20

R101_104 V101 V104 443.8413316284373
L101_104 V101 V104 4.948138267186616e-12
C101_104 V101 V104 -1.5684850960260535e-20

R101_105 V101 V105 84.49549154563454
L101_105 V101 V105 -4.620362015392505e-12
C101_105 V101 V105 -1.8654318531430225e-19

R101_106 V101 V106 -4554.718657661511
L101_106 V101 V106 -3.2703600771548886e-12
C101_106 V101 V106 -3.4833375019059002e-19

R101_107 V101 V107 -261.9988080216042
L101_107 V101 V107 2.2344987975825456e-12
C101_107 V101 V107 2.8993864143155344e-19

R101_108 V101 V108 -266.0834221694199
L101_108 V101 V108 -2.856683570867011e-12
C101_108 V101 V108 -1.1823153189180974e-19

R101_109 V101 V109 395.7253179466926
L101_109 V101 V109 1.436643932392458e-12
C101_109 V101 V109 5.844984219483271e-19

R101_110 V101 V110 -323.0698206744969
L101_110 V101 V110 3.178797976528357e-12
C101_110 V101 V110 3.179353455564849e-19

R101_111 V101 V111 -1445.819994645801
L101_111 V101 V111 -7.615288872154036e-12
C101_111 V101 V111 -9.493986042150687e-20

R101_112 V101 V112 -1477.5425119833035
L101_112 V101 V112 4.78520676931839e-12
C101_112 V101 V112 1.5453260939670648e-19

R101_113 V101 V113 -81.60384684572206
L101_113 V101 V113 1.828667434639479e-11
C101_113 V101 V113 1.463779925029336e-19

R101_114 V101 V114 1220.4815096637176
L101_114 V101 V114 2.2404639510980324e-12
C101_114 V101 V114 3.699484077317445e-19

R101_115 V101 V115 220.7922747266628
L101_115 V101 V115 -2.817318515114752e-12
C101_115 V101 V115 -6.791118186213959e-20

R101_116 V101 V116 212.66880441643806
L101_116 V101 V116 -2.4173618123610523e-10
C101_116 V101 V116 1.6776661734989934e-19

R101_117 V101 V117 433.6298169734325
L101_117 V101 V117 -7.89242205108329e-12
C101_117 V101 V117 7.564153697465515e-20

R101_118 V101 V118 230.23494614931786
L101_118 V101 V118 -1.609072257205236e-12
C101_118 V101 V118 -5.136168962022277e-19

R101_119 V101 V119 -548.7697500845024
L101_119 V101 V119 -1.2314881233419243e-11
C101_119 V101 V119 -1.6042933681718467e-19

R101_120 V101 V120 -291.5436601365692
L101_120 V101 V120 -2.926941188649022e-12
C101_120 V101 V120 -3.6775239630545217e-19

R101_121 V101 V121 110.09252458677878
L101_121 V101 V121 -3.661883659165842e-12
C101_121 V101 V121 -4.984030269381655e-19

R101_122 V101 V122 -372.13986318628207
L101_122 V101 V122 5.518172881390617e-12
C101_122 V101 V122 1.2285355281346638e-19

R101_123 V101 V123 -729.7477398705977
L101_123 V101 V123 1.909171519379526e-12
C101_123 V101 V123 3.374909197866146e-19

R101_124 V101 V124 -3962.0108068566606
L101_124 V101 V124 1.5763686457029216e-12
C101_124 V101 V124 3.3388516816183885e-19

R101_125 V101 V125 1124.433548677204
L101_125 V101 V125 -1.6615459166639232e-12
C101_125 V101 V125 -2.3492265381270803e-19

R101_126 V101 V126 -182.34458888253954
L101_126 V101 V126 3.2253555507194764e-12
C101_126 V101 V126 1.0897935443796889e-19

R101_127 V101 V127 -823.0284947832588
L101_127 V101 V127 -7.544462063457053e-11
C101_127 V101 V127 -3.134458661672384e-20

R101_128 V101 V128 -12558.64819678306
L101_128 V101 V128 -3.430646726552834e-12
C101_128 V101 V128 -5.512104876052885e-20

R101_129 V101 V129 -116.10861647832307
L101_129 V101 V129 1.5023844771876517e-12
C101_129 V101 V129 6.759239436636337e-19

R101_130 V101 V130 258.35506889637895
L101_130 V101 V130 -2.5662312181928334e-12
C101_130 V101 V130 -1.4423257008541242e-19

R101_131 V101 V131 441.7883500207843
L101_131 V101 V131 -3.2692654014450555e-12
C101_131 V101 V131 -1.801117878373909e-19

R101_132 V101 V132 821.0489508814882
L101_132 V101 V132 -3.500978078564252e-12
C101_132 V101 V132 -1.8436212280490378e-19

R101_133 V101 V133 -1169.7165364768505
L101_133 V101 V133 -6.4128310427523885e-12
C101_133 V101 V133 -1.937663130672482e-19

R101_134 V101 V134 440.3391057774347
L101_134 V101 V134 2.2332975724687013e-12
C101_134 V101 V134 1.954440564266602e-19

R101_135 V101 V135 265.5378061970545
L101_135 V101 V135 8.090227459322893e-12
C101_135 V101 V135 1.952521948473165e-19

R101_136 V101 V136 210.36488225979656
L101_136 V101 V136 2.2604384589663676e-12
C101_136 V101 V136 3.5158618354490027e-19

R101_137 V101 V137 97.01514205316613
L101_137 V101 V137 -9.840199179583654e-12
C101_137 V101 V137 -7.349684274259703e-20

R101_138 V101 V138 -449.12960108115686
L101_138 V101 V138 -6.64951560827683e-11
C101_138 V101 V138 -3.19474168190758e-20

R101_139 V101 V139 -175.75406062508907
L101_139 V101 V139 -2.9894238899114797e-12
C101_139 V101 V139 -3.288399817003342e-19

R101_140 V101 V140 -144.0603912490386
L101_140 V101 V140 -3.4782952219904406e-12
C101_140 V101 V140 -2.954268019397268e-19

R101_141 V101 V141 509.2302270814168
L101_141 V101 V141 1.937650107389994e-12
C101_141 V101 V141 1.852953459646139e-19

R101_142 V101 V142 -237.03477076051823
L101_142 V101 V142 -3.631000989042906e-12
C101_142 V101 V142 -1.0201394371591635e-19

R101_143 V101 V143 -349.96832216004765
L101_143 V101 V143 1.8746745336771593e-12
C101_143 V101 V143 2.9719807974416286e-19

R101_144 V101 V144 -286.9633934921727
L101_144 V101 V144 3.814291904330915e-10
C101_144 V101 V144 2.792736828978388e-21

R101_145 V101 V145 -92.33468046802577
L101_145 V101 V145 -3.3761439388344718e-12
C101_145 V101 V145 -1.0581054550075198e-21

R101_146 V101 V146 -335.5888994161712
L101_146 V101 V146 8.132627979376045e-12
C101_146 V101 V146 3.1053655757023965e-20

R101_147 V101 V147 335.91981332231046
L101_147 V101 V147 -1.2547512200778344e-11
C101_147 V101 V147 9.830177798982868e-20

R101_148 V101 V148 251.66105823235856
L101_148 V101 V148 2.34840552857754e-12
C101_148 V101 V148 1.0758511435028389e-19

R101_149 V101 V149 -258.4787522995165
L101_149 V101 V149 -7.803595557101954e-13
C101_149 V101 V149 -7.1799365287371e-19

R101_150 V101 V150 78.41458192839758
L101_150 V101 V150 -3.797252665813942e-11
C101_150 V101 V150 2.8127408006202664e-19

R101_151 V101 V151 224.12589990418027
L101_151 V101 V151 -2.9854306040731348e-12
C101_151 V101 V151 -2.875521493194792e-19

R101_152 V101 V152 572.125687437184
L101_152 V101 V152 -4.858396967727596e-12
C101_152 V101 V152 1.7396637067191122e-20

R101_153 V101 V153 83.48686914820968
L101_153 V101 V153 2.1279944661428572e-12
C101_153 V101 V153 3.286877639424496e-19

R101_154 V101 V154 329.5341156819753
L101_154 V101 V154 4.742331034529665e-12
C101_154 V101 V154 -1.4469481094310736e-19

R101_155 V101 V155 -730.1059391958495
L101_155 V101 V155 -2.558431511291301e-12
C101_155 V101 V155 -2.2780680546046783e-19

R101_156 V101 V156 431.1842133860682
L101_156 V101 V156 1.328080533649611e-11
C101_156 V101 V156 -1.1386175301749982e-19

R101_157 V101 V157 93.36463146172514
L101_157 V101 V157 6.295579564073322e-13
C101_157 V101 V157 8.774049021055579e-19

R101_158 V101 V158 -127.17837840141271
L101_158 V101 V158 -5.398843280417502e-12
C101_158 V101 V158 -9.017540502593921e-20

R101_159 V101 V159 -456.5633044210528
L101_159 V101 V159 2.2266814867900266e-12
C101_159 V101 V159 2.7198444684535826e-19

R101_160 V101 V160 -225.06246659686943
L101_160 V101 V160 4.028689576315725e-11
C101_160 V101 V160 8.878482575983222e-20

R101_161 V101 V161 -120.56094149270302
L101_161 V101 V161 -1.526840426765922e-12
C101_161 V101 V161 -4.413485313947215e-19

R101_162 V101 V162 -145.1197848888191
L101_162 V101 V162 -2.3643023060238504e-12
C101_162 V101 V162 7.495720321795026e-20

R101_163 V101 V163 -168.2049351892314
L101_163 V101 V163 3.359206705154257e-12
C101_163 V101 V163 2.239486778025396e-19

R101_164 V101 V164 -148.4725364869678
L101_164 V101 V164 7.75081751877124e-12
C101_164 V101 V164 -4.950295976008454e-20

R101_165 V101 V165 -217.65196568469491
L101_165 V101 V165 -7.371862140798724e-13
C101_165 V101 V165 -5.231671523271996e-19

R101_166 V101 V166 99.8568068402134
L101_166 V101 V166 -2.8660018978954334e-11
C101_166 V101 V166 -7.05129994806359e-21

R101_167 V101 V167 393.74059987469326
L101_167 V101 V167 -3.5165047581564166e-12
C101_167 V101 V167 -2.4852928422321124e-19

R101_168 V101 V168 639.264889845611
L101_168 V101 V168 -2.2635919450446913e-12
C101_168 V101 V168 -2.1675269090882095e-19

R101_169 V101 V169 109.036207158439
L101_169 V101 V169 1.5132514353166578e-12
C101_169 V101 V169 4.057914275249265e-19

R101_170 V101 V170 774.3761087559708
L101_170 V101 V170 -4.4999813563411015e-12
C101_170 V101 V170 -3.558595860398457e-19

R101_171 V101 V171 200.20620082268556
L101_171 V101 V171 -1.4080526952504981e-12
C101_171 V101 V171 -3.74237968455937e-19

R101_172 V101 V172 225.57546586165137
L101_172 V101 V172 3.615721210612292e-11
C101_172 V101 V172 -6.911375019171955e-20

R101_173 V101 V173 10492.17295939096
L101_173 V101 V173 2.452433080475705e-12
C101_173 V101 V173 3.5848926832365476e-19

R101_174 V101 V174 -130.15616244564725
L101_174 V101 V174 1.3601739425440501e-12
C101_174 V101 V174 5.609284318550943e-19

R101_175 V101 V175 -364.28041751065126
L101_175 V101 V175 2.0524541979543817e-12
C101_175 V101 V175 1.8221580302597805e-19

R101_176 V101 V176 -343.99957063228055
L101_176 V101 V176 2.1487595444873242e-12
C101_176 V101 V176 2.211058328791854e-19

R101_177 V101 V177 -205.06292925750392
L101_177 V101 V177 4.710441062532448e-12
C101_177 V101 V177 -2.630575594073717e-19

R101_178 V101 V178 1824.0804365665376
L101_178 V101 V178 9.63368421042006e-12
C101_178 V101 V178 1.3332598152130648e-19

R101_179 V101 V179 -414.88725460023505
L101_179 V101 V179 2.3180093161623657e-12
C101_179 V101 V179 4.219565497709221e-19

R101_180 V101 V180 -304.70697796367733
L101_180 V101 V180 4.771188624552416e-12
C101_180 V101 V180 2.636480252186762e-19

R101_181 V101 V181 448.22186716479143
L101_181 V101 V181 -1.3580131718587935e-12
C101_181 V101 V181 -4.865117458399238e-19

R101_182 V101 V182 132.32175958643896
L101_182 V101 V182 -1.1678622468568503e-12
C101_182 V101 V182 -3.338900594952878e-19

R101_183 V101 V183 676.1093996368693
L101_183 V101 V183 2.0080787715255306e-12
C101_183 V101 V183 1.944649937585774e-20

R101_184 V101 V184 462.417392737099
L101_184 V101 V184 4.938747456321843e-12
C101_184 V101 V184 -1.192966763469807e-19

R101_185 V101 V185 203.3067736725849
L101_185 V101 V185 -4.210029318288255e-12
C101_185 V101 V185 4.100945892520093e-19

R101_186 V101 V186 -773.9587697106421
L101_186 V101 V186 -3.848957809198018e-11
C101_186 V101 V186 -2.0324485813444731e-19

R101_187 V101 V187 -1508.005231137248
L101_187 V101 V187 -1.2210227512326265e-12
C101_187 V101 V187 -4.347113042302896e-19

R101_188 V101 V188 741.4492235809641
L101_188 V101 V188 -8.058889612720544e-13
C101_188 V101 V188 -4.4534864434653e-19

R101_189 V101 V189 -219.1802245053477
L101_189 V101 V189 1.6703231294859516e-12
C101_189 V101 V189 5.222049360755879e-20

R101_190 V101 V190 -268.55609267675686
L101_190 V101 V190 6.0925340584041785e-12
C101_190 V101 V190 2.712365742674659e-19

R101_191 V101 V191 1027.169623584494
L101_191 V101 V191 -1.1979739410559425e-12
C101_191 V101 V191 -7.056741932129704e-20

R101_192 V101 V192 -561.6793275816945
L101_192 V101 V192 4.926046227762385e-12
C101_192 V101 V192 2.955790671352759e-19

R101_193 V101 V193 -319.4699111943904
L101_193 V101 V193 6.042029640099179e-11
C101_193 V101 V193 1.960665172772513e-19

R101_194 V101 V194 231.07523149269736
L101_194 V101 V194 1.4075746341998156e-12
C101_194 V101 V194 4.1836084183756613e-19

R101_195 V101 V195 1829.99200821371
L101_195 V101 V195 8.339239872686511e-13
C101_195 V101 V195 2.862511294655537e-19

R101_196 V101 V196 753.447921617212
L101_196 V101 V196 1.0676810998614723e-12
C101_196 V101 V196 1.7074350875793053e-19

R101_197 V101 V197 245.33865620619105
L101_197 V101 V197 6.743521068209613e-12
C101_197 V101 V197 -2.2726239268884004e-19

R101_198 V101 V198 278.7037923403493
L101_198 V101 V198 -1.9722130851132237e-11
C101_198 V101 V198 -9.314337555789606e-20

R101_199 V101 V199 -6393.7386108060155
L101_199 V101 V199 2.015568728367735e-12
C101_199 V101 V199 2.1262527995996832e-19

R101_200 V101 V200 -903.1403314129594
L101_200 V101 V200 8.354360682286286e-11
C101_200 V101 V200 -1.650801610436508e-19

R102_102 V102 0 -119.2521218963625
L102_102 V102 0 -2.8242144499862176e-13
C102_102 V102 0 -2.038787198794909e-18

R102_103 V102 V103 -2723.2401076610595
L102_103 V102 V103 2.947700491924763e-12
C102_103 V102 V103 1.4191379576172098e-19

R102_104 V102 V104 -1691.7398366221962
L102_104 V102 V104 1.9692526009473167e-12
C102_104 V102 V104 2.3811865186302674e-19

R102_105 V102 V105 -537.9688081116456
L102_105 V102 V105 -5.891233997857346e-12
C102_105 V102 V105 -1.7065733631770464e-19

R102_106 V102 V106 83.9043386929904
L102_106 V102 V106 2.079657320496314e-12
C102_106 V102 V106 4.0478165292029333e-19

R102_107 V102 V107 584.7716366361815
L102_107 V102 V107 2.544167045317934e-12
C102_107 V102 V107 2.455433961360357e-19

R102_108 V102 V108 441.33402812848885
L102_108 V102 V108 -3.06457317696063e-12
C102_108 V102 V108 -1.6120433200402148e-19

R102_109 V102 V109 -277.3744909989852
L102_109 V102 V109 2.4132576166127905e-12
C102_109 V102 V109 3.6793653363169743e-19

R102_110 V102 V110 -317.96356461922613
L102_110 V102 V110 9.84345931017217e-13
C102_110 V102 V110 6.9829541411052105e-19

R102_111 V102 V111 718.2323857356748
L102_111 V102 V111 -4.7282773305002545e-12
C102_111 V102 V111 -1.2975257532202476e-19

R102_112 V102 V112 1427.1666068794163
L102_112 V102 V112 -1.3059765011489912e-11
C102_112 V102 V112 -4.9093769340823564e-20

R102_113 V102 V113 281.4843739614908
L102_113 V102 V113 1.0201562038171422e-11
C102_113 V102 V113 1.1086666597010261e-19

R102_114 V102 V114 -108.84845751129124
L102_114 V102 V114 -2.178060548670081e-12
C102_114 V102 V114 -3.152629169135012e-19

R102_115 V102 V115 -300.5328131777873
L102_115 V102 V115 -2.2554421539458777e-12
C102_115 V102 V115 -1.7575046477727274e-19

R102_116 V102 V116 -280.6124386417527
L102_116 V102 V116 -5.1020158567187945e-11
C102_116 V102 V116 1.5056586366636295e-19

R102_117 V102 V117 244.54316941611583
L102_117 V102 V117 -4.173147513236548e-12
C102_117 V102 V117 -2.0959887587414854e-19

R102_118 V102 V118 79.54606903728354
L102_118 V102 V118 -1.1908977406453125e-12
C102_118 V102 V118 -7.461382071846205e-19

R102_119 V102 V119 599.4323560021332
L102_119 V102 V119 5.691520928572563e-12
C102_119 V102 V119 1.480345379384558e-20

R102_120 V102 V120 628.6565627657129
L102_120 V102 V120 -7.889484392152823e-12
C102_120 V102 V120 -2.2651837392676547e-19

R102_121 V102 V121 -154.59116732452566
L102_121 V102 V121 -8.726181903817613e-12
C102_121 V102 V121 -4.631709556028693e-20

R102_122 V102 V122 -580.7752949986982
L102_122 V102 V122 1.5225223555688323e-12
C102_122 V102 V122 6.237652683198127e-19

R102_123 V102 V123 368.56605212672935
L102_123 V102 V123 1.4760012132150933e-11
C102_123 V102 V123 1.9751246275348672e-20

R102_124 V102 V124 380.9385799124664
L102_124 V102 V124 3.5674925835086626e-12
C102_124 V102 V124 1.6948265065364123e-19

R102_125 V102 V125 -394.05925052120335
L102_125 V102 V125 9.219100657787506e-12
C102_125 V102 V125 5.006994893898793e-20

R102_126 V102 V126 -101.3518841538901
L102_126 V102 V126 1.6822052449433173e-12
C102_126 V102 V126 4.531758895488908e-19

R102_127 V102 V127 -229.91678308589914
L102_127 V102 V127 4.002716005514122e-11
C102_127 V102 V127 1.1804849312914719e-19

R102_128 V102 V128 -257.6705129767009
L102_128 V102 V128 -6.3169353679101e-12
C102_128 V102 V128 8.282652097376118e-20

R102_129 V102 V129 138.6044860350976
L102_129 V102 V129 1.902932484253044e-12
C102_129 V102 V129 4.419779684411411e-19

R102_130 V102 V130 133.93447074410676
L102_130 V102 V130 -1.1593117951483646e-12
C102_130 V102 V130 -7.281744084794289e-19

R102_131 V102 V131 317.89170850002847
L102_131 V102 V131 2.6727603417349946e-11
C102_131 V102 V131 -8.396504573328581e-20

R102_132 V102 V132 260.9076874228684
L102_132 V102 V132 -1.6656281558109383e-11
C102_132 V102 V132 -2.215565640525536e-19

R102_133 V102 V133 -2944.640341000884
L102_133 V102 V133 -1.8880017379764058e-12
C102_133 V102 V133 -4.448119947853586e-19

R102_134 V102 V134 606.7217835146338
L102_134 V102 V134 2.7912039585602477e-12
C102_134 V102 V134 4.1023788100158375e-19

R102_135 V102 V135 528.6749409073569
L102_135 V102 V135 -3.714906072752107e-12
C102_135 V102 V135 -8.370819197057373e-20

R102_136 V102 V136 294.95071245612763
L102_136 V102 V136 7.311866027342826e-12
C102_136 V102 V136 1.864369870235097e-19

R102_137 V102 V137 -168.5492725277459
L102_137 V102 V137 -1.56797455933448e-12
C102_137 V102 V137 -3.1472497902269413e-19

R102_138 V102 V138 -132.6933595238877
L102_138 V102 V138 3.5784662114200184e-12
C102_138 V102 V138 -1.913186177307406e-20

R102_139 V102 V139 -172.84013562665197
L102_139 V102 V139 -5.0048233840305444e-12
C102_139 V102 V139 -1.1109559505859045e-19

R102_140 V102 V140 -106.91205301550525
L102_140 V102 V140 -2.629302680132795e-12
C102_140 V102 V140 -2.4270337814708938e-19

R102_141 V102 V141 555.6651710572621
L102_141 V102 V141 9.082843412513176e-13
C102_141 V102 V141 7.797040684992192e-19

R102_142 V102 V142 2535.777745249597
L102_142 V102 V142 -5.311614123608095e-12
C102_142 V102 V142 -1.0350785020658677e-19

R102_143 V102 V143 248.73794244300788
L102_143 V102 V143 1.7875520897748876e-12
C102_143 V102 V143 2.8301973291924365e-19

R102_144 V102 V144 219.86396885996945
L102_144 V102 V144 3.4805803927274203e-12
C102_144 V102 V144 1.6225603331520141e-19

R102_145 V102 V145 134.7552400731244
L102_145 V102 V145 1.2447256047138985e-12
C102_145 V102 V145 2.943186853417793e-19

R102_146 V102 V146 55.31722138682436
L102_146 V102 V146 3.593951554518545e-12
C102_146 V102 V146 -3.5573563831730824e-20

R102_147 V102 V147 273.4472522511872
L102_147 V102 V147 4.666710918227895e-12
C102_147 V102 V147 1.3558183683822601e-19

R102_148 V102 V148 278.1089704399575
L102_148 V102 V148 1.790449881460547e-12
C102_148 V102 V148 1.644706658009045e-19

R102_149 V102 V149 -3069.5712452647635
L102_149 V102 V149 -4.281334235521322e-13
C102_149 V102 V149 -1.2231353945860698e-18

R102_150 V102 V150 -101.39413899269965
L102_150 V102 V150 -2.844205609384151e-12
C102_150 V102 V150 6.0034148501166895e-19

R102_151 V102 V151 -296.7634834499829
L102_151 V102 V151 -5.069165942514461e-12
C102_151 V102 V151 -2.08107903211753e-19

R102_152 V102 V152 -298.45362238366613
L102_152 V102 V152 -5.361798872283279e-12
C102_152 V102 V152 -1.6811125559685042e-20

R102_153 V102 V153 -114.92570238048525
L102_153 V102 V153 -2.924483408905192e-12
C102_153 V102 V153 -1.0480480608966852e-19

R102_154 V102 V154 -59.86260944689923
L102_154 V102 V154 -1.2010625984920115e-11
C102_154 V102 V154 -4.95706993096866e-19

R102_155 V102 V155 -361.46898957408484
L102_155 V102 V155 -1.3615916569356162e-12
C102_155 V102 V155 -2.5349560695483603e-19

R102_156 V102 V156 -352.0222210433242
L102_156 V102 V156 -2.388335179623333e-12
C102_156 V102 V156 -2.5669241891429305e-19

R102_157 V102 V157 -155.4059495286098
L102_157 V102 V157 4.979315739205123e-13
C102_157 V102 V157 1.1325440383365716e-18

R102_158 V102 V158 55.358290618514715
L102_158 V102 V158 3.877494791324237e-12
C102_158 V102 V158 4.096506541784559e-20

R102_159 V102 V159 341.87097192629267
L102_159 V102 V159 1.5535183774807226e-11
C102_159 V102 V159 -1.929661028912849e-20

R102_160 V102 V160 332.54840280958507
L102_160 V102 V160 -8.533098734375396e-12
C102_160 V102 V160 -5.809365660484907e-20

R102_161 V102 V161 201.48354444714755
L102_161 V102 V161 7.9465759079446e-12
C102_161 V102 V161 5.737921303482633e-20

R102_162 V102 V162 66.88057876335347
L102_162 V102 V162 -1.926763051313323e-12
C102_162 V102 V162 -1.0613937255283623e-19

R102_163 V102 V163 750.5494043257311
L102_163 V102 V163 1.5406014993496898e-12
C102_163 V102 V163 2.579767533778503e-19

R102_164 V102 V164 826.2248693531157
L102_164 V102 V164 1.6755418832585468e-12
C102_164 V102 V164 4.486242290045716e-20

R102_165 V102 V165 125.25877828150514
L102_165 V102 V165 -1.1844985669984045e-12
C102_165 V102 V165 -5.823627839056127e-19

R102_166 V102 V166 -38.93866591078675
L102_166 V102 V166 -3.571457895941122e-12
C102_166 V102 V166 1.6842377577484218e-19

R102_167 V102 V167 214.09351852844333
L102_167 V102 V167 -9.29976226382797e-11
C102_167 V102 V167 -1.0257706301084006e-20

R102_168 V102 V168 143.27880102304556
L102_168 V102 V168 -1.2651506022806869e-11
C102_168 V102 V168 1.6771495979788053e-19

R102_169 V102 V169 -237.62053357158447
L102_169 V102 V169 -3.650381999290707e-11
C102_169 V102 V169 1.1277711471647683e-19

R102_170 V102 V170 417.7450294927158
L102_170 V102 V170 1.7579296277507384e-12
C102_170 V102 V170 -3.513469358277288e-19

R102_171 V102 V171 -335.41910141321745
L102_171 V102 V171 -1.1151007821613408e-12
C102_171 V102 V171 -4.115719515921343e-19

R102_172 V102 V172 -241.776835709641
L102_172 V102 V172 -2.409482712519883e-12
C102_172 V102 V172 -2.643879306868501e-19

R102_173 V102 V173 -290.50518320961993
L102_173 V102 V173 2.9104299633251136e-12
C102_173 V102 V173 1.2956490901241593e-19

R102_174 V102 V174 43.21305652269133
L102_174 V102 V174 -6.33392116128551e-12
C102_174 V102 V174 1.9923244875231871e-19

R102_175 V102 V175 -380.3260701000531
L102_175 V102 V175 5.174659179829696e-11
C102_175 V102 V175 -6.823171473954553e-20

R102_176 V102 V176 -173.14250922139829
L102_176 V102 V176 -3.6220515033372045e-11
C102_176 V102 V176 -1.191587589133489e-19

R102_177 V102 V177 296.4386979302778
L102_177 V102 V177 4.343867231187897e-12
C102_177 V102 V177 -1.114942740055707e-19

R102_178 V102 V178 -122.95742854402786
L102_178 V102 V178 -2.7545891623935665e-12
C102_178 V102 V178 2.7540144752572773e-19

R102_179 V102 V179 446.78453956219664
L102_179 V102 V179 1.150004870487935e-12
C102_179 V102 V179 4.766221009403456e-19

R102_180 V102 V180 173.09829850925715
L102_180 V102 V180 1.1747585755310436e-12
C102_180 V102 V180 3.8200843782076776e-19

R102_181 V102 V181 3140.6968750747465
L102_181 V102 V181 3.8736672743285885e-11
C102_181 V102 V181 2.0347490138801847e-19

R102_182 V102 V182 -103.83374011112397
L102_182 V102 V182 -1.907209375011891e-12
C102_182 V102 V182 -2.9934617627284777e-19

R102_183 V102 V183 7897.276375012861
L102_183 V102 V183 3.1091752206862244e-12
C102_183 V102 V183 8.881171042659236e-20

R102_184 V102 V184 -2680.2894545896647
L102_184 V102 V184 8.983478151325995e-12
C102_184 V102 V184 -1.3388676167520552e-20

R102_185 V102 V185 -263.0458736688056
L102_185 V102 V185 -4.254753760701463e-12
C102_185 V102 V185 -7.335324354790127e-20

R102_186 V102 V186 205.42326991177626
L102_186 V102 V186 1.9522036919034494e-12
C102_186 V102 V186 3.264584870964647e-21

R102_187 V102 V187 1233.2909179318997
L102_187 V102 V187 -1.7010676104243908e-12
C102_187 V102 V187 -3.6334823757847915e-19

R102_188 V102 V188 -473.98386500411027
L102_188 V102 V188 -1.1233190202269758e-12
C102_188 V102 V188 -2.9578531048698205e-19

R102_189 V102 V189 638.3226175381997
L102_189 V102 V189 -2.112819960395784e-12
C102_189 V102 V189 -3.042371312490272e-19

R102_190 V102 V190 126.76906623780278
L102_190 V102 V190 -3.5507100719159847e-12
C102_190 V102 V190 3.0453881137087703e-19

R102_191 V102 V191 5273.1617676845035
L102_191 V102 V191 -1.1576418931575317e-12
C102_191 V102 V191 -2.9166688377287017e-19

R102_192 V102 V192 2980.109638164392
L102_192 V102 V192 -4.714902517133655e-12
C102_192 V102 V192 -1.65154908616822e-19

R102_193 V102 V193 455.669791035762
L102_193 V102 V193 2.5939840191317385e-12
C102_193 V102 V193 1.9937144090441304e-19

R102_194 V102 V194 -316.94913279902266
L102_194 V102 V194 2.677421745030234e-12
C102_194 V102 V194 8.984577517518739e-20

R102_195 V102 V195 -800.5722960273425
L102_195 V102 V195 9.101780142975791e-13
C102_195 V102 V195 5.673529104177202e-19

R102_196 V102 V196 -22261.41480598771
L102_196 V102 V196 1.3297902970322053e-12
C102_196 V102 V196 3.948045694148476e-19

R102_197 V102 V197 -283.7814031745373
L102_197 V102 V197 1.5110974750728808e-12
C102_197 V102 V197 2.3937409750087335e-19

R102_198 V102 V198 -147.99802702360054
L102_198 V102 V198 1.2262423721749155e-10
C102_198 V102 V198 -1.0815295811198042e-19

R102_199 V102 V199 -2561.779906269578
L102_199 V102 V199 1.7872995259965365e-12
C102_199 V102 V199 1.938814366305424e-19

R102_200 V102 V200 -4272.21712450005
L102_200 V102 V200 2.1370843774445014e-12
C102_200 V102 V200 9.39623898053858e-20

R103_103 V103 0 222.39551446755658
L103_103 V103 0 3.0437467026388874e-12
C103_103 V103 0 -2.2147242012158282e-20

R103_104 V103 V104 -511.63142009553695
L103_104 V103 V104 -7.36374249516974e-12
C103_104 V103 V104 1.2949697589474011e-20

R103_105 V103 V105 -461.64738098436015
L103_105 V103 V105 2.9005205196420456e-12
C103_105 V103 V105 1.4019694838512478e-19

R103_106 V103 V106 751.384340844344
L103_106 V103 V106 1.2110058816031215e-12
C103_106 V103 V106 3.6578652072840324e-19

R103_107 V103 V107 1218.290040097856
L103_107 V103 V107 4.4451812804364775e-12
C103_107 V103 V107 3.5732818873604906e-19

R103_108 V103 V108 476.1045529858388
L103_108 V103 V108 -1.287550452906309e-11
C103_108 V103 V108 -1.464326040949146e-19

R103_109 V103 V109 -958.0767142496586
L103_109 V103 V109 -4.725851367007918e-12
C103_109 V103 V109 -1.2507351737470508e-19

R103_110 V103 V110 505.7256476655131
L103_110 V103 V110 -1.6963380142525373e-12
C103_110 V103 V110 -2.642501198746665e-19

R103_111 V103 V111 131.276140024126
L103_111 V103 V111 8.384116576634924e-13
C103_111 V103 V111 4.593201319898239e-19

R103_112 V103 V112 611.1007826384812
L103_112 V103 V112 3.2035559398637435e-11
C103_112 V103 V112 2.3885829130286253e-20

R103_113 V103 V113 411.5702278308527
L103_113 V103 V113 -9.7404804612628e-12
C103_113 V103 V113 3.983590809885076e-20

R103_114 V103 V114 -709.1985694175834
L103_114 V103 V114 -1.6430799912278309e-12
C103_114 V103 V114 -2.5414890378682777e-19

R103_115 V103 V115 -252.99526761343333
L103_115 V103 V115 3.864793182766391e-12
C103_115 V103 V115 -2.8854483063011947e-19

R103_116 V103 V116 -383.762102781694
L103_116 V103 V116 1.5418890991072317e-11
C103_116 V103 V116 5.983051386290506e-20

R103_117 V103 V117 430.67297906155085
L103_117 V103 V117 2.969405995560325e-12
C103_117 V103 V117 5.75339576488764e-20

R103_118 V103 V118 -311.64534250996945
L103_118 V103 V118 1.4068207180720347e-12
C103_118 V103 V118 4.1794992107944073e-19

R103_119 V103 V119 -679.2151598667177
L103_119 V103 V119 -1.5382177022918398e-12
C103_119 V103 V119 6.778716350759171e-20

R103_120 V103 V120 -809.7440911029652
L103_120 V103 V120 6.640579277202998e-12
C103_120 V103 V120 1.195218925836442e-19

R103_121 V103 V121 -204.02048474546334
L103_121 V103 V121 -7.470572522584017e-12
C103_121 V103 V121 -1.6519812420367142e-19

R103_122 V103 V122 374.34479011424804
L103_122 V103 V122 5.571401875495914e-12
C103_122 V103 V122 3.7343505649382903e-20

R103_123 V103 V123 347.337151261071
L103_123 V103 V123 -1.4571780338962044e-12
C103_123 V103 V123 -4.021227562494582e-19

R103_124 V103 V124 313.33647993140175
L103_124 V103 V124 -3.7619273136894025e-12
C103_124 V103 V124 -1.9131718549883045e-19

R103_125 V103 V125 -293.8752047416768
L103_125 V103 V125 -1.0105379778224118e-11
C103_125 V103 V125 9.887816671514934e-20

R103_126 V103 V126 324.80354191208875
L103_126 V103 V126 -1.1781488027843395e-12
C103_126 V103 V126 -3.767820159838241e-19

R103_127 V103 V127 -582.8983436052307
L103_127 V103 V127 6.123630079999011e-13
C103_127 V103 V127 5.762713804420593e-19

R103_128 V103 V128 715.3272386811002
L103_128 V103 V128 -5.464147020035487e-12
C103_128 V103 V128 -1.4677943740296542e-19

R103_129 V103 V129 121.37457443182889
L103_129 V103 V129 4.65366765109128e-12
C103_129 V103 V129 -3.1820540387078345e-21

R103_130 V103 V130 -325.8068604597615
L103_130 V103 V130 9.152473223286704e-12
C103_130 V103 V130 7.84396295227704e-20

R103_131 V103 V131 466.005515981246
L103_131 V103 V131 -1.3286670627846078e-12
C103_131 V103 V131 -1.927408593000162e-19

R103_132 V103 V132 -245.42583996663106
L103_132 V103 V132 2.1489005172162088e-12
C103_132 V103 V132 4.1180203915018097e-19

R103_133 V103 V133 -2071.311203973623
L103_133 V103 V133 -4.765315111154432e-12
C103_133 V103 V133 -6.06358090286979e-20

R103_134 V103 V134 -421.9242087790102
L103_134 V103 V134 2.1221003484157e-12
C103_134 V103 V134 4.0092340479615425e-19

R103_135 V103 V135 2128.9630487104428
L103_135 V103 V135 -6.989532189164925e-13
C103_135 V103 V135 -9.034107430973065e-19

R103_136 V103 V136 -3776.245104810358
L103_136 V103 V136 -8.798410943329627e-12
C103_136 V103 V136 -5.67984975269446e-20

R103_137 V103 V137 -125.12425919147923
L103_137 V103 V137 -6.662477922556144e-12
C103_137 V103 V137 -3.5789858573740126e-20

R103_138 V103 V138 531.7463781518945
L103_138 V103 V138 -1.5590080460754609e-12
C103_138 V103 V138 -4.46424191221964e-19

R103_139 V103 V139 -163.38934187196224
L103_139 V103 V139 4.806780890716813e-13
C103_139 V103 V139 1.2942380451118446e-18

R103_140 V103 V140 6253.342224133213
L103_140 V103 V140 -2.6649825735403375e-11
C103_140 V103 V140 -4.2288426273449065e-20

R103_141 V103 V141 872.1516967659711
L103_141 V103 V141 1.5074034756941774e-11
C103_141 V103 V141 4.915220785201416e-20

R103_142 V103 V142 280.74212066910286
L103_142 V103 V142 -4.090015435641641e-12
C103_142 V103 V142 -1.1190157221058783e-19

R103_143 V103 V143 137.93867329229
L103_143 V103 V143 -4.9724200691028e-12
C103_143 V103 V143 -1.400489660327748e-19

R103_144 V103 V144 490.10694385700646
L103_144 V103 V144 5.3656722798968784e-11
C103_144 V103 V144 8.357295877432634e-20

R103_145 V103 V145 108.2030885791325
L103_145 V103 V145 1.0331334602239622e-11
C103_145 V103 V145 3.924728232318287e-21

R103_146 V103 V146 368.70756797919194
L103_146 V103 V146 1.3993378959669553e-12
C103_146 V103 V146 2.4387899549844065e-19

R103_147 V103 V147 246.51240896641838
L103_147 V103 V147 -9.954852508976177e-13
C103_147 V103 V147 -8.506806241819159e-19

R103_148 V103 V148 808.8107795480779
L103_148 V103 V148 1.885582293334758e-11
C103_148 V103 V148 -1.0708937727599522e-19

R103_149 V103 V149 -693.8259198953929
L103_149 V103 V149 7.620959801855953e-12
C103_149 V103 V149 -9.680790844282472e-20

R103_150 V103 V150 -124.36125139234734
L103_150 V103 V150 -4.3957411844940554e-12
C103_150 V103 V150 2.451605201056089e-19

R103_151 V103 V151 -87.82714797004354
L103_151 V103 V151 4.420004655266043e-11
C103_151 V103 V151 3.348895999793063e-19

R103_152 V103 V152 982.4332115410677
L103_152 V103 V152 2.0383050935651467e-11
C103_152 V103 V152 8.389605022708119e-21

R103_153 V103 V153 -115.8213970439807
L103_153 V103 V153 -2.972832823364966e-12
C103_153 V103 V153 -8.015123017368497e-20

R103_154 V103 V154 -223.90412565582227
L103_154 V103 V154 -5.0243851665255045e-12
C103_154 V103 V154 -3.1221241953350877e-19

R103_155 V103 V155 3197.3132148294694
L103_155 V103 V155 8.174870122958381e-13
C103_155 V103 V155 3.282695522315208e-19

R103_156 V103 V156 -190.03707084314772
L103_156 V103 V156 -4.467996528313905e-12
C103_156 V103 V156 -3.0235371645534096e-20

R103_157 V103 V157 -183.44658751280525
L103_157 V103 V157 8.931241179210188e-12
C103_157 V103 V157 2.1608583517822477e-19

R103_158 V103 V158 194.43870427160658
L103_158 V103 V158 -2.8482496819907137e-11
C103_158 V103 V158 9.995369145254609e-20

R103_159 V103 V159 93.50617369340183
L103_159 V103 V159 -1.401895131814687e-12
C103_159 V103 V159 -4.915913605325544e-19

R103_160 V103 V160 -1784.9369445408527
L103_160 V103 V160 -1.0929195859112226e-11
C103_160 V103 V160 2.0899235768932328e-20

R103_161 V103 V161 162.68955440763983
L103_161 V103 V161 1.9278442885884057e-12
C103_161 V103 V161 1.6698593170077576e-19

R103_162 V103 V162 188.10623869309924
L103_162 V103 V162 2.1159981261862283e-12
C103_162 V103 V162 1.2202248243705113e-19

R103_163 V103 V163 356.28250873935536
L103_163 V103 V163 -5.952147058073843e-12
C103_163 V103 V163 2.959657147102078e-19

R103_164 V103 V164 223.10813616016011
L103_164 V103 V164 3.708418385884611e-12
C103_164 V103 V164 7.716876223104144e-20

R103_165 V103 V165 257.8750670644352
L103_165 V103 V165 -1.4915879991229787e-12
C103_165 V103 V165 -3.8337311620815113e-19

R103_166 V103 V166 -161.14850801245274
L103_166 V103 V166 -4.6956700876963495e-12
C103_166 V103 V166 -1.0693193426081637e-19

R103_167 V103 V167 -75.91440601834735
L103_167 V103 V167 4.169728732104144e-12
C103_167 V103 V167 2.1175249234779618e-19

R103_168 V103 V168 272.4250640909199
L103_168 V103 V168 5.8164033613894495e-12
C103_168 V103 V168 6.61950426104409e-20

R103_169 V103 V169 -217.66796832491477
L103_169 V103 V169 -2.061736784023709e-12
C103_169 V103 V169 -1.7113602195794943e-19

R103_170 V103 V170 3725.8910435584644
L103_170 V103 V170 -3.338979441312584e-12
C103_170 V103 V170 -8.435399298404127e-20

R103_171 V103 V171 219.8387954897153
L103_171 V103 V171 -5.170972867082201e-11
C103_171 V103 V171 -4.965979365553713e-19

R103_172 V103 V172 -292.25630966492935
L103_172 V103 V172 -1.971185673914361e-12
C103_172 V103 V172 -1.8889861367648508e-19

R103_173 V103 V173 -1658.9931318763743
L103_173 V103 V173 1.1591045786088838e-12
C103_173 V103 V173 3.2396908741924495e-19

R103_174 V103 V174 286.8078668839434
L103_174 V103 V174 4.188335157174335e-12
C103_174 V103 V174 1.1444060881987374e-19

R103_175 V103 V175 162.38072064152465
L103_175 V103 V175 3.08452886376676e-12
C103_175 V103 V175 3.5593626599453117e-19

R103_176 V103 V176 -2284.4840363212325
L103_176 V103 V176 4.07405352705652e-12
C103_176 V103 V176 3.2765141476053255e-20

R103_177 V103 V177 753.0893699900802
L103_177 V103 V177 -4.013741864625806e-12
C103_177 V103 V177 -1.2282671992433442e-19

R103_178 V103 V178 -3263.519591981818
L103_178 V103 V178 8.283434276332155e-12
C103_178 V103 V178 3.583719257917273e-20

R103_179 V103 V179 -227.65646221348106
L103_179 V103 V179 -1.7269269254614555e-12
C103_179 V103 V179 -2.2596626827837315e-20

R103_180 V103 V180 762.4514610844261
L103_180 V103 V180 3.70623233663766e-12
C103_180 V103 V180 7.449418496620747e-20

R103_181 V103 V181 -1720.714351457208
L103_181 V103 V181 7.717243282915281e-12
C103_181 V103 V181 4.711969152449328e-21

R103_182 V103 V182 -344.24376869190996
L103_182 V103 V182 -3.365842720521688e-12
C103_182 V103 V182 -8.450846824977447e-20

R103_183 V103 V183 -435.580821429344
L103_183 V103 V183 8.269530023305535e-12
C103_183 V103 V183 1.7915953439536383e-20

R103_184 V103 V184 -836.6519796657959
L103_184 V103 V184 -2.441762046163698e-12
C103_184 V103 V184 -5.82840052212295e-20

R103_185 V103 V185 -756.7307043233903
L103_185 V103 V185 2.3847841236993657e-11
C103_185 V103 V185 8.384809549416912e-20

R103_186 V103 V186 -4480.5255407413415
L103_186 V103 V186 -3.344527134688623e-12
C103_186 V103 V186 -7.628773233412223e-20

R103_187 V103 V187 279.91022164701
L103_187 V103 V187 1.1387052521561684e-12
C103_187 V103 V187 1.9891801331549056e-19

R103_188 V103 V188 509.5117695265643
L103_188 V103 V188 2.8872253415057717e-12
C103_188 V103 V188 4.888876565520379e-21

R103_189 V103 V189 851.6081966102587
L103_189 V103 V189 -2.0677248345494164e-12
C103_189 V103 V189 -2.2464266892894347e-19

R103_190 V103 V190 577.7481373041992
L103_190 V103 V190 4.017187126227935e-12
C103_190 V103 V190 1.4637465099696572e-19

R103_191 V103 V191 537.6694280723433
L103_191 V103 V191 -1.323379370569231e-12
C103_191 V103 V191 -4.681406307611319e-19

R103_192 V103 V192 2557.611687482507
L103_192 V103 V192 1.8337024461677216e-11
C103_192 V103 V192 -1.3704175044541163e-19

R103_193 V103 V193 1017.0898174766021
L103_193 V103 V193 3.1602141206293916e-12
C103_193 V103 V193 8.420529781095537e-20

R103_194 V103 V194 -508.1434244074347
L103_194 V103 V194 -2.304398795032726e-12
C103_194 V103 V194 -2.0295004644610392e-19

R103_195 V103 V195 -379.34073690916654
L103_195 V103 V195 1.044525700585581e-12
C103_195 V103 V195 7.138312601956421e-19

R103_196 V103 V196 -467.7701382449457
L103_196 V103 V196 -2.3124890551658155e-12
C103_196 V103 V196 6.204561779732557e-20

R103_197 V103 V197 -679.0153478509782
L103_197 V103 V197 2.4156638079308777e-12
C103_197 V103 V197 1.5883117522178822e-19

R103_198 V103 V198 -650.8837876168051
L103_198 V103 V198 -4.804249508823254e-11
C103_198 V103 V198 -3.2720801785038272e-21

R103_199 V103 V199 -594.495919617063
L103_199 V103 V199 3.629891855264777e-12
C103_199 V103 V199 1.0417784819990312e-19

R103_200 V103 V200 1025.1386138056698
L103_200 V103 V200 1.6960418810174932e-12
C103_200 V103 V200 2.1793337679081613e-19

R104_104 V104 0 88.30946401324285
L104_104 V104 0 5.136256739187497e-13
C104_104 V104 0 1.0603158014942956e-18

R104_105 V104 V105 -450.7028209061792
L104_105 V104 V105 2.992799209979517e-12
C104_105 V104 V105 1.0414025005930106e-19

R104_106 V104 V106 430.4204820445126
L104_106 V104 V106 1.5179943723114558e-12
C104_106 V104 V106 2.543239611377003e-19

R104_107 V104 V107 433.36748872521326
L104_107 V104 V107 -4.7224089623493934e-12
C104_107 V104 V107 -1.1921969412753273e-19

R104_108 V104 V108 7866.935003431216
L104_108 V104 V108 1.1589608305776922e-12
C104_108 V104 V108 5.112241025725244e-19

R104_109 V104 V109 -518.0823927444325
L104_109 V104 V109 -3.1528255494628874e-12
C104_109 V104 V109 -1.7516040299258697e-19

R104_110 V104 V110 777.8884829237047
L104_110 V104 V110 -1.7462833857559214e-12
C104_110 V104 V110 -2.288507005856622e-19

R104_111 V104 V111 441.39339380105736
L104_111 V104 V111 -4.479214017554954e-10
C104_111 V104 V111 3.517057412757665e-20

R104_112 V104 V112 140.17422800751373
L104_112 V104 V112 2.1343139573268176e-12
C104_112 V104 V112 1.6453653600124739e-19

R104_113 V104 V113 257.45532497440706
L104_113 V104 V113 -1.0604361036066313e-11
C104_113 V104 V113 8.045593972824862e-20

R104_114 V104 V114 -739.1530172217125
L104_114 V104 V114 -1.6857092353518954e-12
C104_114 V104 V114 -1.797746772051357e-19

R104_115 V104 V115 -272.4160063628813
L104_115 V104 V115 1.3274986799301263e-11
C104_115 V104 V115 6.572965772731341e-20

R104_116 V104 V116 -363.47162989132795
L104_116 V104 V116 7.990497376317807e-12
C104_116 V104 V116 -2.5140314653669907e-19

R104_117 V104 V117 347.3244337109372
L104_117 V104 V117 2.5137500309325675e-12
C104_117 V104 V117 9.109051513001276e-20

R104_118 V104 V118 -273.2112279422893
L104_118 V104 V118 1.8523506982823856e-12
C104_118 V104 V118 3.3331982190941395e-19

R104_119 V104 V119 -689.7008372457304
L104_119 V104 V119 3.3441258623751626e-12
C104_119 V104 V119 2.200492982313527e-19

R104_120 V104 V120 -263.89250111334223
L104_120 V104 V120 -1.5547829270002422e-11
C104_120 V104 V120 4.807201520452958e-19

R104_121 V104 V121 -152.63579396156172
L104_121 V104 V121 -5.5696200099390745e-12
C104_121 V104 V121 -1.9739184638009547e-19

R104_122 V104 V122 432.290757477294
L104_122 V104 V122 4.7814946930778735e-12
C104_122 V104 V122 1.1466926227913474e-19

R104_123 V104 V123 290.184576186497
L104_123 V104 V123 -2.305940117650841e-12
C104_123 V104 V123 -2.1428116032305262e-19

R104_124 V104 V124 232.48602968345432
L104_124 V104 V124 -7.185846740539001e-13
C104_124 V104 V124 -8.35918617555968e-19

R104_125 V104 V125 -267.49295823533555
L104_125 V104 V125 -3.62981803945551e-12
C104_125 V104 V125 5.092351640593306e-20

R104_126 V104 V126 238.35384650192623
L104_126 V104 V126 -1.0441938433305871e-12
C104_126 V104 V126 -3.701247799253826e-19

R104_127 V104 V127 820.6760524202642
L104_127 V104 V127 -1.4581935014239937e-12
C104_127 V104 V127 -2.859907783497507e-19

R104_128 V104 V128 1334.6909276409076
L104_128 V104 V128 6.935111629544159e-13
C104_128 V104 V128 3.446667135923281e-19

R104_129 V104 V129 98.2522473625463
L104_129 V104 V129 2.6573872406161908e-12
C104_129 V104 V129 3.912827984971658e-21

R104_130 V104 V130 -269.15707708380796
L104_130 V104 V130 5.77825125389488e-12
C104_130 V104 V130 1.0162748801085548e-19

R104_131 V104 V131 -256.68963110957526
L104_131 V104 V131 1.187639869999467e-12
C104_131 V104 V131 4.619588699298701e-19

R104_132 V104 V132 -580.6622895354933
L104_132 V104 V132 -2.7648943129827718e-12
C104_132 V104 V132 1.94811301314105e-19

R104_133 V104 V133 -1384.6200179662435
L104_133 V104 V133 -6.283585733907099e-12
C104_133 V104 V133 4.404618172010012e-20

R104_134 V104 V134 -308.204477451863
L104_134 V104 V134 1.6549090626797566e-12
C104_134 V104 V134 5.6366310396957525e-19

R104_135 V104 V135 -3124.2013577734015
L104_135 V104 V135 -6.1653571052685515e-12
C104_135 V104 V135 -1.8616311210999725e-20

R104_136 V104 V136 1872.6310094178982
L104_136 V104 V136 -6.852314106070823e-13
C104_136 V104 V136 -8.49381578760479e-19

R104_137 V104 V137 -112.21471806493332
L104_137 V104 V137 -2.3807277727474236e-12
C104_137 V104 V137 -1.2004493087807927e-19

R104_138 V104 V138 301.7140823568422
L104_138 V104 V138 -1.1938035851027212e-12
C104_138 V104 V138 -5.625567766277531e-19

R104_139 V104 V139 764.7054528035405
L104_139 V104 V139 -3.95593012043026e-12
C104_139 V104 V139 -1.785035652901588e-19

R104_140 V104 V140 -187.11873410767353
L104_140 V104 V140 6.033569768286614e-13
C104_140 V104 V140 1.0757633766862798e-18

R104_141 V104 V141 2705.6221910631007
L104_141 V104 V141 4.247448865549388e-11
C104_141 V104 V141 3.4859621348873214e-20

R104_142 V104 V142 292.83093818532706
L104_142 V104 V142 -3.013645897122171e-12
C104_142 V104 V142 -1.3995274446163213e-19

R104_143 V104 V143 876.6035078498337
L104_143 V104 V143 -1.0439991636609217e-11
C104_143 V104 V143 1.1009795320074958e-19

R104_144 V104 V144 119.87919989369946
L104_144 V104 V144 -4.2466668805845014e-12
C104_144 V104 V144 -2.1060260622493782e-19

R104_145 V104 V145 94.72987619430617
L104_145 V104 V145 3.4968830952267697e-12
C104_145 V104 V145 5.152676773859616e-20

R104_146 V104 V146 327.6511256724147
L104_146 V104 V146 1.1153237675780403e-12
C104_146 V104 V146 2.746732918713532e-19

R104_147 V104 V147 261.24528434809895
L104_147 V104 V147 -5.9953548940384074e-12
C104_147 V104 V147 -2.213883534483328e-19

R104_148 V104 V148 -1208.0699923910242
L104_148 V104 V148 -7.933921930267277e-13
C104_148 V104 V148 -5.761055815680476e-19

R104_149 V104 V149 -3779.3645899314974
L104_149 V104 V149 1.4125378037872335e-11
C104_149 V104 V149 -2.242591821671659e-19

R104_150 V104 V150 -108.82536093002426
L104_150 V104 V150 -3.7306481782941464e-12
C104_150 V104 V150 1.7042497197200736e-19

R104_151 V104 V151 -292.39313103329687
L104_151 V104 V151 4.176683516835007e-12
C104_151 V104 V151 -1.7995194683138263e-20

R104_152 V104 V152 -218.39164875568153
L104_152 V104 V152 1.638312778311927e-12
C104_152 V104 V152 2.315961314842502e-19

R104_153 V104 V153 -97.75273083982326
L104_153 V104 V153 -1.1025894351417275e-11
C104_153 V104 V153 2.693505618783023e-20

R104_154 V104 V154 -209.16306413317358
L104_154 V104 V154 2.992780725876768e-11
C104_154 V104 V154 -2.880971972847044e-19

R104_155 V104 V155 2868.8303737501383
L104_155 V104 V155 3.4574548720025915e-12
C104_155 V104 V155 1.512085357801327e-20

R104_156 V104 V156 -98.27533606660569
L104_156 V104 V156 2.973378160406955e-12
C104_156 V104 V156 4.676534171928383e-19

R104_157 V104 V157 -139.57085067194376
L104_157 V104 V157 -4.753937969258192e-12
C104_157 V104 V157 1.6073407368837572e-19

R104_158 V104 V158 192.30427104049843
L104_158 V104 V158 -7.24873406287075e-12
C104_158 V104 V158 9.474706373352365e-20

R104_159 V104 V159 -301.0989624723302
L104_159 V104 V159 -4.779779726569392e-12
C104_159 V104 V159 4.5865081530857335e-20

R104_160 V104 V160 72.44804811371519
L104_160 V104 V160 -5.828377074919059e-12
C104_160 V104 V160 -4.210046239207128e-19

R104_161 V104 V161 135.90056329034107
L104_161 V104 V161 1.0943986886820747e-12
C104_161 V104 V161 1.6503330122473378e-19

R104_162 V104 V162 168.78007239938685
L104_162 V104 V162 1.6882205965833115e-12
C104_162 V104 V162 1.1244057183399387e-19

R104_163 V104 V163 221.99239354603068
L104_163 V104 V163 1.9682469866378824e-12
C104_163 V104 V163 1.3066119686288364e-19

R104_164 V104 V164 211.4040489088037
L104_164 V104 V164 -5.195324303183819e-12
C104_164 V104 V164 2.3425554732866357e-19

R104_165 V104 V165 219.47965390309457
L104_165 V104 V165 -1.5196482810544818e-12
C104_165 V104 V165 -3.9979866273044724e-19

R104_166 V104 V166 -142.0526570111752
L104_166 V104 V166 -5.182469896866337e-12
C104_166 V104 V166 -1.6890437577432873e-19

R104_167 V104 V167 1225.7443581137743
L104_167 V104 V167 1.3625664316587109e-11
C104_167 V104 V167 2.4839237161636585e-20

R104_168 V104 V168 -88.96863180212166
L104_168 V104 V168 1.8089240690271304e-12
C104_168 V104 V168 1.560256410068831e-19

R104_169 V104 V169 -164.51444639694557
L104_169 V104 V169 -2.1368357864685603e-12
C104_169 V104 V169 -1.7149464578729927e-19

R104_170 V104 V170 -1157.8365436615968
L104_170 V104 V170 -6.17489741127432e-12
C104_170 V104 V170 -7.340265876657683e-20

R104_171 V104 V171 -474.68927013052695
L104_171 V104 V171 -4.364352791390424e-12
C104_171 V104 V171 -2.432418056034856e-19

R104_172 V104 V172 1890.0534809478195
L104_172 V104 V172 -2.008913070130132e-12
C104_172 V104 V172 -3.4489682793402115e-19

R104_173 V104 V173 -1553.7017328869695
L104_173 V104 V173 1.1312636057858445e-12
C104_173 V104 V173 3.607641102208875e-19

R104_174 V104 V174 252.55066456937297
L104_174 V104 V174 8.544433579002126e-12
C104_174 V104 V174 1.4808361351851265e-19

R104_175 V104 V175 -878.4022667436474
L104_175 V104 V175 1.5071402883123866e-11
C104_175 V104 V175 7.053586085829826e-20

R104_176 V104 V176 135.47522485431526
L104_176 V104 V176 2.4541296093773624e-12
C104_176 V104 V176 4.0513359448738146e-19

R104_177 V104 V177 423.00072173731303
L104_177 V104 V177 -6.5093168941772335e-12
C104_177 V104 V177 -1.5899258985189813e-19

R104_178 V104 V178 875.9209432379912
L104_178 V104 V178 1.1921328776558946e-11
C104_178 V104 V178 1.6098337599461738e-20

R104_179 V104 V179 375.73083382545445
L104_179 V104 V179 6.218616242209124e-12
C104_179 V104 V179 7.069786955882477e-20

R104_180 V104 V180 -357.79463738390035
L104_180 V104 V180 -1.3518997367708665e-12
C104_180 V104 V180 -1.1277220704653568e-19

R104_181 V104 V181 -787.8677708260468
L104_181 V104 V181 6.715930234505187e-11
C104_181 V104 V181 -3.324403377284555e-20

R104_182 V104 V182 -234.6394752725133
L104_182 V104 V182 -3.0438204489465165e-12
C104_182 V104 V182 -1.5053154709117333e-19

R104_183 V104 V183 -610.3594750748862
L104_183 V104 V183 -2.3065895513963696e-12
C104_183 V104 V183 -5.481225021156328e-20

R104_184 V104 V184 -381.8802893292031
L104_184 V104 V184 4.8618404858412644e-11
C104_184 V104 V184 -1.4657926876936543e-20

R104_185 V104 V185 -539.6609811284569
L104_185 V104 V185 1.40721030786903e-11
C104_185 V104 V185 1.2786967035873063e-19

R104_186 V104 V186 -959.486326827277
L104_186 V104 V186 -2.5551975928711904e-12
C104_186 V104 V186 -2.0241289567046047e-20

R104_187 V104 V187 7652.168392927576
L104_187 V104 V187 -1.717307423665823e-11
C104_187 V104 V187 1.1193265123261618e-20

R104_188 V104 V188 229.9050113086577
L104_188 V104 V188 6.268446699625981e-13
C104_188 V104 V188 1.279211039559257e-19

R104_189 V104 V189 740.7253703382389
L104_189 V104 V189 -2.2884542650748267e-12
C104_189 V104 V189 -2.172927258271841e-19

R104_190 V104 V190 453.6652876214923
L104_190 V104 V190 2.8554342217879823e-12
C104_190 V104 V190 1.4547663024993078e-19

R104_191 V104 V191 835.7858623203025
L104_191 V104 V191 1.5403238600815802e-12
C104_191 V104 V191 -7.052995578454051e-20

R104_192 V104 V192 799.7224320569229
L104_192 V104 V192 -6.656621110185311e-13
C104_192 V104 V192 -4.795157037760843e-19

R104_193 V104 V193 609.0626748103318
L104_193 V104 V193 6.203896599981234e-12
C104_193 V104 V193 3.3710197024911077e-20

R104_194 V104 V194 -466.4478582552616
L104_194 V104 V194 -1.4600345123769488e-12
C104_194 V104 V194 -2.8491232911167057e-19

R104_195 V104 V195 -537.4015873117711
L104_195 V104 V195 -1.2590524964046447e-12
C104_195 V104 V195 -8.621188270827277e-20

R104_196 V104 V196 -348.403806122924
L104_196 V104 V196 5.693078038663046e-13
C104_196 V104 V196 9.354583748923098e-19

R104_197 V104 V197 -652.1946748233586
L104_197 V104 V197 2.5325822144204163e-12
C104_197 V104 V197 1.5769595889504335e-19

R104_198 V104 V198 -388.8534102800698
L104_198 V104 V198 -1.7552380474857724e-11
C104_198 V104 V198 -8.685151263495624e-20

R104_199 V104 V199 -1060.9050359674773
L104_199 V104 V199 1.8292730310994865e-12
C104_199 V104 V199 2.4193557387666603e-19

R104_200 V104 V200 -6192.2929352515885
L104_200 V104 V200 1.975929130621398e-11
C104_200 V104 V200 -8.893066339744987e-20

R105_105 V105 0 29.899757826432275
L105_105 V105 0 6.835683176978814e-13
C105_105 V105 0 -1.2758031664841658e-18

R105_106 V105 V106 -391.2473126329775
L105_106 V105 V106 -3.3705180641001863e-12
C105_106 V105 V106 -1.3055673686697617e-19

R105_107 V105 V107 171.7768790521696
L105_107 V105 V107 2.19264952375527e-12
C105_107 V105 V107 1.716443320125613e-19

R105_108 V105 V108 146.8692734381728
L105_108 V105 V108 -7.532410322984796e-12
C105_108 V105 V108 -3.9769900245132925e-20

R105_109 V105 V109 804.6288622233074
L105_109 V105 V109 3.232035599146024e-12
C105_109 V105 V109 2.670597508183529e-19

R105_110 V105 V110 167.36414108114437
L105_110 V105 V110 1.1151344243512898e-11
C105_110 V105 V110 6.434666029785467e-20

R105_111 V105 V111 -780.3069962408515
L105_111 V105 V111 -3.937234430921506e-12
C105_111 V105 V111 -1.4129235207754645e-20

R105_112 V105 V112 -660.7843046689549
L105_112 V105 V112 6.408988572946572e-12
C105_112 V105 V112 1.4756758474971777e-19

R105_113 V105 V113 47.39020593814324
L105_113 V105 V113 9.269109393198812e-13
C105_113 V105 V113 5.20970545625579e-19

R105_114 V105 V114 470.34447127484344
L105_114 V105 V114 1.8226073673329475e-12
C105_114 V105 V114 2.584665319607036e-19

R105_115 V105 V115 -240.55246927529112
L105_115 V105 V115 -2.2914188039811796e-12
C105_115 V105 V115 -1.673837474810994e-19

R105_116 V105 V116 -175.80749014088997
L105_116 V105 V116 -5.310239647528032e-12
C105_116 V105 V116 -3.453174707022327e-21

R105_117 V105 V117 -100.91812147691482
L105_117 V105 V117 -7.368946335158698e-12
C105_117 V105 V117 -1.4436599718201524e-19

R105_118 V105 V118 -87.63887865535129
L105_118 V105 V118 -1.2895908886232716e-12
C105_118 V105 V118 -3.445060125589655e-19

R105_119 V105 V119 384.6442436509217
L105_119 V105 V119 1.1092322687201576e-11
C105_119 V105 V119 -1.356619503049773e-19

R105_120 V105 V120 150.53780044804068
L105_120 V105 V120 -6.02389397568726e-12
C105_120 V105 V120 -3.4041218373052114e-19

R105_121 V105 V121 -87.75253055383577
L105_121 V105 V121 -1.0321235807826283e-12
C105_121 V105 V121 -3.0241817513726223e-19

R105_122 V105 V122 182.67953766568948
L105_122 V105 V122 4.152445754374269e-12
C105_122 V105 V122 1.0522959870955803e-19

R105_123 V105 V123 -10910.987176698674
L105_123 V105 V123 2.14338629177036e-12
C105_123 V105 V123 3.297411328235312e-19

R105_124 V105 V124 -422.0085379749916
L105_124 V105 V124 1.5939030730752483e-12
C105_124 V105 V124 4.508432939250723e-19

R105_125 V105 V125 -947.8937861990019
L105_125 V105 V125 -2.8165022147566235e-10
C105_125 V105 V125 5.318873295482924e-20

R105_126 V105 V126 93.74353033229943
L105_126 V105 V126 1.5168553572837264e-12
C105_126 V105 V126 1.9337303566339663e-19

R105_127 V105 V127 283.468357588467
L105_127 V105 V127 -1.2720802373429479e-11
C105_127 V105 V127 -3.074173542573676e-20

R105_128 V105 V128 4146.28889206312
L105_128 V105 V128 -3.7173931068137286e-12
C105_128 V105 V128 2.45523584623426e-20

R105_129 V105 V129 95.53175035118925
L105_129 V105 V129 1.3204623589226108e-12
C105_129 V105 V129 3.1076224594177195e-19

R105_130 V105 V130 -125.88068887162994
L105_130 V105 V130 -1.461028522813613e-12
C105_130 V105 V130 -2.7260487799665255e-19

R105_131 V105 V131 -211.71938780385935
L105_131 V105 V131 -3.3405872087981636e-12
C105_131 V105 V131 -1.8930164302847334e-19

R105_132 V105 V132 -685.185698570108
L105_132 V105 V132 -2.4270302492158507e-12
C105_132 V105 V132 -4.276734465389125e-19

R105_133 V105 V133 370.7581275801671
L105_133 V105 V133 -1.6939056978764932e-12
C105_133 V105 V133 -3.034322632648239e-19

R105_134 V105 V134 -2526.0570287144033
L105_134 V105 V134 2.5074704722441427e-12
C105_134 V105 V134 1.159141276856141e-19

R105_135 V105 V135 -198.3687196415836
L105_135 V105 V135 7.978308265404845e-12
C105_135 V105 V135 2.1650483488417555e-19

R105_136 V105 V136 -131.30660190718677
L105_136 V105 V136 2.8741614251706443e-12
C105_136 V105 V136 3.7252501139046066e-19

R105_137 V105 V137 -70.58514412466602
L105_137 V105 V137 1.1765358405074389e-11
C105_137 V105 V137 8.373006805742975e-20

R105_138 V105 V138 531.9211539966672
L105_138 V105 V138 8.376374188618522e-12
C105_138 V105 V138 1.0960770559799338e-19

R105_139 V105 V139 87.25298259624559
L105_139 V105 V139 -4.396302226136875e-12
C105_139 V105 V139 -3.0346391129574744e-19

R105_140 V105 V140 71.20439262287172
L105_140 V105 V140 2.987339515650026e-11
C105_140 V105 V140 -2.268274409415994e-19

R105_141 V105 V141 -355.95617925928497
L105_141 V105 V141 3.3142769057011922e-12
C105_141 V105 V141 2.730830908268793e-19

R105_142 V105 V142 222.44297288567026
L105_142 V105 V142 -2.1179645577699327e-12
C105_142 V105 V142 -1.1821558912212732e-19

R105_143 V105 V143 -3568.040037863712
L105_143 V105 V143 2.2454848034812104e-12
C105_143 V105 V143 1.6331065508521772e-19

R105_144 V105 V144 467.84370555771727
L105_144 V105 V144 -1.4499579265956651e-11
C105_144 V105 V144 -5.956927395129359e-20

R105_145 V105 V145 110.14677288785943
L105_145 V105 V145 -1.4639112079789834e-11
C105_145 V105 V145 -1.3258305275497724e-20

R105_146 V105 V146 799.3236466904334
L105_146 V105 V146 2.9079259834478783e-12
C105_146 V105 V146 -4.5724701343144844e-20

R105_147 V105 V147 -239.2630904484866
L105_147 V105 V147 -7.134133418179843e-11
C105_147 V105 V147 2.1792265121926643e-19

R105_148 V105 V148 -103.55610490485768
L105_148 V105 V148 4.768577485978105e-12
C105_148 V105 V148 2.3356761728843626e-19

R105_149 V105 V149 89.76371536641506
L105_149 V105 V149 -1.027756232735812e-12
C105_149 V105 V149 -5.854500152160892e-19

R105_150 V105 V150 -76.78027562060491
L105_150 V105 V150 -1.4602267623125098e-11
C105_150 V105 V150 2.1590408797448247e-19

R105_151 V105 V151 -203.38984849859872
L105_151 V105 V151 -2.0486261916346822e-12
C105_151 V105 V151 -2.1334654149973822e-19

R105_152 V105 V152 343.76545730528846
L105_152 V105 V152 -4.581361003171859e-12
C105_152 V105 V152 -1.4483947138420653e-20

R105_153 V105 V153 -72.78455915290617
L105_153 V105 V153 4.214486571543701e-12
C105_153 V105 V153 1.5992468431715908e-19

R105_154 V105 V154 -753.2899184565298
L105_154 V105 V154 -2.3995148248543836e-11
C105_154 V105 V154 -9.55730348406074e-20

R105_155 V105 V155 140.9515393025959
L105_155 V105 V155 -2.708125526109067e-12
C105_155 V105 V155 -1.9755494731011524e-19

R105_156 V105 V156 -242.04206779668232
L105_156 V105 V156 4.830531758718708e-11
C105_156 V105 V156 -1.6338868348586122e-19

R105_157 V105 V157 -53.916785399055485
L105_157 V105 V157 1.0758288632055392e-12
C105_157 V105 V157 6.033028493415663e-19

R105_158 V105 V158 194.30431995352103
L105_158 V105 V158 -1.0622833944665529e-11
C105_158 V105 V158 3.887208530375233e-20

R105_159 V105 V159 -335.45823941360754
L105_159 V105 V159 1.6623143902768572e-12
C105_159 V105 V159 2.202369910489899e-19

R105_160 V105 V160 300.1448623142967
L105_160 V105 V160 2.8929847867038584e-12
C105_160 V105 V160 1.013801269274923e-19

R105_161 V105 V161 114.29168572768062
L105_161 V105 V161 -1.7916540506344749e-12
C105_161 V105 V161 -2.7747701701526334e-19

R105_162 V105 V162 104.646752053576
L105_162 V105 V162 -5.934012555365306e-12
C105_162 V105 V162 -1.2014333675674763e-19

R105_163 V105 V163 89.36766986489637
L105_163 V105 V163 2.454445764031332e-12
C105_163 V105 V163 2.05959018031443e-20

R105_164 V105 V164 100.19066481886782
L105_164 V105 V164 8.409025071757583e-12
C105_164 V105 V164 -1.612911462545706e-19

R105_165 V105 V165 191.66097338052754
L105_165 V105 V165 -1.608237990318036e-12
C105_165 V105 V165 -1.1509021530652795e-19

R105_166 V105 V166 -182.74035729301184
L105_166 V105 V166 -6.265078977920698e-12
C105_166 V105 V166 -4.325537999133911e-20

R105_167 V105 V167 -241.44570090884505
L105_167 V105 V167 -2.403695996953098e-12
C105_167 V105 V167 -9.824772289243023e-20

R105_168 V105 V168 625.7267151074105
L105_168 V105 V168 -1.9379680905585736e-12
C105_168 V105 V168 -4.9406306092703813e-20

R105_169 V105 V169 -82.17913986059435
L105_169 V105 V169 1.5979490328588046e-12
C105_169 V105 V169 4.29982855552861e-19

R105_170 V105 V170 -91.56603156105875
L105_170 V105 V170 -4.038338129820532e-12
C105_170 V105 V170 -4.17680282554681e-20

R105_171 V105 V171 -97.8344665696844
L105_171 V105 V171 -1.2428588357622817e-12
C105_171 V105 V171 -1.3917818856533287e-19

R105_172 V105 V172 -87.97696279463038
L105_172 V105 V172 -7.1286148042222245e-12
C105_172 V105 V172 1.964499720288146e-20

R105_173 V105 V173 -258.86117298934283
L105_173 V105 V173 7.063510432351114e-12
C105_173 V105 V173 -1.6330733346233475e-19

R105_174 V105 V174 93.86449105456089
L105_174 V105 V174 1.4740935863745532e-12
C105_174 V105 V174 3.0866375649551393e-19

R105_175 V105 V175 142.88466902502967
L105_175 V105 V175 2.0022942899605186e-12
C105_175 V105 V175 -5.623865119262233e-20

R105_176 V105 V176 134.8838389300797
L105_176 V105 V176 1.9871799739511144e-12
C105_176 V105 V176 -7.894585541142813e-20

R105_177 V105 V177 138.96519369018944
L105_177 V105 V177 -2.353649568115505e-12
C105_177 V105 V177 -2.1752098844633866e-19

R105_178 V105 V178 284.51067334362483
L105_178 V105 V178 4.575395909678347e-12
C105_178 V105 V178 -8.90421450437368e-21

R105_179 V105 V179 203.16473187514052
L105_179 V105 V179 1.5626638922197112e-12
C105_179 V105 V179 3.1731583584686853e-19

R105_180 V105 V180 144.27622841209762
L105_180 V105 V180 2.126777885667152e-12
C105_180 V105 V180 2.3060777496634715e-19

R105_181 V105 V181 -253.34766202121472
L105_181 V105 V181 -6.5719724140499326e-12
C105_181 V105 V181 1.0025542000155288e-19

R105_182 V105 V182 -90.31857603959894
L105_182 V105 V182 -1.0253294453529459e-12
C105_182 V105 V182 -1.6471862108677352e-19

R105_183 V105 V183 -164.5743156097228
L105_183 V105 V183 8.251061399114149e-12
C105_183 V105 V183 9.732877745942905e-20

R105_184 V105 V184 -128.72391841222137
L105_184 V105 V184 -7.722085364519032e-12
C105_184 V105 V184 -1.4721872621648205e-20

R105_185 V105 V185 -131.13916366401082
L105_185 V105 V185 9.282202036938156e-12
C105_185 V105 V185 1.2620452667155348e-19

R105_186 V105 V186 642.9621283654325
L105_186 V105 V186 -3.3128623818863778e-12
C105_186 V105 V186 -1.744283474564953e-20

R105_187 V105 V187 347.8279592248498
L105_187 V105 V187 -1.4185368373864342e-12
C105_187 V105 V187 -3.407237466164725e-19

R105_188 V105 V188 615.4771787995265
L105_188 V105 V188 -9.39089336510824e-13
C105_188 V105 V188 -2.6405858326192627e-19

R105_189 V105 V189 85.4409271376755
L105_189 V105 V189 2.7401760970962878e-12
C105_189 V105 V189 -1.412223755296379e-19

R105_190 V105 V190 193.69730581987753
L105_190 V105 V190 1.829036701200829e-12
C105_190 V105 V190 1.3057719649835658e-19

R105_191 V105 V191 972.692084238511
L105_191 V105 V191 -2.9880291232128796e-12
C105_191 V105 V191 -1.3641033889158856e-19

R105_192 V105 V192 222.52942972372097
L105_192 V105 V192 1.8720360250513174e-12
C105_192 V105 V192 2.6219924034224872e-20

R105_193 V105 V193 561.3462964316811
L105_193 V105 V193 5.921521728896021e-12
C105_193 V105 V193 1.532110929161527e-19

R105_194 V105 V194 -144.44152152340715
L105_194 V105 V194 1.5734942903363808e-12
C105_194 V105 V194 3.2715891594370015e-19

R105_195 V105 V195 -258.6559362186879
L105_195 V105 V195 1.3090638354747477e-12
C105_195 V105 V195 2.970545218350437e-19

R105_196 V105 V196 -171.60689414397757
L105_196 V105 V196 1.5478580534540087e-12
C105_196 V105 V196 1.5445532838630124e-19

R105_197 V105 V197 -105.70444920785009
L105_197 V105 V197 -2.7825328654172175e-12
C105_197 V105 V197 -1.0111164294856182e-19

R105_198 V105 V198 -261.25746325408073
L105_198 V105 V198 -1.6810071649298024e-12
C105_198 V105 V198 -6.909165178866799e-20

R105_199 V105 V199 -10392.866813926965
L105_199 V105 V199 -9.75908714003906e-12
C105_199 V105 V199 1.2401967819429058e-19

R105_200 V105 V200 649.2531809784382
L105_200 V105 V200 -1.6792812922857116e-12
C105_200 V105 V200 -4.7075069306382437e-20

R106_106 V106 0 53.67345383747519
L106_106 V106 0 -6.618280766391376e-13
C106_106 V106 0 -9.38479169260373e-19

R106_107 V106 V107 1948.3443630281333
L106_107 V106 V107 1.6946324865369296e-12
C106_107 V106 V107 3.021479616844253e-19

R106_108 V106 V108 907.7612452533375
L106_108 V106 V108 2.2028273361048914e-11
C106_108 V106 V108 8.118865967260537e-20

R106_109 V106 V109 223.7900017921446
L106_109 V106 V109 3.846346402622652e-12
C106_109 V106 V109 3.6396631890421056e-19

R106_110 V106 V110 109.43915775940157
L106_110 V106 V110 2.5022217612284094e-12
C106_110 V106 V110 1.6840487950194684e-19

R106_111 V106 V111 -169.65619192340705
L106_111 V106 V111 -4.898858297379894e-12
C106_111 V106 V111 -2.1328147803180265e-20

R106_112 V106 V112 -184.4993684674875
L106_112 V106 V112 6.051563026024911e-12
C106_112 V106 V112 2.1980251652521233e-19

R106_113 V106 V113 747.5320251493125
L106_113 V106 V113 1.3105709128638211e-11
C106_113 V106 V113 -1.6300631065704135e-19

R106_114 V106 V114 62.89405149812103
L106_114 V106 V114 6.047645205161657e-13
C106_114 V106 V114 9.241351456902366e-19

R106_115 V106 V115 197.63818158514593
L106_115 V106 V115 -1.422831330333871e-12
C106_115 V106 V115 -2.198949901946985e-19

R106_116 V106 V116 275.39185246315316
L106_116 V106 V116 -1.925283659427337e-12
C106_116 V106 V116 -1.6969043111890067e-19

R106_117 V106 V117 -153.41321119141347
L106_117 V106 V117 -3.791663417830358e-12
C106_117 V106 V117 1.3255941225958667e-20

R106_118 V106 V118 -41.75737866365526
L106_118 V106 V118 -1.1723978768148972e-12
C106_118 V106 V118 -2.8207568133654477e-19

R106_119 V106 V119 2651.018898673454
L106_119 V106 V119 -3.2317250686526434e-11
C106_119 V106 V119 -2.73576906898928e-19

R106_120 V106 V120 386.1600367199174
L106_120 V106 V120 -4.6960773450484666e-12
C106_120 V106 V120 -4.413152920191894e-19

R106_121 V106 V121 200.08034848372878
L106_121 V106 V121 3.6245411702161727e-12
C106_121 V106 V121 1.7751344159420175e-19

R106_122 V106 V122 347.1071642053252
L106_122 V106 V122 -1.4107556378853816e-12
C106_122 V106 V122 -5.338169724448325e-19

R106_123 V106 V123 -135.94085881836756
L106_123 V106 V123 8.949142831844383e-13
C106_123 V106 V123 7.739198137002964e-19

R106_124 V106 V124 -124.7502667591686
L106_124 V106 V124 8.614990810146969e-13
C106_124 V106 V124 8.67470506369867e-19

R106_125 V106 V125 317.79067227782366
L106_125 V106 V125 -1.4905557279723087e-11
C106_125 V106 V125 -2.430808362427243e-19

R106_126 V106 V126 53.47808566306085
L106_126 V106 V126 9.170148250632507e-13
C106_126 V106 V126 1.5322309950891608e-19

R106_127 V106 V127 124.06222282215323
L106_127 V106 V127 -2.6250904819406265e-12
C106_127 V106 V127 -2.605358080592642e-19

R106_128 V106 V128 171.251462321325
L106_128 V106 V128 -2.5923410046986294e-12
C106_128 V106 V128 -1.3641051394708768e-19

R106_129 V106 V129 -157.74410125157053
L106_129 V106 V129 -2.9122977538824436e-12
C106_129 V106 V129 5.793826603608206e-20

R106_130 V106 V130 -90.12353354856276
L106_130 V106 V130 -2.8086667115596302e-11
C106_130 V106 V130 3.5214561684698273e-19

R106_131 V106 V131 -214.73130427598372
L106_131 V106 V131 -1.832053143429061e-12
C106_131 V106 V131 -3.314258319114538e-19

R106_132 V106 V132 -257.7014518295857
L106_132 V106 V132 -1.325624395215483e-12
C106_132 V106 V132 -5.508997650587955e-19

R106_133 V106 V133 402.50458705524744
L106_133 V106 V133 3.029614524838949e-12
C106_133 V106 V133 6.977738791108077e-20

R106_134 V106 V134 -172.49334322980818
L106_134 V106 V134 -1.2835820407764334e-12
C106_134 V106 V134 -6.059877316581306e-19

R106_135 V106 V135 -136.0667133332822
L106_135 V106 V135 1.1908398640847869e-12
C106_135 V106 V135 7.677755856730114e-19

R106_136 V106 V136 -93.65003646533025
L106_136 V106 V136 1.7190434882707796e-12
C106_136 V106 V136 6.349882664724084e-19

R106_137 V106 V137 520.8786586701859
L106_137 V106 V137 3.618259954606583e-12
C106_137 V106 V137 1.6821101615176542e-19

R106_138 V106 V138 77.59316120404247
L106_138 V106 V138 1.1102817519744908e-12
C106_138 V106 V138 4.392814761437908e-19

R106_139 V106 V139 65.75556997436045
L106_139 V106 V139 -1.2396374311402922e-12
C106_139 V106 V139 -8.657945718211864e-19

R106_140 V106 V140 46.92643114482155
L106_140 V106 V140 -8.442415778340732e-12
C106_140 V106 V140 -6.089592236430271e-19

R106_141 V106 V141 -196.43814671752716
L106_141 V106 V141 -4.590706059108968e-12
C106_141 V106 V141 -9.734355313378082e-20

R106_142 V106 V142 208.37084710190217
L106_142 V106 V142 2.5491461230605128e-12
C106_142 V106 V142 1.4784150120083307e-19

R106_143 V106 V143 -171.1596442386586
L106_143 V106 V143 3.628635130591926e-12
C106_143 V106 V143 7.693168765713714e-20

R106_144 V106 V144 -212.4456031358624
L106_144 V106 V144 -1.4174858971761824e-11
C106_144 V106 V144 2.3461397981598767e-21

R106_145 V106 V145 -635.9235505286631
L106_145 V106 V145 -6.8403485902177605e-12
C106_145 V106 V145 -1.0445145884323464e-19

R106_146 V106 V146 -36.035619372442135
L106_146 V106 V146 -8.332132332573636e-13
C106_146 V106 V146 -2.479954263578272e-19

R106_147 V106 V147 -122.47562525746825
L106_147 V106 V147 5.13599140854876e-12
C106_147 V106 V147 6.944625172693109e-19

R106_148 V106 V148 -83.73003353526518
L106_148 V106 V148 3.3552538529640107e-12
C106_148 V106 V148 4.170937144675028e-19

R106_149 V106 V149 -894.5758661218226
L106_149 V106 V149 3.827574761867089e-11
C106_149 V106 V149 1.2506758509571968e-19

R106_150 V106 V150 473.5087260171624
L106_150 V106 V150 1.7072216573445799e-12
C106_150 V106 V150 -1.5882103228532316e-19

R106_151 V106 V151 383.79897223966987
L106_151 V106 V151 -3.1815628248719486e-12
C106_151 V106 V151 -2.602579346751077e-19

R106_152 V106 V152 147.20991603245383
L106_152 V106 V152 -2.217358222245006e-12
C106_152 V106 V152 -1.3163731951545537e-19

R106_153 V106 V153 141.46586280078873
L106_153 V106 V153 7.01850568762546e-12
C106_153 V106 V153 1.3911793628365078e-19

R106_154 V106 V154 37.56946572476837
L106_154 V106 V154 3.4017981873707915e-12
C106_154 V106 V154 3.580028765033581e-19

R106_155 V106 V155 85.3570904279378
L106_155 V106 V155 -1.6076698106547742e-12
C106_155 V106 V155 -3.032987277124278e-19

R106_156 V106 V156 248.6062446566287
L106_156 V106 V156 2.154589332494063e-12
C106_156 V106 V156 -2.026701946843775e-19

R106_157 V106 V157 131.83526416896504
L106_157 V106 V157 3.88345234536196e-12
C106_157 V106 V157 -7.528608967189688e-20

R106_158 V106 V158 -53.438846359962405
L106_158 V106 V158 -3.0865340972325773e-12
C106_158 V106 V158 -2.286431259847179e-19

R106_159 V106 V159 -106.06921441505094
L106_159 V106 V159 1.0806632624432245e-12
C106_159 V106 V159 4.298484844627916e-19

R106_160 V106 V160 -219.84480437764094
L106_160 V106 V160 3.240439943370847e-12
C106_160 V106 V160 2.5652138224379953e-19

R106_161 V106 V161 -403.5188482194045
L106_161 V106 V161 -1.587217583505406e-12
C106_161 V106 V161 -2.530602883452661e-19

R106_162 V106 V162 -47.64608498131778
L106_162 V106 V162 -1.4904081979657358e-12
C106_162 V106 V162 -1.08115101634785e-19

R106_163 V106 V163 -2420.679441113313
L106_163 V106 V163 -1.7805687232538678e-12
C106_163 V106 V163 -3.0837575186958583e-19

R106_164 V106 V164 -434.5479073022223
L106_164 V106 V164 -2.449570065259533e-12
C106_164 V106 V164 -2.5992463562465073e-19

R106_165 V106 V165 -78.66555228681776
L106_165 V106 V165 2.9428527020982156e-12
C106_165 V106 V165 2.895143480775089e-19

R106_166 V106 V166 43.19208742758403
L106_166 V106 V166 1.1234871743208048e-12
C106_166 V106 V166 2.4067043581038815e-19

R106_167 V106 V167 -209.53470241382655
L106_167 V106 V167 -5.011641872199908e-12
C106_167 V106 V167 -1.161927688502213e-19

R106_168 V106 V168 -358.56757790313117
L106_168 V106 V168 -1.7280597126327472e-12
C106_168 V106 V168 -1.708141992378562e-19

R106_169 V106 V169 1139.2729786231164
L106_169 V106 V169 2.2380742967121073e-12
C106_169 V106 V169 2.543399546334552e-19

R106_170 V106 V170 245.18007810046586
L106_170 V106 V170 -2.535557400511845e-12
C106_170 V106 V170 -3.54283893487081e-20

R106_171 V106 V171 530.4019519486743
L106_171 V106 V171 2.1657459214990205e-12
C106_171 V106 V171 3.408036888196441e-19

R106_172 V106 V172 459.3938333503132
L106_172 V106 V172 1.0705431323145277e-12
C106_172 V106 V172 2.7804199329494557e-19

R106_173 V106 V173 118.20021608049503
L106_173 V106 V173 -1.9916750952059514e-12
C106_173 V106 V173 -1.9922544708085713e-19

R106_174 V106 V174 -42.72534263013787
L106_174 V106 V174 -3.371289408707239e-12
C106_174 V106 V174 1.0208373478365332e-20

R106_175 V106 V175 564.4061434777323
L106_175 V106 V175 -2.3491494651495096e-12
C106_175 V106 V175 -3.1374879780432557e-19

R106_176 V106 V176 213.32748860244618
L106_176 V106 V176 -2.3431407742513794e-12
C106_176 V106 V176 -2.466578122037351e-19

R106_177 V106 V177 -214.01715605006922
L106_177 V106 V177 2.323156742019437e-12
C106_177 V106 V177 1.8358077628782515e-19

R106_178 V106 V178 542.6597975147736
L106_178 V106 V178 1.9977507143959202e-12
C106_178 V106 V178 -6.626213679492054e-20

R106_179 V106 V179 680.6431965984362
L106_179 V106 V179 5.587033849515776e-12
C106_179 V106 V179 1.5354267447111072e-19

R106_180 V106 V180 -466.92592379763147
L106_180 V106 V180 2.1174677316187964e-10
C106_180 V106 V180 1.8987050189234974e-19

R106_181 V106 V181 -502.4429620287764
L106_181 V106 V181 -2.1458756982160647e-12
C106_181 V106 V181 -3.21504570573477e-19

R106_182 V106 V182 89.83546347560569
L106_182 V106 V182 -3.72380766761212e-11
C106_182 V106 V182 6.078983182237435e-20

R106_183 V106 V183 -549.8610234053716
L106_183 V106 V183 1.8123621542013087e-12
C106_183 V106 V183 -2.305291560796072e-20

R106_184 V106 V184 -1300.313041145935
L106_184 V106 V184 1.5680457664245903e-12
C106_184 V106 V184 -3.8135660388414593e-20

R106_185 V106 V185 169.1862260818407
L106_185 V106 V185 -5.825569375617324e-12
C106_185 V106 V185 4.471715777307809e-20

R106_186 V106 V186 -447.5311432315701
L106_186 V106 V186 4.188480411089975e-12
C106_186 V106 V186 7.025270930036708e-20

R106_187 V106 V187 -645.4393391856794
L106_187 V106 V187 -1.550755330354563e-12
C106_187 V106 V187 -2.6221835681060257e-19

R106_188 V106 V188 819.1871986954955
L106_188 V106 V188 -8.658892611477007e-13
C106_188 V106 V188 -1.809732864909121e-19

R106_189 V106 V189 -320.9419339967358
L106_189 V106 V189 1.1036074764252428e-12
C106_189 V106 V189 4.640333355078062e-19

R106_190 V106 V190 -78.59061764235909
L106_190 V106 V190 1.8792807077823768e-11
C106_190 V106 V190 -1.0904033334840675e-19

R106_191 V106 V191 -1485.3972917737117
L106_191 V106 V191 -1.2981565003330144e-11
C106_191 V106 V191 4.815663203615156e-19

R106_192 V106 V192 1189.1257022103794
L106_192 V106 V192 1.6444749864375895e-12
C106_192 V106 V192 5.478791560384285e-19

R106_193 V106 V193 -601.3897549259949
L106_193 V106 V193 -5.630383339918173e-12
C106_193 V106 V193 -1.236892575090804e-19

R106_194 V106 V194 210.44305454572896
L106_194 V106 V194 4.62638298428451e-12
C106_194 V106 V194 3.0503091798566e-19

R106_195 V106 V195 689.908892950076
L106_195 V106 V195 3.902038838819425e-12
C106_195 V106 V195 -5.094885747616398e-19

R106_196 V106 V196 -487.007754905252
L106_196 V106 V196 -7.349886340753718e-12
C106_196 V106 V196 -6.330339301134596e-19

R106_197 V106 V197 185.83475277539952
L106_197 V106 V197 -1.6255168049507031e-12
C106_197 V106 V197 -3.188626913397703e-19

R106_198 V106 V198 137.6544135426106
L106_198 V106 V198 -1.0049022907647122e-11
C106_198 V106 V198 8.998365829292543e-20

R106_199 V106 V199 -1023.8569546280406
L106_199 V106 V199 -2.8860414930701936e-12
C106_199 V106 V199 -2.103375393136855e-19

R106_200 V106 V200 397.3491253019281
L106_200 V106 V200 -2.7187052456608536e-12
C106_200 V106 V200 -1.9693402517076658e-19

R107_107 V107 0 -135.98698279977881
L107_107 V107 0 3.297377907711442e-13
C107_107 V107 0 2.2158833714296765e-18

R107_108 V107 V108 -427.35562884116155
L107_108 V107 V108 6.039987055718772e-12
C107_108 V107 V108 7.365512060247959e-20

R107_109 V107 V109 266.1380886797383
L107_109 V107 V109 -1.857032693032293e-12
C107_109 V107 V109 -4.273584926950171e-19

R107_110 V107 V110 -311.4491660421913
L107_110 V107 V110 -2.9302750979540717e-12
C107_110 V107 V110 -1.7343550324737861e-19

R107_111 V107 V111 127.1588604167105
L107_111 V107 V111 -6.916643824205374e-12
C107_111 V107 V111 -2.879050308997339e-19

R107_112 V107 V112 -2017.263727700115
L107_112 V107 V112 -5.525694590905836e-11
C107_112 V107 V112 7.86173839151172e-20

R107_113 V107 V113 -81.88797400525044
L107_113 V107 V113 -2.286239676052709e-12
C107_113 V107 V113 -3.6050325140850624e-20

R107_114 V107 V114 -1183.6032743183705
L107_114 V107 V114 -1.420993035636333e-12
C107_114 V107 V114 -4.088733560201911e-19

R107_115 V107 V115 103.4347365011359
L107_115 V107 V115 5.899258821276688e-13
C107_115 V107 V115 9.374586808526205e-19

R107_116 V107 V116 334.6099579769685
L107_116 V107 V116 9.284116488428995e-11
C107_116 V107 V116 -1.360909822756206e-19

R107_117 V107 V117 -592.8257349653502
L107_117 V107 V117 2.677099743745636e-12
C107_117 V107 V117 2.342076299451665e-19

R107_118 V107 V118 193.22600771831773
L107_118 V107 V118 1.3811413750658242e-12
C107_118 V107 V118 3.679647697881418e-19

R107_119 V107 V119 -66.90475492850058
L107_119 V107 V119 -2.6337280260000416e-12
C107_119 V107 V119 4.0052288707393463e-20

R107_120 V107 V120 -754.843551646336
L107_120 V107 V120 6.230071588782786e-12
C107_120 V107 V120 1.8341348404546367e-19

R107_121 V107 V121 85.7864972690278
L107_121 V107 V121 2.5130234893170005e-12
C107_121 V107 V121 -1.240095490715709e-20

R107_122 V107 V122 -772.3903937496237
L107_122 V107 V122 -1.405733701699785e-11
C107_122 V107 V122 -4.452909509972282e-20

R107_123 V107 V123 127.04335092182825
L107_123 V107 V123 -1.0070479676409516e-12
C107_123 V107 V123 -8.234366594985137e-19

R107_124 V107 V124 -1409.6918809679805
L107_124 V107 V124 -5.0522663497586355e-12
C107_124 V107 V124 -5.643798564370161e-20

R107_125 V107 V125 596.4517299141575
L107_125 V107 V125 -4.919781387387251e-12
C107_125 V107 V125 -8.365408982033231e-20

R107_126 V107 V126 -181.55791089660354
L107_126 V107 V126 -1.4737386905088907e-12
C107_126 V107 V126 -2.4548732139883283e-19

R107_127 V107 V127 168.5820197186838
L107_127 V107 V127 3.2579044049649923e-12
C107_127 V107 V127 1.199775471640706e-19

R107_128 V107 V128 863.5327199609898
L107_128 V107 V128 -8.82303077289304e-12
C107_128 V107 V128 -1.9075549941585224e-19

R107_129 V107 V129 -84.00737911189393
L107_129 V107 V129 -1.2760047116910369e-12
C107_129 V107 V129 -4.056644456238726e-19

R107_130 V107 V130 309.14821029926907
L107_130 V107 V130 1.3839760006168344e-12
C107_130 V107 V130 3.168805037425028e-19

R107_131 V107 V131 -115.48544126059672
L107_131 V107 V131 3.19416378443138e-12
C107_131 V107 V131 4.2300711129693282e-19

R107_132 V107 V132 -648.1536198294616
L107_132 V107 V132 2.245188240844914e-12
C107_132 V107 V132 3.917469918549527e-19

R107_133 V107 V133 -1160.0387655939958
L107_133 V107 V133 1.7789570713067965e-12
C107_133 V107 V133 4.439682566644121e-19

R107_134 V107 V134 -733.0593516595834
L107_134 V107 V134 -1.9095197715467835e-12
C107_134 V107 V134 -3.4652608616193845e-19

R107_135 V107 V135 89.09103323000063
L107_135 V107 V135 -2.2743785265745567e-11
C107_135 V107 V135 -4.955496561470599e-19

R107_136 V107 V136 -1745.021067326436
L107_136 V107 V136 1.654656822320102e-11
C107_136 V107 V136 -2.1973375314334535e-20

R107_137 V107 V137 95.12402724192813
L107_137 V107 V137 1.3358017574579313e-12
C107_137 V107 V137 2.988034182839608e-19

R107_138 V107 V138 1580.9503095096638
L107_138 V107 V138 -2.1601317633740988e-11
C107_138 V107 V138 9.202547047208096e-20

R107_139 V107 V139 -93.9063697043272
L107_139 V107 V139 5.080218061020207e-12
C107_139 V107 V139 6.072728957163796e-19

R107_140 V107 V140 -3541.3627834900235
L107_140 V107 V140 -3.693567852431653e-12
C107_140 V107 V140 -3.305859547462376e-20

R107_141 V107 V141 252.9464950050874
L107_141 V107 V141 -9.60218662172099e-13
C107_141 V107 V141 -7.93576050683124e-19

R107_142 V107 V142 450.75506745179695
L107_142 V107 V142 1.7861968994368043e-12
C107_142 V107 V142 1.3877416850986012e-19

R107_143 V107 V143 -127.42339734484815
L107_143 V107 V143 -1.0403506289686612e-12
C107_143 V107 V143 -2.9250115064957406e-19

R107_144 V107 V144 3096.734567791178
L107_144 V107 V144 -1.1049091564040535e-11
C107_144 V107 V144 -8.346545251068723e-20

R107_145 V107 V145 -75.23630693858037
L107_145 V107 V145 -1.2274682206589648e-12
C107_145 V107 V145 -2.4955419366761243e-19

R107_146 V107 V146 -134.18398586600279
L107_146 V107 V146 -1.7493999921631596e-12
C107_146 V107 V146 4.45793708007255e-21

R107_147 V107 V147 83.78469417131132
L107_147 V107 V147 1.5596058992832804e-12
C107_147 V107 V147 -3.38250207154564e-19

R107_148 V107 V148 -182.78026354616551
L107_148 V107 V148 -3.352865900348245e-12
C107_148 V107 V148 -2.4483137979935354e-20

R107_149 V107 V149 -467.86156175112643
L107_149 V107 V149 4.722808910955771e-13
C107_149 V107 V149 1.1116271422543108e-18

R107_150 V107 V150 251.44171027595124
L107_150 V107 V150 -1.568450150244004e-11
C107_150 V107 V150 -6.05135463573735e-19

R107_151 V107 V151 62.178989515938476
L107_151 V107 V151 1.584049729232468e-12
C107_151 V107 V151 1.8920636202593575e-19

R107_152 V107 V152 685.4714671511332
L107_152 V107 V152 -4.783241396824155e-11
C107_152 V107 V152 -5.135764094329161e-20

R107_153 V107 V153 139.28541742513661
L107_153 V107 V153 3.93291012625101e-12
C107_153 V107 V153 4.673988137557247e-20

R107_154 V107 V154 125.20494735435682
L107_154 V107 V154 3.45716193680028e-12
C107_154 V107 V154 3.9602360554602455e-19

R107_155 V107 V155 -64.30504135324495
L107_155 V107 V155 3.0643886613368545e-12
C107_155 V107 V155 5.132215964568646e-19

R107_156 V107 V156 224.37440901713697
L107_156 V107 V156 2.9259922849289387e-12
C107_156 V107 V156 1.2008108298293683e-19

R107_157 V107 V157 79.0189403695427
L107_157 V107 V157 -5.967976730344692e-13
C107_157 V107 V157 -9.314558243672515e-19

R107_158 V107 V158 -626.935365483748
L107_158 V107 V158 2.4347431674427293e-12
C107_158 V107 V158 7.054171944977481e-20

R107_159 V107 V159 -78.68183294548635
L107_159 V107 V159 -9.993077036159175e-13
C107_159 V107 V159 -2.1073714632136335e-19

R107_160 V107 V160 427.3654167329795
L107_160 V107 V160 3.177260970307059e-12
C107_160 V107 V160 1.4774618063156589e-19

R107_161 V107 V161 -127.30963616716569
L107_161 V107 V161 3.996011779885875e-11
C107_161 V107 V161 -4.116587340041751e-20

R107_162 V107 V162 -148.90684347573236
L107_162 V107 V162 3.792671131609607e-12
C107_162 V107 V162 1.4599638286090418e-19

R107_163 V107 V163 -544.6601701992358
L107_163 V107 V163 1.9676068662434638e-12
C107_163 V107 V163 4.334707081213285e-20

R107_164 V107 V164 -122.94522394951008
L107_164 V107 V164 -2.2604010193780768e-12
C107_164 V107 V164 -1.1520482652945448e-20

R107_165 V107 V165 -103.01988723193607
L107_165 V107 V165 1.6465685783054197e-12
C107_165 V107 V165 3.850942492159086e-19

R107_166 V107 V166 534.9190622192757
L107_166 V107 V166 -3.16329804060792e-12
C107_166 V107 V166 -1.9183920334068813e-19

R107_167 V107 V167 67.19700447546059
L107_167 V107 V167 -5.718983992398503e-12
C107_167 V107 V167 -1.8907472560470773e-19

R107_168 V107 V168 -490.1230620105997
L107_168 V107 V168 1.2779766408739746e-11
C107_168 V107 V168 -1.6076060909996742e-19

R107_169 V107 V169 169.1842949365023
L107_169 V107 V169 9.599843444881495e-12
C107_169 V107 V169 -6.969124796575257e-20

R107_170 V107 V170 778.3758106579337
L107_170 V107 V170 2.5223547258409122e-12
C107_170 V107 V170 2.72183563730836e-19

R107_171 V107 V171 759.3276458830837
L107_171 V107 V171 4.517843394972486e-12
C107_171 V107 V171 3.0219323286319288e-19

R107_172 V107 V172 239.32279922199004
L107_172 V107 V172 2.836446879281505e-12
C107_172 V107 V172 1.9039460403371109e-19

R107_173 V107 V173 204.766006906839
L107_173 V107 V173 -5.0674015943828856e-12
C107_173 V107 V173 -2.656547766193014e-20

R107_174 V107 V174 1216.5865419970073
L107_174 V107 V174 2.4635815539758455e-11
C107_174 V107 V174 -2.3681071594922647e-19

R107_175 V107 V175 -88.37731551617253
L107_175 V107 V175 1.2123694548375831e-12
C107_175 V107 V175 4.2514152228402044e-19

R107_176 V107 V176 -875.153655241512
L107_176 V107 V176 1.297915533599454e-10
C107_176 V107 V176 1.2688016041491266e-19

R107_177 V107 V177 -233.68722292439605
L107_177 V107 V177 -3.266471549543302e-12
C107_177 V107 V177 -9.77541277818618e-21

R107_178 V107 V178 533915.3759066514
L107_178 V107 V178 -1.7982069598976102e-12
C107_178 V107 V178 -1.1592826598571088e-19

R107_179 V107 V179 -152.58760851850548
L107_179 V107 V179 -1.3458946384569515e-12
C107_179 V107 V179 -6.292657548447686e-19

R107_180 V107 V180 -4989.860499004577
L107_180 V107 V180 -1.433956125730236e-12
C107_180 V107 V180 -3.201310981255708e-19

R107_181 V107 V181 1573.0499215262685
L107_181 V107 V181 3.91451233282868e-12
C107_181 V107 V181 -1.978568906043535e-19

R107_182 V107 V182 3402.320448274511
L107_182 V107 V182 9.558171091310259e-13
C107_182 V107 V182 2.8665507645131294e-19

R107_183 V107 V183 70.5677510708007
L107_183 V107 V183 -1.3553177206336843e-12
C107_183 V107 V183 -1.7991023151759993e-20

R107_184 V107 V184 1757.27541926219
L107_184 V107 V184 -4.043045327419115e-12
C107_184 V107 V184 -4.098538438729267e-20

R107_185 V107 V185 306.69990423207554
L107_185 V107 V185 1.7121052886219095e-11
C107_185 V107 V185 1.3928128012596273e-19

R107_186 V107 V186 -2132.688828984411
L107_186 V107 V186 -4.377234593531635e-12
C107_186 V107 V186 -2.173343310209261e-19

R107_187 V107 V187 -1237.5824691344178
L107_187 V107 V187 7.671054991701855e-13
C107_187 V107 V187 5.017294449113888e-19

R107_188 V107 V188 -828.4085905633525
L107_188 V107 V188 1.065587061601194e-12
C107_188 V107 V188 2.6867738086778173e-19

R107_189 V107 V189 -398.3720781653228
L107_189 V107 V189 7.3171004626555e-12
C107_189 V107 V189 2.0399663652052605e-19

R107_190 V107 V190 -8834.157013803908
L107_190 V107 V190 -3.651570362052586e-12
C107_190 V107 V190 -2.2129665289359813e-19

R107_191 V107 V191 -93.33312880083177
L107_191 V107 V191 2.009534211876813e-12
C107_191 V107 V191 -6.589749033116893e-20

R107_192 V107 V192 -1176.1905503111548
L107_192 V107 V192 3.929009539223431e-12
C107_192 V107 V192 1.558296500136911e-19

R107_193 V107 V193 -687.3360141111999
L107_193 V107 V193 -1.380183352978776e-11
C107_193 V107 V193 -1.1658929656372766e-19

R107_194 V107 V194 731.1291528858524
L107_194 V107 V194 1.1468572061822477e-11
C107_194 V107 V194 -4.0497992540427627e-20

R107_195 V107 V195 123.56877333676545
L107_195 V107 V195 -9.133267473676977e-13
C107_195 V107 V195 -8.75944542585326e-20

R107_196 V107 V196 563.8737786105869
L107_196 V107 V196 -8.994961480845415e-13
C107_196 V107 V196 -5.074285934752278e-19

R107_197 V107 V197 300.63067666913884
L107_197 V107 V197 -2.108083331974636e-12
C107_197 V107 V197 -2.5414801778470504e-19

R107_198 V107 V198 1020.0943861272632
L107_198 V107 V198 4.82586380049398e-12
C107_198 V107 V198 6.509215934590105e-20

R107_199 V107 V199 191.8548948610176
L107_199 V107 V199 -4.277692290848817e-12
C107_199 V107 V199 -9.13658587591176e-20

R107_200 V107 V200 481.48006544478307
L107_200 V107 V200 -1.682021081571895e-11
C107_200 V107 V200 2.173905866085371e-20

R108_108 V108 0 -41.268002758891754
L108_108 V108 0 6.541279433051434e-13
C108_108 V108 0 6.854092405232883e-19

R108_109 V108 V109 413.0820791559943
L108_109 V108 V109 2.572089518280536e-11
C108_109 V108 V109 -3.1807048416503625e-20

R108_110 V108 V110 -229.42930532308606
L108_110 V108 V110 5.037308808271264e-12
C108_110 V108 V110 1.6900826806640896e-19

R108_111 V108 V111 -772.2081373672107
L108_111 V108 V111 1.3743446855484133e-11
C108_111 V108 V111 7.904551392440462e-20

R108_112 V108 V112 92.34847524231357
L108_112 V108 V112 1.4885313962598233e-11
C108_112 V108 V112 -2.3222035515424403e-19

R108_113 V108 V113 -79.39566825165345
L108_113 V108 V113 -3.1401180619128344e-11
C108_113 V108 V113 1.3211044863538888e-19

R108_114 V108 V114 -2885.104236736687
L108_114 V108 V114 -2.006940221855256e-11
C108_114 V108 V114 -1.3202170208869284e-19

R108_115 V108 V115 782.8278185312323
L108_115 V108 V115 -4.145307445452803e-12
C108_115 V108 V115 -1.1151561404861872e-19

R108_116 V108 V116 75.2149199016201
L108_116 V108 V116 1.2306452132270248e-12
C108_116 V108 V116 5.551752173280305e-19

R108_117 V108 V117 -1385.5299710289476
L108_117 V108 V117 -2.433639202819017e-11
C108_117 V108 V117 2.811126653068932e-20

R108_118 V108 V118 159.41444623718712
L108_118 V108 V118 -7.88762619358339e-12
C108_118 V108 V118 -8.796002981693689e-20

R108_119 V108 V119 549.4285987787371
L108_119 V108 V119 8.726163058038396e-11
C108_119 V108 V119 -9.743295848797133e-21

R108_120 V108 V120 -48.755730018137285
L108_120 V108 V120 -1.6620934392323743e-12
C108_120 V108 V120 -3.607035736152102e-20

R108_121 V108 V121 105.83427043453196
L108_121 V108 V121 -9.983648227645135e-12
C108_121 V108 V121 -1.469557999185073e-19

R108_122 V108 V122 -278.49154010906415
L108_122 V108 V122 1.1296208826020312e-11
C108_122 V108 V122 1.0420225161121021e-19

R108_123 V108 V123 -327.553944882292
L108_123 V108 V123 2.947184014901387e-12
C108_123 V108 V123 1.9302980736391311e-19

R108_124 V108 V124 107.55072872209747
L108_124 V108 V124 2.8107333305298914e-12
C108_124 V108 V124 -3.662333327047938e-19

R108_125 V108 V125 2586.8192655394564
L108_125 V108 V125 -1.019708135770352e-11
C108_125 V108 V125 -5.472613300651454e-20

R108_126 V108 V126 -166.2738860539482
L108_126 V108 V126 5.643699683061413e-12
C108_126 V108 V126 6.025340217645099e-20

R108_127 V108 V127 -237.30016716494367
L108_127 V108 V127 -1.5556553716149522e-11
C108_127 V108 V127 -5.657981392758761e-20

R108_128 V108 V128 128.5339922009864
L108_128 V108 V128 -4.250406383778826e-12
C108_128 V108 V128 -5.0644983630502916e-20

R108_129 V108 V129 -97.86995615083808
L108_129 V108 V129 -1.7339051344830734e-11
C108_129 V108 V129 5.40218474287238e-20

R108_130 V108 V130 224.91548228536448
L108_130 V108 V130 1.7078802127341214e-10
C108_130 V108 V130 -5.919729439407209e-21

R108_131 V108 V131 164.25380605332907
L108_131 V108 V131 -5.4921675900448105e-12
C108_131 V108 V131 -1.0040110728529422e-19

R108_132 V108 V132 -92.15534681016669
L108_132 V108 V132 1.6519276950175523e-11
C108_132 V108 V132 3.3262926305701986e-19

R108_133 V108 V133 -708.9988121051085
L108_133 V108 V133 2.3341182299033085e-11
C108_133 V108 V133 1.2654657300273778e-19

R108_134 V108 V134 -520.4912797880859
L108_134 V108 V134 -2.0823321768663045e-11
C108_134 V108 V134 -1.1750102100696814e-20

R108_135 V108 V135 -390.5454855262488
L108_135 V108 V135 3.693194844265068e-12
C108_135 V108 V135 2.248493820293419e-19

R108_136 V108 V136 100.44311728174678
L108_136 V108 V136 1.770268484158524e-12
C108_136 V108 V136 -1.684738052286653e-19

R108_137 V108 V137 95.08634536603267
L108_137 V108 V137 2.619535419177654e-12
C108_137 V108 V137 1.5041772137588175e-20

R108_138 V108 V138 2015.445495149338
L108_138 V108 V138 4.623932437285529e-12
C108_138 V108 V138 6.123037598770607e-20

R108_139 V108 V139 -1408.6399176412924
L108_139 V108 V139 -3.659073285179969e-12
C108_139 V108 V139 -2.0823226872620353e-19

R108_140 V108 V140 -139.5350273436151
L108_140 V108 V140 -1.3279148547886636e-12
C108_140 V108 V140 1.0916551790528848e-19

R108_141 V108 V141 345.7923768552257
L108_141 V108 V141 -1.7468768346497863e-11
C108_141 V108 V141 -1.9904912523072844e-19

R108_142 V108 V142 1166.9999896897782
L108_142 V108 V142 -4.823538959717364e-11
C108_142 V108 V142 -1.2839885314441845e-20

R108_143 V108 V143 709.4223577597978
L108_143 V108 V143 3.871342393868059e-12
C108_143 V108 V143 2.730071623577021e-20

R108_144 V108 V144 -72.20298643041578
L108_144 V108 V144 -4.572006415445327e-12
C108_144 V108 V144 -7.351312203166919e-21

R108_145 V108 V145 -73.20888409762202
L108_145 V108 V145 -1.8216518495984114e-12
C108_145 V108 V145 1.334489786334893e-20

R108_146 V108 V146 -120.14925605848752
L108_146 V108 V146 -3.849171852755466e-12
C108_146 V108 V146 6.783546399614256e-21

R108_147 V108 V147 -230.43688923780047
L108_147 V108 V147 -3.785840672427545e-11
C108_147 V108 V147 1.2060038087229567e-19

R108_148 V108 V148 41.944071699281714
L108_148 V108 V148 1.3149897765145115e-12
C108_148 V108 V148 -1.872972968646915e-19

R108_149 V108 V149 -437.73932682934856
L108_149 V108 V149 -8.065769576686409e-12
C108_149 V108 V149 1.0569175523060715e-20

R108_150 V108 V150 152.39822687418447
L108_150 V108 V150 2.135418644737395e-11
C108_150 V108 V150 -1.576582045351715e-19

R108_151 V108 V151 1275.1124541713023
L108_151 V108 V151 -2.996533104614629e-12
C108_151 V108 V151 -1.1925862109540833e-19

R108_152 V108 V152 144.38618438656184
L108_152 V108 V152 2.3723906213084675e-12
C108_152 V108 V152 7.484023172724885e-20

R108_153 V108 V153 112.32598868174667
L108_153 V108 V153 2.4677780177302177e-12
C108_153 V108 V153 1.6323468436209394e-19

R108_154 V108 V154 141.49122165324962
L108_154 V108 V154 4.15442063965113e-12
C108_154 V108 V154 8.544231040570811e-20

R108_155 V108 V155 203.18425162965784
L108_155 V108 V155 -1.662043382017926e-11
C108_155 V108 V155 -1.6177705513576938e-20

R108_156 V108 V156 -505.62436753756646
L108_156 V108 V156 -1.4448521454543104e-12
C108_156 V108 V156 7.564322378145844e-20

R108_157 V108 V157 74.46443564119012
L108_157 V108 V157 3.794694629543555e-12
C108_157 V108 V157 -1.3085654862296845e-19

R108_158 V108 V158 2451.8129141627214
L108_158 V108 V158 1.060790495122329e-11
C108_158 V108 V158 -4.9834338704175e-21

R108_159 V108 V159 169.60947898057844
L108_159 V108 V159 2.2325357458664267e-12
C108_159 V108 V159 8.940052300022495e-20

R108_160 V108 V160 -40.97143900145648
L108_160 V108 V160 -2.50897081086703e-12
C108_160 V108 V160 3.886005358159174e-20

R108_161 V108 V161 -144.0922964584266
L108_161 V108 V161 -2.7073101310813735e-12
C108_161 V108 V161 -1.0598769379764806e-19

R108_162 V108 V162 -137.26929084399072
L108_162 V108 V162 -3.074353659024671e-12
C108_162 V108 V162 -3.720272035484263e-21

R108_163 V108 V163 -145.91260220081253
L108_163 V108 V163 -3.5483067505612243e-12
C108_163 V108 V163 -4.981948922261316e-20

R108_164 V108 V164 142.35244752815177
L108_164 V108 V164 1.1900234940343411e-12
C108_164 V108 V164 2.987335828069492e-20

R108_165 V108 V165 -131.41792915806192
L108_165 V108 V165 -2.182683641229116e-12
C108_165 V108 V165 -3.958809359549971e-20

R108_166 V108 V166 291.2169971018966
L108_166 V108 V166 -4.053826636899622e-12
C108_166 V108 V166 -1.1972588914244202e-19

R108_167 V108 V167 566.9501451781039
L108_167 V108 V167 -9.687717706644245e-11
C108_167 V108 V167 -4.421595981550363e-20

R108_168 V108 V168 131.69744594243025
L108_168 V108 V168 -2.1348370255484087e-12
C108_168 V108 V168 -2.076145071909156e-19

R108_169 V108 V169 176.21630454994227
L108_169 V108 V169 2.1608395770954432e-12
C108_169 V108 V169 1.0973810938859595e-19

R108_170 V108 V170 309.182455816534
L108_170 V108 V170 3.662732180935392e-12
C108_170 V108 V170 2.926714400497888e-20

R108_171 V108 V171 344.5507794197308
L108_171 V108 V171 -9.974393621883405e-10
C108_171 V108 V171 -4.851471091624894e-21

R108_172 V108 V172 226.33328075532384
L108_172 V108 V172 -4.454826155469665e-12
C108_172 V108 V172 1.403242484369702e-19

R108_173 V108 V173 176.1873237305217
L108_173 V108 V173 1.4023736786495125e-11
C108_173 V108 V173 2.4632246125543095e-20

R108_174 V108 V174 -339.7499302543513
L108_174 V108 V174 7.484948839042004e-12
C108_174 V108 V174 4.2334235302802146e-20

R108_175 V108 V175 2492.279726150975
L108_175 V108 V175 -1.1833367412328403e-11
C108_175 V108 V175 5.096795459557564e-21

R108_176 V108 V176 -105.3842641302543
L108_176 V108 V176 1.8916288538418842e-12
C108_176 V108 V176 2.257027089388602e-19

R108_177 V108 V177 -344.06267135383797
L108_177 V108 V177 -5.704503627402835e-12
C108_177 V108 V177 -8.674259904936272e-20

R108_178 V108 V178 1874.5229377141702
L108_178 V108 V178 -9.588784760534254e-12
C108_178 V108 V178 4.6596899355339474e-20

R108_179 V108 V179 572.4467175064026
L108_179 V108 V179 8.045403159053626e-12
C108_179 V108 V179 6.354264955758205e-20

R108_180 V108 V180 -69.96787236702782
L108_180 V108 V180 -4.9771426779610744e-11
C108_180 V108 V180 -1.9039678125519673e-19

R108_181 V108 V181 -1620.5312595640298
L108_181 V108 V181 -1.731204534421423e-11
C108_181 V108 V181 -1.3206973656100834e-19

R108_182 V108 V182 540.3114813009502
L108_182 V108 V182 -9.436926164403238e-12
C108_182 V108 V182 -5.2075466125061445e-20

R108_183 V108 V183 -245.35515142664275
L108_183 V108 V183 5.426957792313836e-12
C108_183 V108 V183 -4.20926793945853e-20

R108_184 V108 V184 61.501653639060635
L108_184 V108 V184 5.869744876440146e-11
C108_184 V108 V184 1.1121225896272397e-19

R108_185 V108 V185 221.24887814311342
L108_185 V108 V185 -1.0665906285199034e-11
C108_185 V108 V185 1.1494493147582993e-19

R108_186 V108 V186 -978.8646542589374
L108_186 V108 V186 -4.652146231354953e-12
C108_186 V108 V186 -6.033037597412434e-20

R108_187 V108 V187 -374.16651973100466
L108_187 V108 V187 -2.6340005220010064e-12
C108_187 V108 V187 -6.119825116102142e-22

R108_188 V108 V188 380.6501865201258
L108_188 V108 V188 -5.074688663707589e-12
C108_188 V108 V188 -9.248082054370896e-20

R108_189 V108 V189 -616.8175694352282
L108_189 V108 V189 2.8821422169811845e-12
C108_189 V108 V189 8.296297007044766e-20

R108_190 V108 V190 1772.3412212971853
L108_190 V108 V190 1.3230645375895671e-11
C108_190 V108 V190 -2.151567133671389e-20

R108_191 V108 V191 203.95881968926167
L108_191 V108 V191 -8.199545248504854e-12
C108_191 V108 V191 4.143038392281081e-20

R108_192 V108 V192 -70.54797349481386
L108_192 V108 V192 4.607169839544833e-12
C108_192 V108 V192 4.7486080500199183e-20

R108_193 V108 V193 -193.4216080290921
L108_193 V108 V193 7.322006524962366e-12
C108_193 V108 V193 1.6798910815638703e-20

R108_194 V108 V194 525.6959243252157
L108_194 V108 V194 2.4757086147770717e-12
C108_194 V108 V194 5.131709232862813e-20

R108_195 V108 V195 -1318.3873850811212
L108_195 V108 V195 2.8618320515441133e-12
C108_195 V108 V195 -1.5838199718005736e-19

R108_196 V108 V196 92.18683210909337
L108_196 V108 V196 8.831296078823908e-10
C108_196 V108 V196 9.820946277331778e-20

R108_197 V108 V197 416.6111979259637
L108_197 V108 V197 -4.117948767457166e-12
C108_197 V108 V197 -9.190923873052394e-20

R108_198 V108 V198 404.69282138613414
L108_198 V108 V198 -9.03932858842252e-12
C108_198 V108 V198 -4.56408474346234e-20

R108_199 V108 V199 272.122077269963
L108_199 V108 V199 -1.7912432229405193e-11
C108_199 V108 V199 -4.302099627705827e-20

R108_200 V108 V200 314.70836558308895
L108_200 V108 V200 -9.370914695435065e-12
C108_200 V108 V200 -2.9391084575360837e-20

R109_109 V109 0 -332.73784795663886
L109_109 V109 0 4.007755735876162e-13
C109_109 V109 0 2.2065645554887702e-18

R109_110 V109 V110 -17207.582130131246
L109_110 V109 V110 -3.5443739971671464e-12
C109_110 V109 V110 -2.8029493250607066e-19

R109_111 V109 V111 1752.2662477026238
L109_111 V109 V111 -1.0305003172535409e-11
C109_111 V109 V111 5.238002647453762e-20

R109_112 V109 V112 701.9153991715891
L109_112 V109 V112 -4.161301147057856e-12
C109_112 V109 V112 -1.8396669920770452e-19

R109_113 V109 V113 264.551030529223
L109_113 V109 V113 2.314284547322179e-12
C109_113 V109 V113 -6.22948453995961e-20

R109_114 V109 V114 -239.9813435642794
L109_114 V109 V114 -2.2582693726274484e-12
C109_114 V109 V114 -4.045271470870434e-19

R109_115 V109 V115 -223.20453466534335
L109_115 V109 V115 1.714784331210593e-12
C109_115 V109 V115 3.120926190412967e-19

R109_116 V109 V116 -246.39872114131467
L109_116 V109 V116 3.1402069575072104e-12
C109_116 V109 V116 1.0046935688958541e-19

R109_117 V109 V117 151.4828707921113
L109_117 V109 V117 2.0477003061001775e-12
C109_117 V109 V117 2.9976345222283817e-19

R109_118 V109 V118 260.0148299896315
L109_118 V109 V118 1.587160529008625e-12
C109_118 V109 V118 5.393926676398672e-19

R109_119 V109 V119 433.9641868106092
L109_119 V109 V119 -1.1911112818948562e-08
C109_119 V109 V119 1.2667885202210026e-19

R109_120 V109 V120 687.5724307310455
L109_120 V109 V120 8.942995520414374e-12
C109_120 V109 V120 3.9153312309756154e-19

R109_121 V109 V121 -122.26844406655357
L109_121 V109 V121 5.893183489576062e-12
C109_121 V109 V121 1.2963105901914136e-19

R109_122 V109 V122 -2097.2889768703017
L109_122 V109 V122 -6.3992400343692705e-12
C109_122 V109 V122 -8.789584568001405e-20

R109_123 V109 V123 695.4233020188481
L109_123 V109 V123 -2.296261346174148e-12
C109_123 V109 V123 -4.174604472161418e-19

R109_124 V109 V124 530.1761674269068
L109_124 V109 V124 -1.715074932414388e-12
C109_124 V109 V124 -6.749275486277674e-19

R109_125 V109 V125 -356.0877515752134
L109_125 V109 V125 -3.4244280518833863e-12
C109_125 V109 V125 -3.868866638475859e-20

R109_126 V109 V126 -732.9636689084152
L109_126 V109 V126 -1.5784580099373749e-12
C109_126 V109 V126 -2.833409733355154e-19

R109_127 V109 V127 -724.0455128535364
L109_127 V109 V127 -1.1769252522318475e-11
C109_127 V109 V127 -2.3206640348352705e-20

R109_128 V109 V128 -1216.8683570101662
L109_128 V109 V128 1.6767380400517732e-11
C109_128 V109 V128 8.225879106827196e-21

R109_129 V109 V129 111.2334210000833
L109_129 V109 V129 -1.5353653622355543e-12
C109_129 V109 V129 -5.712100909742846e-19

R109_130 V109 V130 535.174975037746
L109_130 V109 V130 1.606131607498315e-12
C109_130 V109 V130 3.1076375393849187e-19

R109_131 V109 V131 1098.4672261099086
L109_131 V109 V131 2.8354589198279114e-12
C109_131 V109 V131 3.203088430745252e-19

R109_132 V109 V132 4284.1247623008385
L109_132 V109 V132 1.967440646518785e-12
C109_132 V109 V132 5.703165683126229e-19

R109_133 V109 V133 -6231.068787815138
L109_133 V109 V133 2.4261143488046296e-12
C109_133 V109 V133 4.524356257778056e-19

R109_134 V109 V134 -425.6537882998021
L109_134 V109 V134 -2.7416996363708893e-12
C109_134 V109 V134 -1.0552634844460541e-19

R109_135 V109 V135 -359.500305305487
L109_135 V109 V135 -7.425044943728946e-12
C109_135 V109 V135 -2.4415952986681597e-19

R109_136 V109 V136 -648.0726107919494
L109_136 V109 V136 -3.946180431149071e-12
C109_136 V109 V136 -5.558411148551716e-19

R109_137 V109 V137 -119.94872742046047
L109_137 V109 V137 2.1854325793297232e-12
C109_137 V109 V137 1.761053726227598e-19

R109_138 V109 V138 38017.84235259057
L109_138 V109 V138 -2.2674173301243368e-11
C109_138 V109 V138 -9.210088981969233e-20

R109_139 V109 V139 2011.8426543463104
L109_139 V109 V139 6.20315424623458e-12
C109_139 V109 V139 3.552310889571168e-19

R109_140 V109 V140 -1194.8630213127306
L109_140 V109 V140 1.2149093502526201e-11
C109_140 V109 V140 5.142950629207628e-19

R109_141 V109 V141 -1523.1004340366835
L109_141 V109 V141 -1.2126682189685519e-12
C109_141 V109 V141 -5.0948499413766345e-19

R109_142 V109 V142 315.00244244755487
L109_142 V109 V142 4.404999145038323e-12
C109_142 V109 V142 5.618371387058398e-20

R109_143 V109 V143 169.18050000526705
L109_143 V109 V143 -3.615236876799479e-12
C109_143 V109 V143 -2.492050535921923e-19

R109_144 V109 V144 189.48326159635766
L109_144 V109 V144 -1.8356256558228587e-11
C109_144 V109 V144 -9.078114185297593e-20

R109_145 V109 V145 76.92499267622138
L109_145 V109 V145 -9.703110732233776e-12
C109_145 V109 V145 -1.4266060712381724e-19

R109_146 V109 V146 131.3736488163526
L109_146 V109 V146 5.6559609534301274e-11
C109_146 V109 V146 1.0034314734071918e-19

R109_147 V109 V147 -965.7465029300503
L109_147 V109 V147 -8.83671774219654e-12
C109_147 V109 V147 -2.961750052884339e-19

R109_148 V109 V148 1165.8563872895895
L109_148 V109 V148 -2.1738284842367076e-12
C109_148 V109 V148 -3.918998896683283e-19

R109_149 V109 V149 -410.8337181482786
L109_149 V109 V149 6.642040003604008e-13
C109_149 V109 V149 8.115453403291073e-19

R109_150 V109 V150 -82.19689940241337
L109_150 V109 V150 -8.510443050979192e-12
C109_150 V109 V150 -4.494800027370477e-19

R109_151 V109 V151 -128.39306552831565
L109_151 V109 V151 3.0983921156133036e-11
C109_151 V109 V151 2.336920925590286e-19

R109_152 V109 V152 -162.6857016918125
L109_152 V109 V152 3.950564616829009e-12
C109_152 V109 V152 9.810340869806054e-20

R109_153 V109 V153 -90.9293235526114
L109_153 V109 V153 -5.3390921365179355e-12
C109_153 V109 V153 -7.178490338477917e-20

R109_154 V109 V154 -130.16698180557825
L109_154 V109 V154 -1.9658993562584948e-11
C109_154 V109 V154 2.1662186622509248e-19

R109_155 V109 V155 652.6850651021301
L109_155 V109 V155 1.8039272387925975e-12
C109_155 V109 V155 3.4838809701849416e-19

R109_156 V109 V156 -692.2279568238428
L109_156 V109 V156 -2.1057704995609955e-11
C109_156 V109 V156 3.1687509300027356e-19

R109_157 V109 V157 -205.71721225404013
L109_157 V109 V157 -6.168492060753133e-13
C109_157 V109 V157 -8.98048338511822e-19

R109_158 V109 V158 89.63201900841318
L109_158 V109 V158 4.104818525938039e-12
C109_158 V109 V158 7.204987480660775e-20

R109_159 V109 V159 157.85813759869714
L109_159 V109 V159 -7.635967932926032e-12
C109_159 V109 V159 -2.1910955769512175e-19

R109_160 V109 V160 148.35211806707864
L109_160 V109 V160 4.2732789908214355e-12
C109_160 V109 V160 -9.64063465532641e-20

R109_161 V109 V161 125.60246569276433
L109_161 V109 V161 1.6381823084135086e-12
C109_161 V109 V161 2.6869887974682233e-19

R109_162 V109 V162 159.96886191564306
L109_162 V109 V162 2.1729608919067055e-12
C109_162 V109 V162 9.552432748734696e-20

R109_163 V109 V163 3303.051100140908
L109_163 V109 V163 -1.0296821470876305e-11
C109_163 V109 V163 -8.18255738387658e-20

R109_164 V109 V164 488.5663966443021
L109_164 V109 V164 -8.205273800461275e-12
C109_164 V109 V164 1.1946404309246526e-19

R109_165 V109 V165 211.5675628882964
L109_165 V109 V165 8.553163623482313e-12
C109_165 V109 V165 3.091982834146064e-19

R109_166 V109 V166 -63.74187307248995
L109_166 V109 V166 -2.739213059506154e-12
C109_166 V109 V166 -1.6971594297318506e-19

R109_167 V109 V167 -405.6539476246608
L109_167 V109 V167 -1.2999866211035902e-11
C109_167 V109 V167 6.237309454265166e-20

R109_168 V109 V168 -418.3525311826756
L109_168 V109 V168 3.271899679057077e-11
C109_168 V109 V168 -3.189919264779785e-20

R109_169 V109 V169 -169.4709046310901
L109_169 V109 V169 1.3410843639068578e-11
C109_169 V109 V169 -3.2215534389399436e-19

R109_170 V109 V170 151.93089525248922
L109_170 V109 V170 3.1344007797233323e-12
C109_170 V109 V170 2.449894439382954e-19

R109_171 V109 V171 958.3683528211424
L109_171 V109 V171 2.0548052251147732e-12
C109_171 V109 V171 2.3126008312988173e-19

R109_172 V109 V172 716.1351791433649
L109_172 V109 V172 2.5860344910950563e-11
C109_172 V109 V172 8.525155376745313e-20

R109_173 V109 V173 675.3972759753505
L109_173 V109 V173 9.829764961930234e-12
C109_173 V109 V173 -2.2391084668200274e-20

R109_174 V109 V174 126.39965313507828
L109_174 V109 V174 -9.101350948503258e-12
C109_174 V109 V174 -3.257112788479294e-19

R109_175 V109 V175 -1572.4595740926238
L109_175 V109 V175 7.099956698311852e-12
C109_175 V109 V175 1.1450282561372456e-19

R109_176 V109 V176 -704.2258545835077
L109_176 V109 V176 5.029971416787554e-12
C109_176 V109 V176 2.054852823604754e-19

R109_177 V109 V177 448.03448330522076
L109_177 V109 V177 -2.0987063289913003e-12
C109_177 V109 V177 4.888924663480418e-20

R109_178 V109 V178 -180.33888846839085
L109_178 V109 V178 -3.489001956504598e-12
C109_178 V109 V178 -9.876225427511621e-20

R109_179 V109 V179 736.9064998635189
L109_179 V109 V179 -2.3039578377403276e-12
C109_179 V109 V179 -4.482931085403239e-19

R109_180 V109 V180 1529.204676056674
L109_180 V109 V180 -2.5606628574998727e-12
C109_180 V109 V180 -4.19579374433072e-19

R109_181 V109 V181 1721.5949855531505
L109_181 V109 V181 2.932650683444649e-12
C109_181 V109 V181 2.390875661732981e-20

R109_182 V109 V182 -256.4227419795631
L109_182 V109 V182 1.741987325621453e-12
C109_182 V109 V182 2.565063120410627e-19

R109_183 V109 V183 3854.113960887596
L109_183 V109 V183 -2.3727356093654675e-12
C109_183 V109 V183 -7.886517595917184e-20

R109_184 V109 V184 583.2667849413361
L109_184 V109 V184 -3.3196724844549506e-12
C109_184 V109 V184 7.923349132690176e-20

R109_185 V109 V185 -318.7080428815103
L109_185 V109 V185 8.282890009959111e-12
C109_185 V109 V185 -6.994734460153414e-21

R109_186 V109 V186 484.01979976389725
L109_186 V109 V186 -2.9356858622337977e-12
C109_186 V109 V186 -2.4049993524455478e-21

R109_187 V109 V187 -1258.660870681371
L109_187 V109 V187 1.938124557541588e-12
C109_187 V109 V187 4.761563565524223e-19

R109_188 V109 V188 -312.94389744007395
L109_188 V109 V188 1.0757987546133991e-12
C109_188 V109 V188 3.640869856707863e-19

R109_189 V109 V189 -687.9033312258692
L109_189 V109 V189 -4.302188910807163e-12
C109_189 V109 V189 9.286169187658504e-20

R109_190 V109 V190 456.9048373968428
L109_190 V109 V190 -1.562008412772054e-10
C109_190 V109 V190 -2.4431248391520615e-19

R109_191 V109 V191 -849.215809420634
L109_191 V109 V191 1.3785579936930542e-12
C109_191 V109 V191 3.929162390543426e-20

R109_192 V109 V192 -116122.9169488673
L109_192 V109 V192 1.2008661953554011e-11
C109_192 V109 V192 -1.804751297326561e-19

R109_193 V109 V193 244.58365085075573
L109_193 V109 V193 2.799051942308199e-12
C109_193 V109 V193 -1.8522364236181186e-19

R109_194 V109 V194 -641.1500110779355
L109_194 V109 V194 1.616465907999114e-11
C109_194 V109 V194 -3.1192530232957175e-19

R109_195 V109 V195 1096.4483816527581
L109_195 V109 V195 -1.0045915835962844e-12
C109_195 V109 V195 -3.4578968801358153e-19

R109_196 V109 V196 947.0321032971696
L109_196 V109 V196 -1.5530158648481947e-12
C109_196 V109 V196 -2.9791768782825396e-20

R109_197 V109 V197 -20563.525402804127
L109_197 V109 V197 -2.756957744016057e-12
C109_197 V109 V197 -1.0329660571011604e-20

R109_198 V109 V198 -272.4890101972552
L109_198 V109 V198 -5.422684485487052e-12
C109_198 V109 V198 5.655175027802501e-21

R109_199 V109 V199 -1588.1161539277416
L109_199 V109 V199 -2.8857707419767974e-12
C109_199 V109 V199 -1.2441065690509374e-19

R109_200 V109 V200 1875.6190645063823
L109_200 V109 V200 -7.45976186095159e-12
C109_200 V109 V200 6.796374330247139e-20

R110_110 V110 0 -56.4240509739214
L110_110 V110 0 4.138823764008006e-13
C110_110 V110 0 1.3908338559046393e-18

R110_111 V110 V111 696.5626186247978
L110_111 V110 V111 3.836018247380607e-12
C110_111 V110 V111 9.793999802932903e-20

R110_112 V110 V112 445.6286531227443
L110_112 V110 V112 4.936786756351648e-12
C110_112 V110 V112 7.657824729564098e-20

R110_113 V110 V113 -123.55162038485422
L110_113 V110 V113 -7.48708684610761e-11
C110_113 V110 V113 9.16762779963414e-20

R110_114 V110 V114 -164.93072733359378
L110_114 V110 V114 1.2065277350619965e-11
C110_114 V110 V114 2.555006371297014e-19

R110_115 V110 V115 956.7271489081224
L110_115 V110 V115 2.4575163742446526e-12
C110_115 V110 V115 1.4697618332021909e-19

R110_116 V110 V116 496.10597221623004
L110_116 V110 V116 -7.414514453795906e-12
C110_116 V110 V116 -1.5658263701685386e-19

R110_117 V110 V117 628.7575403978517
L110_117 V110 V117 1.3922279712440166e-11
C110_117 V110 V117 2.865603660786022e-20

R110_118 V110 V118 56.035414214077626
L110_118 V110 V118 9.133496087120772e-13
C110_118 V110 V118 5.762545696304984e-19

R110_119 V110 V119 -1461.4614517510843
L110_119 V110 V119 -5.1379765815461954e-12
C110_119 V110 V119 3.374366681645878e-20

R110_120 V110 V120 -363.12861198639064
L110_120 V110 V120 -4.756382052282748e-11
C110_120 V110 V120 1.6190079425793495e-19

R110_121 V110 V121 176.42455271784374
L110_121 V110 V121 -1.8686299730998385e-11
C110_121 V110 V121 -5.16162447445305e-20

R110_122 V110 V122 -209.7320858923292
L110_122 V110 V122 -2.2585179914592277e-12
C110_122 V110 V122 -4.385917631339575e-19

R110_123 V110 V123 475.21652079914304
L110_123 V110 V123 -3.0469028000407115e-12
C110_123 V110 V123 -2.576915193753684e-19

R110_124 V110 V124 356.9484726729028
L110_124 V110 V124 -1.2180620906015131e-11
C110_124 V110 V124 -8.401702695071236e-20

R110_125 V110 V125 1446.625918722196
L110_125 V110 V125 9.773648824122397e-11
C110_125 V110 V125 9.550135934677575e-20

R110_126 V110 V126 -65.44953674778337
L110_126 V110 V126 -1.1070705989347511e-12
C110_126 V110 V126 -9.91827693808691e-20

R110_127 V110 V127 -205.9587706542177
L110_127 V110 V127 5.769965169026292e-12
C110_127 V110 V127 1.2581178544883207e-19

R110_128 V110 V128 -279.5622347909199
L110_128 V110 V128 3.011984951850861e-11
C110_128 V110 V128 -2.881702229960276e-20

R110_129 V110 V129 -137.0928248801603
L110_129 V110 V129 -1.4672252168985516e-11
C110_129 V110 V129 -2.075181068746094e-19

R110_130 V110 V130 108.81872177674728
L110_130 V110 V130 1.7119007059529652e-12
C110_130 V110 V130 1.6684638742178586e-19

R110_131 V110 V131 220.82607718354893
L110_131 V110 V131 2.843503664034835e-11
C110_131 V110 V131 4.98063789309543e-20

R110_132 V110 V132 206.02964106949094
L110_132 V110 V132 2.0887185872006908e-11
C110_132 V110 V132 1.0791817429946373e-19

R110_133 V110 V133 -1972.5301655807446
L110_133 V110 V133 -9.276880087434617e-12
C110_133 V110 V133 1.3021579289872574e-19

R110_134 V110 V134 142.5320639615033
L110_134 V110 V134 6.966585370773579e-12
C110_134 V110 V134 -4.415592550884566e-20

R110_135 V110 V135 192.411350038949
L110_135 V110 V135 -6.264743616109602e-12
C110_135 V110 V135 -2.9860393603494827e-19

R110_136 V110 V136 123.40956744492675
L110_136 V110 V136 2.6119195019669906e-11
C110_136 V110 V136 -1.2142304288039536e-19

R110_137 V110 V137 119.41840658487277
L110_137 V110 V137 3.863374889084002e-12
C110_137 V110 V137 1.3570343323223456e-19

R110_138 V110 V138 -106.0624496884073
L110_138 V110 V138 -2.2406764820437904e-12
C110_138 V110 V138 -4.040276253334907e-20

R110_139 V110 V139 -93.60116778006935
L110_139 V110 V139 2.616361623126995e-12
C110_139 V110 V139 5.096158157465438e-19

R110_140 V110 V140 -64.3537695849424
L110_140 V110 V140 -8.222555866966452e-12
C110_140 V110 V140 2.2410112219490707e-19

R110_141 V110 V141 260.6829538010961
L110_141 V110 V141 -4.1109138902978315e-12
C110_141 V110 V141 -3.407882904324666e-19

R110_142 V110 V142 -135.76619404226173
L110_142 V110 V142 -2.933593161062278e-12
C110_142 V110 V142 -1.227540030949172e-19

R110_143 V110 V143 411.48219788713595
L110_143 V110 V143 -2.2647495723922176e-12
C110_143 V110 V143 -2.1377675319891218e-19

R110_144 V110 V144 1497.9521715327232
L110_144 V110 V144 -5.809512566023143e-12
C110_144 V110 V144 -1.1763268956812733e-19

R110_145 V110 V145 -91.74638651115686
L110_145 V110 V145 -1.8161791126301694e-12
C110_145 V110 V145 -1.5720471755902683e-19

R110_146 V110 V146 107.29646461037252
L110_146 V110 V146 1.4522095595435691e-12
C110_146 V110 V146 1.779585506384019e-19

R110_147 V110 V147 405.47773763745204
L110_147 V110 V147 -8.99410574097362e-12
C110_147 V110 V147 -3.534303475577937e-19

R110_148 V110 V148 119.9706817439253
L110_148 V110 V148 -1.7165235777910384e-11
C110_148 V110 V148 -1.0815813801825559e-19

R110_149 V110 V149 -2240.7255111470836
L110_149 V110 V149 8.607694940513768e-13
C110_149 V110 V149 5.729128112322721e-19

R110_150 V110 V150 59.45436639823132
L110_150 V110 V150 5.038942535472608e-12
C110_150 V110 V150 -2.1544685144949046e-19

R110_151 V110 V151 1895.4758005448987
L110_151 V110 V151 6.360525784136386e-12
C110_151 V110 V151 2.276552235702083e-19

R110_152 V110 V152 -158.46536538381994
L110_152 V110 V152 1.4918423473195803e-11
C110_152 V110 V152 3.246237242335784e-20

R110_153 V110 V153 142.22910701754884
L110_153 V110 V153 7.067344238339092e-12
C110_153 V110 V153 5.0301200135815176e-20

R110_154 V110 V154 -108.43040554798287
L110_154 V110 V154 -3.8828593008642025e-12
C110_154 V110 V154 1.302683550127055e-19

R110_155 V110 V155 -140.4350455937287
L110_155 V110 V155 1.6063744777380427e-12
C110_155 V110 V155 2.638869336527395e-19

R110_156 V110 V156 252.1656367895628
L110_156 V110 V156 1.5113741724822315e-11
C110_156 V110 V156 1.1486517533845884e-19

R110_157 V110 V157 214.87803819940675
L110_157 V110 V157 -9.77019729878036e-13
C110_157 V110 V157 -4.969997000036566e-19

R110_158 V110 V158 -177.81705945303838
L110_158 V110 V158 -3.841875228385679e-12
C110_158 V110 V158 2.758387950561472e-20

R110_159 V110 V159 115.97711956697952
L110_159 V110 V159 -3.1806693324938896e-12
C110_159 V110 V159 -1.4873799670121703e-19

R110_160 V110 V160 288.79267328495746
L110_160 V110 V160 4.807335203789975e-12
C110_160 V110 V160 1.0126458389319673e-20

R110_161 V110 V161 -103.67990182618306
L110_161 V110 V161 4.181467286192534e-11
C110_161 V110 V161 -1.663160523659557e-20

R110_162 V110 V162 -1154.1179799131999
L110_162 V110 V162 1.2510628822353486e-12
C110_162 V110 V162 1.4204803790954081e-19

R110_163 V110 V163 -160.87035700753574
L110_163 V110 V163 -5.591749252777404e-12
C110_163 V110 V163 -1.4140959646911867e-20

R110_164 V110 V164 -168.93518757762726
L110_164 V110 V164 -3.662729299413499e-12
C110_164 V110 V164 1.4796969298334786e-20

R110_165 V110 V165 538.740230849548
L110_165 V110 V165 2.2653542769885227e-12
C110_165 V110 V165 2.4222341207939935e-19

R110_166 V110 V166 72.91344742246916
L110_166 V110 V166 9.677117386147871e-12
C110_166 V110 V166 -1.9883189913347308e-19

R110_167 V110 V167 -934.0196356653871
L110_167 V110 V167 8.859829502878575e-12
C110_167 V110 V167 3.1910572240117827e-20

R110_168 V110 V168 -143.43281337619277
L110_168 V110 V168 6.594775119688193e-12
C110_168 V110 V168 -4.982219477512715e-20

R110_169 V110 V169 88.10459641001464
L110_169 V110 V169 1.0207049615291824e-11
C110_169 V110 V169 -1.0915826636157065e-20

R110_170 V110 V170 -278.3158124515776
L110_170 V110 V170 -1.4755646944071287e-12
C110_170 V110 V170 1.9683847287389634e-19

R110_171 V110 V171 180.26121437183147
L110_171 V110 V171 2.813996906888726e-12
C110_171 V110 V171 9.515966674024328e-20

R110_172 V110 V172 130.91365050896079
L110_172 V110 V172 6.171948520619173e-12
C110_172 V110 V172 6.195331762249042e-20

R110_173 V110 V173 -130.51387927927985
L110_173 V110 V173 -3.7958371859685556e-12
C110_173 V110 V173 -1.0236612337315769e-19

R110_174 V110 V174 -91.57353655944914
L110_174 V110 V174 2.62080224512355e-12
C110_174 V110 V174 2.910458825797536e-20

R110_175 V110 V175 915.9574021383537
L110_175 V110 V175 3.4855247602540538e-12
C110_175 V110 V175 1.9493883168088816e-19

R110_176 V110 V176 771.014571472515
L110_176 V110 V176 2.4606165301754863e-11
C110_176 V110 V176 8.551415514181462e-20

R110_177 V110 V177 -415.7270159101664
L110_177 V110 V177 -2.723735284178926e-12
C110_177 V110 V177 -5.782478719436607e-20

R110_178 V110 V178 194.9859575162403
L110_178 V110 V178 6.862640897774961e-12
C110_178 V110 V178 -2.4348918363629364e-19

R110_179 V110 V179 -187.24132419890725
L110_179 V110 V179 -1.917656774723268e-12
C110_179 V110 V179 -3.281845666963647e-19

R110_180 V110 V180 -150.48724541066758
L110_180 V110 V180 -2.0471196632303194e-12
C110_180 V110 V180 -2.227626954273833e-19

R110_181 V110 V181 204.61466946074796
L110_181 V110 V181 2.329237206010775e-12
C110_181 V110 V181 8.26770456402759e-20

R110_182 V110 V182 113.84498438505786
L110_182 V110 V182 -8.90227236673935e-11
C110_182 V110 V182 1.6764772639584913e-19

R110_183 V110 V183 494.5790342532113
L110_183 V110 V183 -3.701972604118466e-12
C110_183 V110 V183 -1.382703009653123e-20

R110_184 V110 V184 475.94789716452647
L110_184 V110 V184 -2.434148422333292e-11
C110_184 V110 V184 -4.751931502724173e-21

R110_185 V110 V185 5124.837271135104
L110_185 V110 V185 6.004785238795934e-12
C110_185 V110 V185 1.8022980541271628e-20

R110_186 V110 V186 -583.9264053789816
L110_186 V110 V186 2.2884861083548212e-11
C110_186 V110 V186 4.323334323617648e-20

R110_187 V110 V187 -5773.766967906868
L110_187 V110 V187 1.3635822997204819e-12
C110_187 V110 V187 2.6265134287048767e-19

R110_188 V110 V188 -2291.5726066990305
L110_188 V110 V188 1.2762930879696261e-12
C110_188 V110 V188 1.6187387124910287e-19

R110_189 V110 V189 -895.0048347321728
L110_189 V110 V189 -4.968601240583714e-12
C110_189 V110 V189 -3.22184572382381e-20

R110_190 V110 V190 -507.5179241202982
L110_190 V110 V190 1.1632187738399733e-10
C110_190 V110 V190 -1.8667893721756682e-19

R110_191 V110 V191 -3738.6492720037922
L110_191 V110 V191 3.5604762830348004e-12
C110_191 V110 V191 -7.896731648626336e-20

R110_192 V110 V192 -631.5164996371074
L110_192 V110 V192 -2.3644802464098816e-11
C110_192 V110 V192 -2.791573929769216e-20

R110_193 V110 V193 -413.3830171249432
L110_193 V110 V193 -3.333709602644305e-11
C110_193 V110 V193 -3.391354148740516e-20

R110_194 V110 V194 412.8945000601722
L110_194 V110 V194 -3.5815793356253165e-12
C110_194 V110 V194 -2.618986880948847e-21

R110_195 V110 V195 735.4795751738335
L110_195 V110 V195 -2.479176004530746e-12
C110_195 V110 V195 2.3536249608015943e-20

R110_196 V110 V196 336.8571087593061
L110_196 V110 V196 -2.9048790847167904e-12
C110_196 V110 V196 -1.13510185131644e-19

R110_197 V110 V197 1906.7835895745932
L110_197 V110 V197 -5.0361938818521376e-12
C110_197 V110 V197 -6.806563851070591e-20

R110_198 V110 V198 200.29420875217158
L110_198 V110 V198 -2.7641106707659696e-11
C110_198 V110 V198 5.270824996181285e-21

R110_199 V110 V199 454.2326556397004
L110_199 V110 V199 -1.0889761998295162e-11
C110_199 V110 V199 -3.6547949910544246e-20

R110_200 V110 V200 -290.24852885245053
L110_200 V110 V200 -6.089048928441828e-10
C110_200 V110 V200 -1.6959971614761298e-20

R111_111 V111 0 665.9262443289572
L111_111 V111 0 2.0910982012266022e-12
C111_111 V111 0 -1.7251137388141556e-19

R111_112 V111 V112 -263.67362964658446
L111_112 V111 V112 2.8019598851118283e-08
C111_112 V111 V112 1.4076616489332576e-19

R111_113 V111 V113 336.31297105060514
L111_113 V111 V113 3.2848834882362263e-12
C111_113 V111 V113 -5.226663519872406e-20

R111_114 V111 V114 204.4495311600494
L111_114 V111 V114 9.310749684938176e-12
C111_114 V111 V114 -1.4182095039357717e-20

R111_115 V111 V115 491.2078058068298
L111_115 V111 V115 1.2244981223515187e-12
C111_115 V111 V115 4.563657799179112e-19

R111_116 V111 V116 247.71947866598816
L111_116 V111 V116 -1.8802677663942503e-11
C111_116 V111 V116 -1.3681568012932468e-19

R111_117 V111 V117 -443.0820062449161
L111_117 V111 V117 -1.3313385275154256e-10
C111_117 V111 V117 5.213371293417341e-20

R111_118 V111 V118 -355.6158831976623
L111_118 V111 V118 -2.6862216548414958e-12
C111_118 V111 V118 -1.479796239981134e-19

R111_119 V111 V119 78.61143711072499
L111_119 V111 V119 1.5126214752704793e-12
C111_119 V111 V119 -4.935671421438211e-20

R111_120 V111 V120 1197.9539964823457
L111_120 V111 V120 -1.7314931546494177e-11
C111_120 V111 V120 -1.3461088131603138e-19

R111_121 V111 V121 1454.9703622919483
L111_121 V111 V121 -7.130102044720821e-12
C111_121 V111 V121 -8.252856301470321e-21

R111_122 V111 V122 -433.9677158055619
L111_122 V111 V122 1.1492269064874376e-10
C111_122 V111 V122 4.216166866368789e-20

R111_123 V111 V123 -74.67781328871231
L111_123 V111 V123 -1.1122662774167133e-12
C111_123 V111 V123 -2.1235889918085883e-19

R111_124 V111 V124 -205.27919785913235
L111_124 V111 V124 4.1634383610095374e-12
C111_124 V111 V124 3.729698408785806e-19

R111_125 V111 V125 510.56325524684866
L111_125 V111 V125 -7.150938061793902e-12
C111_125 V111 V125 -6.544634184848824e-20

R111_126 V111 V126 1702.0549379837798
L111_126 V111 V126 4.136602757192745e-12
C111_126 V111 V126 8.217600393394863e-20

R111_127 V111 V127 -277.8149070401675
L111_127 V111 V127 -2.209538499850054e-12
C111_127 V111 V127 4.253538029379151e-20

R111_128 V111 V128 -2731.144027218014
L111_128 V111 V128 -4.744189185907795e-12
C111_128 V111 V128 -1.0967253079468412e-19

R111_129 V111 V129 -268.2191344756932
L111_129 V111 V129 -1.0285797098540412e-11
C111_129 V111 V129 5.233983808910796e-20

R111_130 V111 V130 439.43786088151603
L111_130 V111 V130 4.821292300249556e-10
C111_130 V111 V130 -3.4269482258605385e-20

R111_131 V111 V131 119.52323597401555
L111_131 V111 V131 1.194790369468567e-12
C111_131 V111 V131 9.03583593088733e-20

R111_132 V111 V132 180.88598970444846
L111_132 V111 V132 5.2225452783982776e-12
C111_132 V111 V132 -8.267594828548205e-20

R111_133 V111 V133 389.41825872178475
L111_133 V111 V133 3.425586450405437e-12
C111_133 V111 V133 -1.0353794915407305e-20

R111_134 V111 V134 322.1530145041471
L111_134 V111 V134 -1.1424895742993992e-11
C111_134 V111 V134 -1.5806209707054562e-19

R111_135 V111 V135 -119.78617334442666
L111_135 V111 V135 -3.250251632382739e-12
C111_135 V111 V135 -6.985942956967251e-20

R111_136 V111 V136 5160.424311827513
L111_136 V111 V136 3.6759872596615326e-12
C111_136 V111 V136 2.391353090541946e-19

R111_137 V111 V137 331.9024603801819
L111_137 V111 V137 4.644501904132382e-12
C111_137 V111 V137 4.473046973718023e-20

R111_138 V111 V138 -406.0374210072817
L111_138 V111 V138 1.3380396496679016e-11
C111_138 V111 V138 1.311619772233522e-19

R111_139 V111 V139 81.07779317249678
L111_139 V111 V139 4.6620127022472334e-12
C111_139 V111 V139 -2.49612603270215e-21

R111_140 V111 V140 5106.18024962119
L111_140 V111 V140 -3.3522112728382457e-12
C111_140 V111 V140 -2.729767526895857e-19

R111_141 V111 V141 -221.01649768281297
L111_141 V111 V141 -2.191620130640766e-12
C111_141 V111 V141 -4.893573258101311e-20

R111_142 V111 V142 -185.32327581845072
L111_142 V111 V142 -3.2421710951435235e-09
C111_142 V111 V142 5.8377164029893e-20

R111_143 V111 V143 -251.76614289546694
L111_143 V111 V143 -2.350706278544568e-11
C111_143 V111 V143 1.6306415630240255e-20

R111_144 V111 V144 -320.03444778289287
L111_144 V111 V144 -3.2447160842444766e-08
C111_144 V111 V144 3.95852362130825e-20

R111_145 V111 V145 -321.104052621797
L111_145 V111 V145 -3.775094520606e-12
C111_145 V111 V145 -3.469358649795437e-20

R111_146 V111 V146 6767.702004051978
L111_146 V111 V146 -8.355653660999338e-12
C111_146 V111 V146 -4.6982688786338905e-20

R111_147 V111 V147 -103.01680406661383
L111_147 V111 V147 -2.1418473160880173e-12
C111_147 V111 V147 4.3807187631371224e-20

R111_148 V111 V148 723.9961852474465
L111_148 V111 V148 2.175248407935816e-11
C111_148 V111 V148 1.3737877765040412e-19

R111_149 V111 V149 393.9319738719082
L111_149 V111 V149 2.160051440129889e-12
C111_149 V111 V149 7.243060517709073e-20

R111_150 V111 V150 149.00855512477116
L111_150 V111 V150 1.0551310530439505e-11
C111_150 V111 V150 -7.494826204869715e-20

R111_151 V111 V151 -465.9742773688695
L111_151 V111 V151 6.301849727524369e-12
C111_151 V111 V151 -4.806549147214322e-20

R111_152 V111 V152 -682.0993166282993
L111_152 V111 V152 -4.693385061677095e-12
C111_152 V111 V152 -5.414814150723994e-20

R111_153 V111 V153 135.71830527534829
L111_153 V111 V153 2.6604185773532582e-12
C111_153 V111 V153 1.3444212069561418e-20

R111_154 V111 V154 340.52751123981466
L111_154 V111 V154 7.679866724328817e-12
C111_154 V111 V154 6.842761914180601e-20

R111_155 V111 V155 45.8211821672471
L111_155 V111 V155 2.2473070347341414e-12
C111_155 V111 V155 6.194061451371662e-20

R111_156 V111 V156 260.04522587808964
L111_156 V111 V156 3.5268588409394153e-12
C111_156 V111 V156 -1.017511626781167e-19

R111_157 V111 V157 1298.0283696213253
L111_157 V111 V157 -3.330874662419381e-12
C111_157 V111 V157 1.0956054922442986e-20

R111_158 V111 V158 -134.91501712382356
L111_158 V111 V158 1.85043290261583e-11
C111_158 V111 V158 -1.6897563246659064e-20

R111_159 V111 V159 -112.2158402818318
L111_159 V111 V159 -2.3136165751693814e-12
C111_159 V111 V159 -1.2182649599642724e-20

R111_160 V111 V160 -894.8307080893712
L111_160 V111 V160 4.9835096825489345e-12
C111_160 V111 V160 8.89624875717839e-20

R111_161 V111 V161 -212.32986952526733
L111_161 V111 V161 -3.2853381279140583e-12
C111_161 V111 V161 -7.398517588043387e-20

R111_162 V111 V162 -211.44387486064124
L111_162 V111 V162 -9.975302080594082e-12
C111_162 V111 V162 2.262744713082971e-20

R111_163 V111 V163 -141.13010870110725
L111_163 V111 V163 3.200762371870308e-12
C111_163 V111 V163 9.017998675392054e-20

R111_164 V111 V164 -183.83144878976375
L111_164 V111 V164 -4.9180247479803e-12
C111_164 V111 V164 -2.2707921204015996e-20

R111_165 V111 V165 -631.5088647748739
L111_165 V111 V165 2.3810021304961504e-10
C111_165 V111 V165 3.745865545051253e-20

R111_166 V111 V166 133.53268468280342
L111_166 V111 V166 -2.0010165325705073e-11
C111_166 V111 V166 4.2346855798502475e-20

R111_167 V111 V167 146.19756808128153
L111_167 V111 V167 1.474717964156028e-11
C111_167 V111 V167 -1.7132568932116074e-19

R111_168 V111 V168 812.2175447999608
L111_168 V111 V168 -6.117582349505336e-12
C111_168 V111 V168 -5.527968031686205e-20

R111_169 V111 V169 275.38547183300744
L111_169 V111 V169 2.9662759290762445e-12
C111_169 V111 V169 5.884387835557219e-20

R111_170 V111 V170 1247.8910001901647
L111_170 V111 V170 7.392619630586208e-12
C111_170 V111 V170 -2.2519756081995253e-20

R111_171 V111 V171 -894.7567095478008
L111_171 V111 V171 -2.4612791844658705e-12
C111_171 V111 V171 1.1006512198822377e-19

R111_172 V111 V172 312.60364301113833
L111_172 V111 V172 3.628426933521392e-12
C111_172 V111 V172 4.99152938580881e-20

R111_173 V111 V173 -803.18130372248
L111_173 V111 V173 -5.1348659967776e-12
C111_173 V111 V173 -1.3576891609794783e-21

R111_174 V111 V174 -193.10311637081378
L111_174 V111 V174 5.294796280596227e-12
C111_174 V111 V174 -6.234934070930606e-21

R111_175 V111 V175 -297.18866474019615
L111_175 V111 V175 2.475933248520374e-12
C111_175 V111 V175 7.524034360341286e-20

R111_176 V111 V176 -831.9768591448322
L111_176 V111 V176 4.428489279338959e-11
C111_176 V111 V176 -6.711342707203644e-20

R111_177 V111 V177 -529.1661278807948
L111_177 V111 V177 -5.980733510445337e-11
C111_177 V111 V177 1.3075049644575704e-20

R111_178 V111 V178 -349.53128891210196
L111_178 V111 V178 -3.4016284659769013e-12
C111_178 V111 V178 2.6742561090699865e-20

R111_179 V111 V179 86.52896575214265
L111_179 V111 V179 2.3228218682592877e-12
C111_179 V111 V179 -8.297870428528785e-20

R111_180 V111 V180 -416.1423716009573
L111_180 V111 V180 -4.568094842405891e-12
C111_180 V111 V180 6.503503864384095e-20

R111_181 V111 V181 555.5771508911466
L111_181 V111 V181 -1.1446219868880949e-11
C111_181 V111 V181 -1.0121828043205624e-19

R111_182 V111 V182 136.83112040526433
L111_182 V111 V182 4.480508893095188e-12
C111_182 V111 V182 2.1240946514300397e-20

R111_183 V111 V183 -115.0645403360645
L111_183 V111 V183 -1.8206107018505184e-12
C111_183 V111 V183 4.334007211464225e-21

R111_184 V111 V184 524.0163861064561
L111_184 V111 V184 6.318587450982157e-12
C111_184 V111 V184 -2.0436047618417782e-20

R111_185 V111 V185 736.9714825788534
L111_185 V111 V185 -1.482162660772404e-11
C111_185 V111 V185 3.818038323219313e-20

R111_186 V111 V186 566.3610056677783
L111_186 V111 V186 6.6912178614779624e-12
C111_186 V111 V186 -6.789777599944607e-20

R111_187 V111 V187 -274.78287131308537
L111_187 V111 V187 -9.176332441757475e-12
C111_187 V111 V187 4.721315801795044e-20

R111_188 V111 V188 2616.307590967317
L111_188 V111 V188 -4.119952124360509e-12
C111_188 V111 V188 -7.971391532196495e-20

R111_189 V111 V189 -515.1441396828711
L111_189 V111 V189 2.6761519940410672e-12
C111_189 V111 V189 1.0585364887683051e-19

R111_190 V111 V190 -175.5198227393419
L111_190 V111 V190 -4.483169095833418e-12
C111_190 V111 V190 -1.335176281923387e-20

R111_191 V111 V191 164.34446866246893
L111_191 V111 V191 1.9163416600696764e-12
C111_191 V111 V191 -4.3283861965360585e-22

R111_192 V111 V192 -1018.1184530018353
L111_192 V111 V192 3.4120338025829366e-12
C111_192 V111 V192 1.8493934396458878e-19

R111_193 V111 V193 -2784.9000813987923
L111_193 V111 V193 -2.719320171857314e-11
C111_193 V111 V193 -7.767344453124796e-21

R111_194 V111 V194 306.1530010290942
L111_194 V111 V194 1.8369565441228324e-12
C111_194 V111 V194 1.3755340182044068e-19

R111_195 V111 V195 -276.4660889224094
L111_195 V111 V195 -1.5072481889446992e-12
C111_195 V111 V195 1.8029215967818943e-20

R111_196 V111 V196 -1154.7011492658662
L111_196 V111 V196 -6.471782621251424e-12
C111_196 V111 V196 -2.743892887975227e-19

R111_197 V111 V197 1488.0708303731449
L111_197 V111 V197 -3.747892859145864e-12
C111_197 V111 V197 -8.464039594848228e-20

R111_198 V111 V198 370.6053161406613
L111_198 V111 V198 2.9643753220362365e-10
C111_198 V111 V198 9.591815740522868e-21

R111_199 V111 V199 -771.6151241300338
L111_199 V111 V199 2.3466470036759676e-11
C111_199 V111 V199 4.1083317286348953e-20

R111_200 V111 V200 -2132.5071964957997
L111_200 V111 V200 -4.79289982534816e-12
C111_200 V111 V200 -8.965545008897026e-21

R112_112 V112 0 181.35131287170503
L112_112 V112 0 4.263925390174368e-13
C112_112 V112 0 1.4123158360244784e-18

R112_113 V112 V113 366.564659452715
L112_113 V112 V113 -6.523946498119702e-11
C112_113 V112 V113 -1.4277131874676123e-19

R112_114 V112 V114 288.52394204271025
L112_114 V112 V114 -2.3635755736074925e-12
C112_114 V112 V114 -2.7832129464592784e-19

R112_115 V112 V115 212.5437336733286
L112_115 V112 V115 -5.78657366260245e-12
C112_115 V112 V115 -2.3947490661789555e-19

R112_116 V112 V116 -418.61744553254283
L112_116 V112 V116 9.356912557915359e-13
C112_116 V112 V116 6.101084485778856e-19

R112_117 V112 V117 -359.7568841422046
L112_117 V112 V117 1.7124495810603934e-11
C112_117 V112 V117 1.0323394636324787e-19

R112_118 V112 V118 -386.0742406573114
L112_118 V112 V118 -3.1999473479739674e-11
C112_118 V112 V118 6.224271899440163e-20

R112_119 V112 V119 9737.584076091982
L112_119 V112 V119 7.2133441224993135e-12
C112_119 V112 V119 1.2765432419441927e-19

R112_120 V112 V120 64.63669008611448
L112_120 V112 V120 9.424935220476914e-13
C112_120 V112 V120 4.049202093941491e-19

R112_121 V112 V121 437.36795113194256
L112_121 V112 V121 5.883167382847463e-12
C112_121 V112 V121 7.125273456963807e-20

R112_122 V112 V122 -4579.429900762084
L112_122 V112 V122 5.4681956201857866e-12
C112_122 V112 V122 1.5049873744762792e-19

R112_123 V112 V123 -308.11932656710945
L112_123 V112 V123 3.2024999921577455e-12
C112_123 V112 V123 2.951007481985474e-19

R112_124 V112 V124 -81.87377222347689
L112_124 V112 V124 -4.353222536195973e-13
C112_124 V112 V124 -1.1240368925291034e-18

R112_125 V112 V125 309.6040012025473
L112_125 V112 V125 -1.9024098747648793e-11
C112_125 V112 V125 -3.9164648372566175e-20

R112_126 V112 V126 2019.7323181300906
L112_126 V112 V126 -6.007137756914284e-12
C112_126 V112 V126 -4.304532966257742e-20

R112_127 V112 V127 328.7614803892907
L112_127 V112 V127 -1.822888328829353e-12
C112_127 V112 V127 -3.9252652177397172e-19

R112_128 V112 V128 -165.1858789638803
L112_128 V112 V128 4.214260118500533e-12
C112_128 V112 V128 2.9132793281665215e-19

R112_129 V112 V129 -201.28337136213057
L112_129 V112 V129 -2.98090082980625e-12
C112_129 V112 V129 -9.990962686955065e-20

R112_130 V112 V130 949.2548721066305
L112_130 V112 V130 8.61688499910509e-12
C112_130 V112 V130 2.52718519348351e-20

R112_131 V112 V131 -1533.2371115291648
L112_131 V112 V131 4.888611240984064e-12
C112_131 V112 V131 1.5503009279420285e-19

R112_132 V112 V132 85.73772976243997
L112_132 V112 V132 8.468531561454178e-13
C112_132 V112 V132 3.0228164792240663e-19

R112_133 V112 V133 475.1748762286985
L112_133 V112 V133 2.4175519618744982e-12
C112_133 V112 V133 1.4317611663844641e-19

R112_134 V112 V134 256.4914375959409
L112_134 V112 V134 6.84467618579124e-12
C112_134 V112 V134 1.0409622243700335e-19

R112_135 V112 V135 1286.3273728244958
L112_135 V112 V135 1.565993517719936e-12
C112_135 V112 V135 4.363161607451448e-19

R112_136 V112 V136 -170.98670377290532
L112_136 V112 V136 -9.100850892721377e-13
C112_136 V112 V136 -6.450592003223172e-19

R112_137 V112 V137 301.3759902239737
L112_137 V112 V137 2.1512447080818672e-10
C112_137 V112 V137 -9.665931254487728e-20

R112_138 V112 V138 -346.40947486985414
L112_138 V112 V138 -3.698334646756919e-12
C112_138 V112 V138 -1.0810852091246622e-19

R112_139 V112 V139 1145.4879746106078
L112_139 V112 V139 -1.1349261759834177e-12
C112_139 V112 V139 -5.695556805759199e-19

R112_140 V112 V140 154.79982407716588
L112_140 V112 V140 1.2727471966108011e-12
C112_140 V112 V140 6.348485443118409e-19

R112_141 V112 V141 -353.6199544691208
L112_141 V112 V141 -2.268519494033466e-12
C112_141 V112 V141 -7.040275961357563e-20

R112_142 V112 V142 -209.60386922528116
L112_142 V112 V142 -1.541022078300006e-11
C112_142 V112 V142 3.943885085950887e-20

R112_143 V112 V143 -352.0906627274768
L112_143 V112 V143 -6.063569911062493e-11
C112_143 V112 V143 5.617260285902464e-20

R112_144 V112 V144 981.7769203827729
L112_144 V112 V144 -1.0001385011040361e-11
C112_144 V112 V144 -8.168630080917734e-20

R112_145 V112 V145 -371.95209267764733
L112_145 V112 V145 -1.644639939524359e-11
C112_145 V112 V145 6.888618815036948e-20

R112_146 V112 V146 519.0998413286408
L112_146 V112 V146 3.6375525119556907e-12
C112_146 V112 V146 2.5004173065804263e-20

R112_147 V112 V147 -1767.2738859936283
L112_147 V112 V147 1.9084150731679792e-11
C112_147 V112 V147 1.8094009021753437e-19

R112_148 V112 V148 -67.76008463640399
L112_148 V112 V148 -7.738500063508533e-13
C112_148 V112 V148 -3.482023086250731e-19

R112_149 V112 V149 1677.6028353500283
L112_149 V112 V149 1.6802795888441703e-12
C112_149 V112 V149 1.2258924732717102e-19

R112_150 V112 V150 192.46632048542128
L112_150 V112 V150 -6.259913987504423e-12
C112_150 V112 V150 -1.4998619713835273e-19

R112_151 V112 V151 2254.1373876325165
L112_151 V112 V151 6.861281387863345e-12
C112_151 V112 V151 -3.97655424112772e-20

R112_152 V112 V152 604.2079736067627
L112_152 V112 V152 9.989598913234499e-13
C112_152 V112 V152 1.0666246940801746e-19

R112_153 V112 V153 137.1940061393514
L112_153 V112 V153 2.4960425205631532e-12
C112_153 V112 V153 -6.219413964449355e-20

R112_154 V112 V154 375.8857392542829
L112_154 V112 V154 2.7924066483914305e-12
C112_154 V112 V154 3.550725313236259e-20

R112_155 V112 V155 318.50867142449056
L112_155 V112 V155 -4.134144444732593e-11
C112_155 V112 V155 -1.393685615186904e-19

R112_156 V112 V156 87.34795294913962
L112_156 V112 V156 9.888350678568838e-12
C112_156 V112 V156 3.2298382659286896e-19

R112_157 V112 V157 4340.608117429298
L112_157 V112 V157 -1.1281779498715043e-12
C112_157 V112 V157 -3.110153083914911e-19

R112_158 V112 V158 -126.11650722753383
L112_158 V112 V158 -1.1961884645228682e-11
C112_158 V112 V158 1.5773416950273343e-20

R112_159 V112 V159 -531.705442163408
L112_159 V112 V159 3.191793673537113e-12
C112_159 V112 V159 1.5717336651296358e-19

R112_160 V112 V160 2064.4105832713326
L112_160 V112 V160 -2.163048950000449e-12
C112_160 V112 V160 -2.1285631677661554e-19

R112_161 V112 V161 -228.529017416138
L112_161 V112 V161 5.735879389683436e-12
C112_161 V112 V161 1.5374157555430022e-19

R112_162 V112 V162 -320.0480904832518
L112_162 V112 V162 1.307029404035719e-11
C112_162 V112 V162 3.8253077299630176e-21

R112_163 V112 V163 -374.9669385516785
L112_163 V112 V163 -3.3473290320240097e-12
C112_163 V112 V163 -1.5032131800895375e-19

R112_164 V112 V164 -69.53316525130583
L112_164 V112 V164 -8.886070664601495e-12
C112_164 V112 V164 1.391830759168896e-19

R112_165 V112 V165 -448.6206436344439
L112_165 V112 V165 1.0013923944911999e-11
C112_165 V112 V165 6.653194822605681e-20

R112_166 V112 V166 173.5913551260501
L112_166 V112 V166 -7.58207728852357e-12
C112_166 V112 V166 -4.1956518501853045e-20

R112_167 V112 V167 -272.22003896252835
L112_167 V112 V167 -1.759887633636682e-10
C112_167 V112 V167 8.158338700176447e-20

R112_168 V112 V168 77.40931329130296
L112_168 V112 V168 1.3407981691134884e-12
C112_168 V112 V168 -4.16488807561242e-21

R112_169 V112 V169 236.66173316454496
L112_169 V112 V169 3.0888976492612356e-11
C112_169 V112 V169 -2.2684713156310614e-19

R112_170 V112 V170 1828.4396929593831
L112_170 V112 V170 3.879990663717225e-12
C112_170 V112 V170 2.5180905366332682e-20

R112_171 V112 V171 258.4764303148811
L112_171 V112 V171 1.6781372777595812e-12
C112_171 V112 V171 1.0495274445786325e-19

R112_172 V112 V172 -348.21433859985177
L112_172 V112 V172 -1.2118555081304066e-12
C112_172 V112 V172 -3.21947658267853e-20

R112_173 V112 V173 -507.6827221294923
L112_173 V112 V173 -7.816819731916768e-12
C112_173 V112 V173 5.2310715649656134e-20

R112_174 V112 V174 -331.7395384533275
L112_174 V112 V174 -3.4114198911608856e-11
C112_174 V112 V174 -1.1428193054307104e-19

R112_175 V112 V175 -6348.337104988347
L112_175 V112 V175 -2.2273264268877024e-12
C112_175 V112 V175 -2.0713145540079546e-19

R112_176 V112 V176 -208.15529320176955
L112_176 V112 V176 2.1522145448277046e-12
C112_176 V112 V176 3.265970722762375e-19

R112_177 V112 V177 -345.03220825354384
L112_177 V112 V177 -2.4041446156129594e-11
C112_177 V112 V177 5.602798386022251e-20

R112_178 V112 V178 -283.22885481702826
L112_178 V112 V178 -2.159896729817728e-12
C112_178 V112 V178 3.766404097558091e-21

R112_179 V112 V179 -341.86939028114966
L112_179 V112 V179 -2.2442276571359242e-12
C112_179 V112 V179 1.4572351742382207e-20

R112_180 V112 V180 83.28407775015867
L112_180 V112 V180 2.685835999212737e-12
C112_180 V112 V180 -3.3133714134144326e-19

R112_181 V112 V181 388.2347215372174
L112_181 V112 V181 8.422681728132664e-11
C112_181 V112 V181 1.866020480438614e-20

R112_182 V112 V182 166.85519036949862
L112_182 V112 V182 2.8652300483524868e-12
C112_182 V112 V182 4.4343588012398946e-20

R112_183 V112 V183 386.6636268882081
L112_183 V112 V183 5.991829323680516e-12
C112_183 V112 V183 -8.570432138066661e-20

R112_184 V112 V184 -138.49463737229445
L112_184 V112 V184 -1.1420099769321872e-12
C112_184 V112 V184 3.3318342147546653e-20

R112_185 V112 V185 1235.365152169251
L112_185 V112 V185 2.021959549478724e-11
C112_185 V112 V185 -5.141449774603287e-20

R112_186 V112 V186 629.1664804424422
L112_186 V112 V186 -7.238288140480826e-10
C112_186 V112 V186 3.275719176286307e-20

R112_187 V112 V187 980.4025536390753
L112_187 V112 V187 -1.01027400212668e-11
C112_187 V112 V187 -3.838494515482535e-20

R112_188 V112 V188 -278.56814484158207
L112_188 V112 V188 8.686756202170043e-13
C112_188 V112 V188 3.350609279921864e-19

R112_189 V112 V189 -471.8246966319073
L112_189 V112 V189 -1.683024102688148e-11
C112_189 V112 V189 -9.182757108416442e-21

R112_190 V112 V190 -199.25656919701166
L112_190 V112 V190 -3.4108284270077958e-12
C112_190 V112 V190 -6.479138699720075e-20

R112_191 V112 V191 -394.67114153128165
L112_191 V112 V191 1.8241573996332883e-12
C112_191 V112 V191 2.748243736469693e-19

R112_192 V112 V192 155.73628788123096
L112_192 V112 V192 -4.966096343810167e-12
C112_192 V112 V192 -3.428130974233835e-19

R112_193 V112 V193 748.4149192207933
L112_193 V112 V193 -4.4784510223307014e-11
C112_193 V112 V193 -8.565760202708282e-20

R112_194 V112 V194 411.76277687936096
L112_194 V112 V194 -2.615411160124742e-11
C112_194 V112 V194 -2.128280758304608e-19

R112_195 V112 V195 806.1277162644845
L112_195 V112 V195 -1.2492871031603778e-12
C112_195 V112 V195 -5.5282045755671215e-19

R112_196 V112 V196 -187.75501158028706
L112_196 V112 V196 4.6192641355145877e-11
C112_196 V112 V196 5.181513535410348e-19

R112_197 V112 V197 896.2910079578647
L112_197 V112 V197 -3.4034896968404654e-11
C112_197 V112 V197 9.662983148332918e-20

R112_198 V112 V198 671.1212350873438
L112_198 V112 V198 2.0603632960143387e-11
C112_198 V112 V198 -7.486609814167795e-20

R112_199 V112 V199 -352.8768835076013
L112_199 V112 V199 -8.689582350224078e-12
C112_199 V112 V199 -4.336462342178372e-20

R112_200 V112 V200 -9559.56750192971
L112_200 V112 V200 -1.6192846270819578e-11
C112_200 V112 V200 -4.6528848114952975e-20

R113_113 V113 0 -35.73540386493601
L113_113 V113 0 -2.5771599436767017e-12
C113_113 V113 0 6.884118548566624e-19

R113_114 V113 V114 -1132.3462237939573
L113_114 V113 V114 -3.2739474491935235e-12
C113_114 V113 V114 -4.812002861043486e-20

R113_115 V113 V115 102.96462839469307
L113_115 V113 V115 2.3655623044644343e-12
C113_115 V113 V115 1.1732973175496767e-19

R113_116 V113 V116 86.41570186848116
L113_116 V113 V116 5.357393074259364e-12
C113_116 V113 V116 -8.780374324328805e-20

R113_117 V113 V117 179.8702854993219
L113_117 V113 V117 1.4703069794683734e-12
C113_117 V113 V117 3.9764707993528456e-19

R113_118 V113 V118 66.21984224805524
L113_118 V113 V118 1.5334339639289902e-12
C113_118 V113 V118 1.8193002509334534e-19

R113_119 V113 V119 -166.6831780062465
L113_119 V113 V119 -5.0350195866520525e-12
C113_119 V113 V119 1.1689110587245076e-19

R113_120 V113 V120 -90.14914107896936
L113_120 V113 V120 3.5437424639498316e-10
C113_120 V113 V120 2.641437134050023e-19

R113_121 V113 V121 50.4708412258759
L113_121 V113 V121 8.937793406884109e-13
C113_121 V113 V121 4.629813739371218e-19

R113_122 V113 V122 -136.57729230399653
L113_122 V113 V122 -2.513506087077349e-12
C113_122 V113 V122 -2.347845215533564e-19

R113_123 V113 V123 -2602.0551906259507
L113_123 V113 V123 -3.9085584723077945e-12
C113_123 V113 V123 -2.3025720679421404e-19

R113_124 V113 V124 446.50490851461416
L113_124 V113 V124 -2.5744354277539394e-12
C113_124 V113 V124 -2.0549149051773822e-19

R113_125 V113 V125 -791.2429096944537
L113_125 V113 V125 -1.096109717148648e-11
C113_125 V113 V125 -8.683564141568069e-20

R113_126 V113 V126 -63.259617841992615
L113_126 V113 V126 -1.7131013371231168e-12
C113_126 V113 V126 -3.254485241016664e-20

R113_127 V113 V127 -270.7539597702981
L113_127 V113 V127 -2.543139872207886e-10
C113_127 V113 V127 3.613746268631332e-20

R113_128 V113 V128 945.3719210690815
L113_128 V113 V128 5.651614812745455e-12
C113_128 V113 V128 -4.1286905480185295e-20

R113_129 V113 V129 -52.89461378699368
L113_129 V113 V129 -1.0617431823730032e-12
C113_129 V113 V129 -3.474852880912e-19

R113_130 V113 V130 83.19111876204747
L113_130 V113 V130 1.2654526438647725e-12
C113_130 V113 V130 2.846408523612913e-19

R113_131 V113 V131 156.68967370595053
L113_131 V113 V131 4.792273538839742e-12
C113_131 V113 V131 5.528576353507228e-20

R113_132 V113 V132 388.44565836123695
L113_132 V113 V132 3.2249034909750493e-12
C113_132 V113 V132 1.8840290188197165e-19

R113_133 V113 V133 1208.326640987706
L113_133 V113 V133 1.472700970975711e-12
C113_133 V113 V133 1.438527941384307e-19

R113_134 V113 V134 711.6153165459219
L113_134 V113 V134 -2.188546285623832e-12
C113_134 V113 V134 -3.5639888130836996e-19

R113_135 V113 V135 131.4156145418475
L113_135 V113 V135 6.711323638840315e-12
C113_135 V113 V135 -3.771568906464081e-20

R113_136 V113 V136 105.61403337694566
L113_136 V113 V136 -7.798107168552691e-12
C113_136 V113 V136 -1.0399910254062514e-19

R113_137 V113 V137 57.82977637338717
L113_137 V113 V137 -4.072372012050207e-11
C113_137 V113 V137 -2.1713306223740237e-20

R113_138 V113 V138 -201.6659736881069
L113_138 V113 V138 -6.117245984320434e-12
C113_138 V113 V138 9.708650906098563e-20

R113_139 V113 V139 -62.808901415595955
L113_139 V113 V139 -8.96619230750031e-12
C113_139 V113 V139 1.2054231370540898e-19

R113_140 V113 V140 -53.54926523355272
L113_140 V113 V140 -3.258629778968001e-12
C113_140 V113 V140 -8.103953731696304e-20

R113_141 V113 V141 170.46886657387518
L113_141 V113 V141 -6.80830374534086e-12
C113_141 V113 V141 -4.331973957423762e-20

R113_142 V113 V142 -401.4170421390314
L113_142 V113 V142 1.4806122091457801e-12
C113_142 V113 V142 2.0705906942245444e-19

R113_143 V113 V143 -1941.2035882474331
L113_143 V113 V143 -2.7048315458301995e-12
C113_143 V113 V143 -1.784027674305642e-19

R113_144 V113 V144 -571.6280270166294
L113_144 V113 V144 1.0216265701613187e-11
C113_144 V113 V144 1.0943014774414916e-19

R113_145 V113 V145 -51.94107737567301
L113_145 V113 V145 4.84320295104307e-12
C113_145 V113 V145 -4.614495103260606e-21

R113_146 V113 V146 -230.18410575229865
L113_146 V113 V146 -1.9237836820596e-12
C113_146 V113 V146 -1.1605654805032634e-19

R113_147 V113 V147 151.80401401947063
L113_147 V113 V147 3.76064812661543e-12
C113_147 V113 V147 3.82013135899405e-20

R113_148 V113 V148 103.15827577674224
L113_148 V113 V148 1.9578223390897556e-11
C113_148 V113 V148 4.0409074141574435e-20

R113_149 V113 V149 -106.561202266035
L113_149 V113 V149 3.8096329619266995e-12
C113_149 V113 V149 5.444229615737384e-19

R113_150 V113 V150 60.063622344524376
L113_150 V113 V150 5.108399041121909e-12
C113_150 V113 V150 -1.8682669296766488e-19

R113_151 V113 V151 134.5472117328255
L113_151 V113 V151 1.9242377369193897e-12
C113_151 V113 V151 1.8232640662461603e-19

R113_152 V113 V152 -941.2599283778749
L113_152 V113 V152 9.821399012762028e-12
C113_152 V113 V152 -9.561017321816981e-20

R113_153 V113 V153 62.159822877258435
L113_153 V113 V153 -3.2166484474315344e-11
C113_153 V113 V153 -3.111543168555745e-19

R113_154 V113 V154 154.21653523634393
L113_154 V113 V154 8.225039224792321e-12
C113_154 V113 V154 1.7028243856885874e-19

R113_155 V113 V155 -171.02669420927478
L113_155 V113 V155 3.4971170310068575e-11
C113_155 V113 V155 5.0508112322769366e-20

R113_156 V113 V156 155.73795128062486
L113_156 V113 V156 1.7527273508235623e-11
C113_156 V113 V156 7.669481078939068e-21

R113_157 V113 V157 39.709619120976384
L113_157 V113 V157 -3.3513551586254315e-12
C113_157 V113 V157 -5.815243660297739e-19

R113_158 V113 V158 -124.96634475026175
L113_158 V113 V158 3.806622113866983e-11
C113_158 V113 V158 -1.2114531126909648e-19

R113_159 V113 V159 5512.029758637693
L113_159 V113 V159 -2.1800807919525244e-12
C113_159 V113 V159 -1.3062765338602142e-19

R113_160 V113 V160 -210.71361966423322
L113_160 V113 V160 -3.0638177788029912e-12
C113_160 V113 V160 2.421427297529246e-20

R113_161 V113 V161 -55.76017837813185
L113_161 V113 V161 -3.6142457609562102e-12
C113_161 V113 V161 3.1698500849497985e-19

R113_162 V113 V162 -61.853362877636386
L113_162 V113 V162 -1.4985498367549282e-11
C113_162 V113 V162 4.983847799365011e-20

R113_163 V113 V163 -65.82081909053129
L113_163 V113 V163 -1.8988488639824537e-12
C113_163 V113 V163 -1.5313214493980733e-19

R113_164 V113 V164 -59.35545174358807
L113_164 V113 V164 -4.238467580434343e-12
C113_164 V113 V164 4.659530884977249e-20

R113_165 V113 V165 -76.5231719769733
L113_165 V113 V165 8.171175275815033e-13
C113_165 V113 V165 4.0329709123791205e-19

R113_166 V113 V166 80.07582164205134
L113_166 V113 V166 1.8240451815061892e-12
C113_166 V113 V166 2.3813427535676524e-19

R113_167 V113 V167 130.55808941117675
L113_167 V113 V167 2.291597258579025e-12
C113_167 V113 V167 1.2413731647739974e-19

R113_168 V113 V168 421.2411094226966
L113_168 V113 V168 2.6654093109567634e-12
C113_168 V113 V168 8.959212967140089e-20

R113_169 V113 V169 52.42257640289314
L113_169 V113 V169 -1.331918069354611e-12
C113_169 V113 V169 -5.964945487133451e-19

R113_170 V113 V170 86.85166341657404
L113_170 V113 V170 -1.404186294766384e-11
C113_170 V113 V170 -1.7805115850417025e-21

R113_171 V113 V171 77.79524515748165
L113_171 V113 V171 1.2808004731884842e-12
C113_171 V113 V171 2.6157156297438455e-19

R113_172 V113 V172 67.84532590883833
L113_172 V113 V172 4.5681716266277295e-12
C113_172 V113 V172 2.3987058701936804e-20

R113_173 V113 V173 579.6456520442389
L113_173 V113 V173 -3.0324569270154094e-12
C113_173 V113 V173 6.886471189998341e-20

R113_174 V113 V174 -75.69521661517398
L113_174 V113 V174 -1.8207833774423216e-12
C113_174 V113 V174 -4.3360058285849426e-19

R113_175 V113 V175 -118.58152129811282
L113_175 V113 V175 -2.3477259859120812e-12
C113_175 V113 V175 -1.1030795243313198e-19

R113_176 V113 V176 -108.41223908125949
L113_176 V113 V176 -2.3264264206774924e-12
C113_176 V113 V176 -1.5646395408112462e-19

R113_177 V113 V177 -106.10877188825283
L113_177 V113 V177 1.4890279863517223e-12
C113_177 V113 V177 3.8999742044755087e-19

R113_178 V113 V178 -159.77496124415086
L113_178 V113 V178 -4.9692882148070955e-12
C113_178 V113 V178 1.3288109351269972e-20

R113_179 V113 V179 -130.90375133369147
L113_179 V113 V179 -1.379679473563396e-12
C113_179 V113 V179 -2.908659243293889e-19

R113_180 V113 V180 -84.24071163214406
L113_180 V113 V180 -1.878312450814566e-12
C113_180 V113 V180 -8.386554751317037e-20

R113_181 V113 V181 157.35775204705828
L113_181 V113 V181 -2.205010130555387e-12
C113_181 V113 V181 -8.076395857821795e-20

R113_182 V113 V182 59.92165067018631
L113_182 V113 V182 1.0207083353798388e-12
C113_182 V113 V182 2.295102730604513e-19

R113_183 V113 V183 118.43203356259424
L113_183 V113 V183 5.4620344282806795e-11
C113_183 V113 V183 -9.745599860045995e-20

R113_184 V113 V184 91.35122257538539
L113_184 V113 V184 3.5679383550289925e-12
C113_184 V113 V184 -1.4145417074942318e-20

R113_185 V113 V185 163.5422938481423
L113_185 V113 V185 6.7534017771410545e-12
C113_185 V113 V185 -2.223155464355394e-19

R113_186 V113 V186 488.5530545107252
L113_186 V113 V186 2.1476219125929544e-12
C113_186 V113 V186 9.59842249756752e-20

R113_187 V113 V187 -353.41970623453903
L113_187 V113 V187 1.2096046800350323e-12
C113_187 V113 V187 3.1762852870005083e-19

R113_188 V113 V188 6165.7748617622065
L113_188 V113 V188 9.819567161744804e-13
C113_188 V113 V188 3.1878075716354366e-19

R113_189 V113 V189 -115.6888957024554
L113_189 V113 V189 3.133630229506453e-12
C113_189 V113 V189 2.6835946327556156e-19

R113_190 V113 V190 -94.73138429755868
L113_190 V113 V190 -1.6740711631931632e-12
C113_190 V113 V190 -1.6476451117126685e-19

R113_191 V113 V191 -194.32361164826278
L113_191 V113 V191 4.9874861349585e-12
C113_191 V113 V191 2.741379290764066e-19

R113_192 V113 V192 -102.29083529672042
L113_192 V113 V192 -2.040070254356824e-12
C113_192 V113 V192 4.802921700231111e-20

R113_193 V113 V193 -241.0539446467649
L113_193 V113 V193 -1.3939108414868449e-12
C113_193 V113 V193 -2.7300555496865484e-19

R113_194 V113 V194 132.1464292050989
L113_194 V113 V194 -1.8132536030892038e-12
C113_194 V113 V194 -3.3909632797045744e-19

R113_195 V113 V195 158.59902325194
L113_195 V113 V195 -1.5992925139483068e-12
C113_195 V113 V195 -4.20249338637281e-19

R113_196 V113 V196 125.570244070385
L113_196 V113 V196 -1.8158296072670932e-12
C113_196 V113 V196 -4.242890096477289e-19

R113_197 V113 V197 111.44753684523445
L113_197 V113 V197 -9.904818150676237e-12
C113_197 V113 V197 8.220744120452834e-20

R113_198 V113 V198 100.45325143751847
L113_198 V113 V198 1.7325489840467903e-12
C113_198 V113 V198 1.1296002408044241e-19

R113_199 V113 V199 193.34693421030175
L113_199 V113 V199 -3.942009692608162e-11
C113_199 V113 V199 -2.543319680359912e-19

R113_200 V113 V200 353.00652866865414
L113_200 V113 V200 2.781843051260814e-12
C113_200 V113 V200 5.954468219901909e-20

R114_114 V114 0 -60.44734441716447
L114_114 V114 0 1.3810368568436173e-12
C114_114 V114 0 7.303557378367244e-19

R114_115 V114 V115 -259.88370405616655
L114_115 V114 V115 1.3524170644033492e-12
C114_115 V114 V115 3.1228055329408936e-19

R114_116 V114 V116 -325.68540691158205
L114_116 V114 V116 1.5138951231269416e-12
C114_116 V114 V116 2.2996050050931656e-19

R114_117 V114 V117 177.25489096235043
L114_117 V114 V117 3.030837524301157e-12
C114_117 V114 V117 9.712164163397727e-20

R114_118 V114 V118 53.572982712077376
L114_118 V114 V118 1.0762302098403462e-12
C114_118 V114 V118 3.5291895586639264e-19

R114_119 V114 V119 42909.25295175281
L114_119 V114 V119 1.75729077891841e-11
C114_119 V114 V119 2.559800633768559e-19

R114_120 V114 V120 -946.1379958590659
L114_120 V114 V120 3.890429882990837e-12
C114_120 V114 V120 4.655906770279983e-19

R114_121 V114 V121 -223.20429436886548
L114_121 V114 V121 -6.4119279222256225e-09
C114_121 V114 V121 -2.2406011268562533e-20

R114_122 V114 V122 -424.9565917784154
L114_122 V114 V122 1.2138110032083216e-12
C114_122 V114 V122 6.976393311493257e-19

R114_123 V114 V123 186.86029353392075
L114_123 V114 V123 -8.975154477300554e-13
C114_123 V114 V123 -7.721714298291735e-19

R114_124 V114 V124 183.85380628987957
L114_124 V114 V124 -6.702396279065961e-13
C114_124 V114 V124 -9.716037953226041e-19

R114_125 V114 V125 -453.98243045639515
L114_125 V114 V125 2.5842289237709915e-11
C114_125 V114 V125 1.4340121271005839e-19

R114_126 V114 V126 -68.09809435603214
L114_126 V114 V126 -9.32851018062998e-13
C114_126 V114 V126 -4.423977408621091e-19

R114_127 V114 V127 -150.81597418922004
L114_127 V114 V127 5.243256611316829e-12
C114_127 V114 V127 1.6469094401481864e-19

R114_128 V114 V128 -212.68829388331088
L114_128 V114 V128 2.1972470799869666e-12
C114_128 V114 V128 1.0594443186791196e-19

R114_129 V114 V129 199.22090119667072
L114_129 V114 V129 -1.3453927092841233e-11
C114_129 V114 V129 -2.3025295684836224e-19

R114_130 V114 V130 110.32056953108064
L114_130 V114 V130 2.84635472206499e-11
C114_130 V114 V130 -1.4336472740586177e-19

R114_131 V114 V131 218.06037645350875
L114_131 V114 V131 1.4937945988746144e-12
C114_131 V114 V131 4.251980912896127e-19

R114_132 V114 V132 248.35888145939242
L114_132 V114 V132 1.0403656276197638e-12
C114_132 V114 V132 7.493158658977366e-19

R114_133 V114 V133 -503.63791487983303
L114_133 V114 V133 5.7588341738640606e-11
C114_133 V114 V133 1.0892866801252392e-19

R114_134 V114 V134 258.6057249455748
L114_134 V114 V134 2.0762152812801345e-12
C114_134 V114 V134 4.734272628997102e-19

R114_135 V114 V135 190.36909860177386
L114_135 V114 V135 -1.4071320165923497e-12
C114_135 V114 V135 -6.527551391319826e-19

R114_136 V114 V136 137.56882232883652
L114_136 V114 V136 -1.1650903933851797e-12
C114_136 V114 V136 -6.965139492638958e-19

R114_137 V114 V137 -515.3508531386867
L114_137 V114 V137 -3.818478551225004e-12
C114_137 V114 V137 -1.0769891569652287e-19

R114_138 V114 V138 -103.28901007735423
L114_138 V114 V138 -1.4052922531425242e-12
C114_138 V114 V138 -4.562263298459118e-19

R114_139 V114 V139 -81.63106850150837
L114_139 V114 V139 1.8503388520576886e-12
C114_139 V114 V139 6.8716832044322925e-19

R114_140 V114 V140 -61.4490701434628
L114_140 V114 V140 4.746958154675803e-12
C114_140 V114 V140 5.072360780959099e-19

R114_141 V114 V141 260.1422948892122
L114_141 V114 V141 -9.408334770790477e-12
C114_141 V114 V141 -9.304394170207285e-20

R114_142 V114 V142 -292.99007955332235
L114_142 V114 V142 -4.7638103849646586e-11
C114_142 V114 V142 7.344412766982002e-20

R114_143 V114 V143 181.5364541963959
L114_143 V114 V143 -3.533413737221884e-12
C114_143 V114 V143 -9.789156878958887e-20

R114_144 V114 V144 202.81410466186816
L114_144 V114 V144 6.013843918504811e-12
C114_144 V114 V144 4.97590664165342e-20

R114_145 V114 V145 411.3962731721969
L114_145 V114 V145 2.7014293006923277e-12
C114_145 V114 V145 1.0317894826101821e-19

R114_146 V114 V146 45.331506374217035
L114_146 V114 V146 1.2128632397282256e-12
C114_146 V114 V146 1.0049108625220114e-19

R114_147 V114 V147 169.80522605361102
L114_147 V114 V147 -5.8972147657376435e-12
C114_147 V114 V147 -5.981556588198705e-19

R114_148 V114 V148 128.1810744428493
L114_148 V114 V148 -1.5310957603430292e-12
C114_148 V114 V148 -4.406928036293137e-19

R114_149 V114 V149 3750.403091968012
L114_149 V114 V149 3.663344255926166e-12
C114_149 V114 V149 2.0758110238151206e-19

R114_150 V114 V150 -379.7124482706295
L114_150 V114 V150 -2.0082928767008887e-12
C114_150 V114 V150 -2.6511171535500704e-20

R114_151 V114 V151 -376.8909236040732
L114_151 V114 V151 2.847552219760709e-12
C114_151 V114 V151 2.7708590708233896e-19

R114_152 V114 V152 -157.16314050406004
L114_152 V114 V152 1.908290198028213e-12
C114_152 V114 V152 1.0913462945844482e-19

R114_153 V114 V153 -151.74520101066335
L114_153 V114 V153 -3.3931290984794235e-12
C114_153 V114 V153 -2.242638290829418e-19

R114_154 V114 V154 -47.82158575627377
L114_154 V114 V154 -6.4151469827395e-12
C114_154 V114 V154 -1.7140771059451233e-19

R114_155 V114 V155 -110.30704341101793
L114_155 V114 V155 1.719039707321403e-12
C114_155 V114 V155 3.137901251153139e-19

R114_156 V114 V156 -594.3867055325187
L114_156 V114 V156 -5.094261707989507e-12
C114_156 V114 V156 2.8580475866956907e-19

R114_157 V114 V157 -186.91527537276028
L114_157 V114 V157 -1.8438383596657313e-12
C114_157 V114 V157 -2.719521302423618e-19

R114_158 V114 V158 67.77037107630584
L114_158 V114 V158 1.39704603899426e-12
C114_158 V114 V158 2.293900022344392e-19

R114_159 V114 V159 123.05683174478236
L114_159 V114 V159 -1.2567364121905209e-12
C114_159 V114 V159 -4.0001247514169215e-19

R114_160 V114 V160 202.0510454263096
L114_160 V114 V160 -2.826540121903983e-12
C114_160 V114 V160 -2.7848370014186754e-19

R114_161 V114 V161 427.5720721043483
L114_161 V114 V161 1.2221442049494922e-12
C114_161 V114 V161 3.8489043247221434e-19

R114_162 V114 V162 60.032105699283115
L114_162 V114 V162 8.110046683049052e-12
C114_162 V114 V162 6.664564415166978e-21

R114_163 V114 V163 -1269.1183778449065
L114_163 V114 V163 2.651877836891148e-12
C114_163 V114 V163 2.1237499315848314e-19

R114_164 V114 V164 -3290.4175291777537
L114_164 V114 V164 3.668867542584501e-12
C114_164 V114 V164 2.7302733758130344e-19

R114_165 V114 V165 109.2403431546345
L114_165 V114 V165 -6.470390430262479e-12
C114_165 V114 V165 -1.4658832386838913e-19

R114_166 V114 V166 -51.49179147958555
L114_166 V114 V166 -1.1978860186646958e-12
C114_166 V114 V166 -1.1823051656653282e-19

R114_167 V114 V167 254.83077505195598
L114_167 V114 V167 3.1742266685837587e-12
C114_167 V114 V167 1.4165014171747932e-19

R114_168 V114 V168 354.7912609879198
L114_168 V114 V168 1.3138674214182214e-12
C114_168 V114 V168 1.5311068269702732e-19

R114_169 V114 V169 -1388.8081801179524
L114_169 V114 V169 -1.679252094868373e-12
C114_169 V114 V169 -4.33110434122365e-19

R114_170 V114 V170 -491.9616683132707
L114_170 V114 V170 1.11524001359579e-12
C114_170 V114 V170 8.557654169706788e-20

R114_171 V114 V171 -2165.1806883661698
L114_171 V114 V171 -9.75643770654004e-12
C114_171 V114 V171 -1.913229998745775e-19

R114_172 V114 V172 -2458.9725370181195
L114_172 V114 V172 -1.1747506818478593e-12
C114_172 V114 V172 -2.264540378293327e-19

R114_173 V114 V173 -174.5640396671815
L114_173 V114 V173 1.597294614192313e-12
C114_173 V114 V173 2.20237464111859e-19

R114_174 V114 V174 52.39623032653756
L114_174 V114 V174 -4.584245876741775e-12
C114_174 V114 V174 -2.264748320430642e-19

R114_175 V114 V175 -428.0610084599818
L114_175 V114 V175 8.807648961725353e-12
C114_175 V114 V175 2.304614225336068e-19

R114_176 V114 V176 -197.3885459018641
L114_176 V114 V176 3.3404850752513813e-12
C114_176 V114 V176 2.332010879089682e-19

R114_177 V114 V177 384.1501397154306
L114_177 V114 V177 -3.567495785154753e-12
C114_177 V114 V177 -3.141123881487097e-20

R114_178 V114 V178 -362.55938575958027
L114_178 V114 V178 -1.7806945421621296e-12
C114_178 V114 V178 1.3431460629308983e-19

R114_179 V114 V179 -599.4209333015586
L114_179 V114 V179 -7.261938094750882e-12
C114_179 V114 V179 -2.449334879784552e-19

R114_180 V114 V180 611.3793210360407
L114_180 V114 V180 1.7891237276004175e-11
C114_180 V114 V180 -2.5671755205664916e-19

R114_181 V114 V181 372.32980867167817
L114_181 V114 V181 4.3098395882224816e-12
C114_181 V114 V181 1.65901740969411e-19

R114_182 V114 V182 -116.26167761287246
L114_182 V114 V182 1.7740616973725904e-12
C114_182 V114 V182 7.918918627095255e-21

R114_183 V114 V183 374.71195700664117
L114_183 V114 V183 -2.2817062775437886e-12
C114_183 V114 V183 -1.6421980867293363e-20

R114_184 V114 V184 636.0278131242326
L114_184 V114 V184 -1.92959937111384e-12
C114_184 V114 V184 5.404458921789963e-20

R114_185 V114 V185 -227.58325663820466
L114_185 V114 V185 2.955828284318957e-12
C114_185 V114 V185 -4.356587333404106e-20

R114_186 V114 V186 333.86759991522854
L114_186 V114 V186 -1.5160960521321868e-12
C114_186 V114 V186 -1.593795037371592e-19

R114_187 V114 V187 962.5283319318504
L114_187 V114 V187 1.8545459516435555e-12
C114_187 V114 V187 3.6120523024495515e-19

R114_188 V114 V188 -505.9350925388044
L114_188 V114 V188 7.628216793886855e-13
C114_188 V114 V188 3.01188811612487e-19

R114_189 V114 V189 1446.8869547318823
L114_189 V114 V189 -1.5771046977557305e-12
C114_189 V114 V189 -2.61640782518861e-19

R114_190 V114 V190 111.15367253031425
L114_190 V114 V190 -6.9898589512424124e-12
C114_190 V114 V190 1.101646835879937e-19

R114_191 V114 V191 -1066.019150928197
L114_191 V114 V191 2.153185778458832e-12
C114_191 V114 V191 -2.811333388530075e-19

R114_192 V114 V192 -840.6655813030668
L114_192 V114 V192 -2.189483604514261e-12
C114_192 V114 V192 -4.708090021621246e-19

R114_193 V114 V193 418.6785072174013
L114_193 V114 V193 3.517342344037739e-11
C114_193 V114 V193 -1.0836808137499687e-20

R114_194 V114 V194 -262.8992581162801
L114_194 V114 V194 -3.4709030780462948e-12
C114_194 V114 V194 -4.383548742649217e-19

R114_195 V114 V195 -174058.72768694328
L114_195 V114 V195 -1.8491193786549433e-12
C114_195 V114 V195 1.9743685794546942e-19

R114_196 V114 V196 446.1648165051814
L114_196 V114 V196 1.745998209559842e-11
C114_196 V114 V196 4.527041226413051e-19

R114_197 V114 V197 -274.407323157074
L114_197 V114 V197 1.8194917826493072e-12
C114_197 V114 V197 2.921449822262286e-19

R114_198 V114 V198 -196.42180237125731
L114_198 V114 V198 4.35565375527848e-12
C114_198 V114 V198 -3.575414836605102e-21

R114_199 V114 V199 998.1157700569652
L114_199 V114 V199 4.30047193258892e-12
C114_199 V114 V199 1.4361109479869892e-19

R114_200 V114 V200 -772.4863114383791
L114_200 V114 V200 4.102118877268766e-12
C114_200 V114 V200 1.805207585077442e-19

R115_115 V115 0 -737.2076232304449
L115_115 V115 0 -3.426239640409248e-13
C115_115 V115 0 -1.7680674099580215e-18

R115_116 V115 V116 -170.88580186239133
L115_116 V115 V116 5.4385828003724135e-12
C115_116 V115 V116 2.5747773580074123e-19

R115_117 V115 V117 465.7215298118392
L115_117 V115 V117 -1.533146533532536e-12
C115_117 V115 V117 -3.3502272235902846e-19

R115_118 V115 V118 -1562.1671440938312
L115_118 V115 V118 -1.2503279663031624e-12
C115_118 V115 V118 -2.831224741539512e-19

R115_119 V115 V119 95.65951304191454
L115_119 V115 V119 2.2011008001417476e-12
C115_119 V115 V119 1.1670601211611398e-19

R115_120 V115 V120 3178.95272672334
L115_120 V115 V120 -6.625710962082421e-12
C115_120 V115 V120 -2.3795343265575842e-20

R115_121 V115 V121 -90.0959185852353
L115_121 V115 V121 -3.9703214007860785e-12
C115_121 V115 V121 8.366098392121295e-20

R115_122 V115 V122 422.9847143056528
L115_122 V115 V122 1.7184622052362738e-11
C115_122 V115 V122 4.2807726152808125e-20

R115_123 V115 V123 10659.782379639772
L115_123 V115 V123 4.3628851749661413e-13
C115_123 V115 V123 9.770801207047684e-19

R115_124 V115 V124 195.02402564719495
L115_124 V115 V124 -4.011839969073808e-12
C115_124 V115 V124 -3.4459140705365675e-19

R115_125 V115 V125 -1303.0703278724943
L115_125 V115 V125 2.5637456433112194e-12
C115_125 V115 V125 1.4652544271452408e-19

R115_126 V115 V126 283.5813776623708
L115_126 V115 V126 1.2116154563307598e-12
C115_126 V115 V126 2.2015252027933513e-19

R115_127 V115 V127 -120.56843306239459
L115_127 V115 V127 -8.4408077784699e-13
C115_127 V115 V127 -3.7973160231480573e-19

R115_128 V115 V128 -411.9926714367319
L115_128 V115 V128 1.940813353094398e-12
C115_128 V115 V128 3.269536856367539e-19

R115_129 V115 V129 90.23006738869051
L115_129 V115 V129 1.257206527683276e-12
C115_129 V115 V129 2.8317943988327353e-19

R115_130 V115 V130 -225.7682784793323
L115_130 V115 V130 -1.2724705188229852e-12
C115_130 V115 V130 -2.646522313082244e-19

R115_131 V115 V131 137.65951908927894
L115_131 V115 V131 -1.6550540155045809e-12
C115_131 V115 V131 -4.1597582766971625e-19

R115_132 V115 V132 -6496.931707986302
L115_132 V115 V132 -1.2970097837573496e-12
C115_132 V115 V132 -3.1105940961730627e-19

R115_133 V115 V133 -526.1620201165292
L115_133 V115 V133 -1.161857790003749e-12
C115_133 V115 V133 -3.729983219747813e-19

R115_134 V115 V134 1402.5352488133137
L115_134 V115 V134 2.1794007233058774e-12
C115_134 V115 V134 3.49042276413461e-19

R115_135 V115 V135 -228.24617044762664
L115_135 V115 V135 7.57017495335653e-13
C115_135 V115 V135 7.698799337478208e-19

R115_136 V115 V136 336.42804487329596
L115_136 V115 V136 -1.9443857860048435e-12
C115_136 V115 V136 -2.7465795826815153e-19

R115_137 V115 V137 -118.553095244473
L115_137 V115 V137 -1.1989802589159544e-12
C115_137 V115 V137 -3.151037192700583e-19

R115_138 V115 V138 -1423.3036700951543
L115_138 V115 V138 5.483021567966485e-12
C115_138 V115 V138 -1.1561042945799414e-19

R115_139 V115 V139 1367.3650956112851
L115_139 V115 V139 -5.703839831633375e-13
C115_139 V115 V139 -8.052665384174698e-19

R115_140 V115 V140 -238.33895427731326
L115_140 V115 V140 1.3148288359299717e-12
C115_140 V115 V140 3.7948912235457907e-19

R115_141 V115 V141 -5406.664339289711
L115_141 V115 V141 6.808568912851341e-13
C115_141 V115 V141 7.1860845902861605e-19

R115_142 V115 V142 -894.9756920584192
L115_142 V115 V142 -1.8058651072555982e-12
C115_142 V115 V142 -1.4117399925097635e-19

R115_143 V115 V143 113.76746672900977
L115_143 V115 V143 9.937067378443678e-13
C115_143 V115 V143 2.0057013422939327e-19

R115_144 V115 V144 815.3549240308371
L115_144 V115 V144 1.8686435726310424e-11
C115_144 V115 V144 -4.9864752453868115e-21

R115_145 V115 V145 98.50555126135927
L115_145 V115 V145 1.0731347519933718e-12
C115_145 V115 V145 2.802553432008483e-19

R115_146 V115 V146 97.12524868892504
L115_146 V115 V146 1.854170101304134e-12
C115_146 V115 V146 4.346057202283398e-22

R115_147 V115 V147 -134.5759826334056
L115_147 V115 V147 1.864810500351883e-12
C115_147 V115 V147 4.9461900283075005e-19

R115_148 V115 V148 141.1506985778215
L115_148 V115 V148 -9.28080118342727e-12
C115_148 V115 V148 -1.173104613638795e-19

R115_149 V115 V149 445.0952424314446
L115_149 V115 V149 -3.872668710792723e-13
C115_149 V115 V149 -9.823169199846664e-19

R115_150 V115 V150 -190.8594768302676
L115_150 V115 V150 1.0012628072796543e-11
C115_150 V115 V150 5.031915028805828e-19

R115_151 V115 V151 -203.81177997212228
L115_151 V115 V151 -1.4413925507745854e-12
C115_151 V115 V151 -2.547390175016558e-19

R115_152 V115 V152 -834.8640560526544
L115_152 V115 V152 2.4903451349800583e-12
C115_152 V115 V152 1.0815637756757841e-19

R115_153 V115 V153 -105.0288892646185
L115_153 V115 V153 -3.028897804710367e-12
C115_153 V115 V153 -7.649396466851072e-20

R115_154 V115 V154 -85.37918978294591
L115_154 V115 V154 -3.610939630809695e-12
C115_154 V115 V154 -3.4978785387265386e-19

R115_155 V115 V155 -108.53170824953395
L115_155 V115 V155 -6.278771037619204e-13
C115_155 V115 V155 -4.593644317349118e-19

R115_156 V115 V156 -159.7020829085633
L115_156 V115 V156 -2.179644908862245e-12
C115_156 V115 V156 2.6894670477932516e-20

R115_157 V115 V157 -76.81090183074554
L115_157 V115 V157 5.696785957991092e-13
C115_157 V115 V157 7.000562415727898e-19

R115_158 V115 V158 123.1745003347785
L115_158 V115 V158 -2.308235529081832e-12
C115_158 V115 V158 -4.007894630749621e-20

R115_159 V115 V159 61.46878157847038
L115_159 V115 V159 5.363453140018419e-13
C115_159 V115 V159 3.192555625450022e-19

R115_160 V115 V160 -570.0227195196437
L115_160 V115 V160 -2.315169593595786e-12
C115_160 V115 V160 -2.7309950663069443e-19

R115_161 V115 V161 104.072587276939
L115_161 V115 V161 6.163699565419074e-12
C115_161 V115 V161 1.160795366172234e-19

R115_162 V115 V162 86.10687341615736
L115_162 V115 V162 -3.131576345484103e-12
C115_162 V115 V162 -1.7123836507377295e-19

R115_163 V115 V163 111.69196320379857
L115_163 V115 V163 -2.0801589456649242e-12
C115_163 V115 V163 -2.008430484930254e-19

R115_164 V115 V164 72.68843703573475
L115_164 V115 V164 1.8236620713302733e-12
C115_164 V115 V164 5.705676380346887e-20

R115_165 V115 V165 84.9268813365807
L115_165 V115 V165 -1.926977355460023e-12
C115_165 V115 V165 -2.6517543298689565e-19

R115_166 V115 V166 -110.96782964459572
L115_166 V115 V166 3.098570838349725e-12
C115_166 V115 V166 1.3681499811014996e-19

R115_167 V115 V167 -94.18692457122249
L115_167 V115 V167 -1.001095158062666e-11
C115_167 V115 V167 2.5656314928407565e-19

R115_168 V115 V168 -483.32754578282567
L115_168 V115 V168 2.0377744457528074e-11
C115_168 V115 V168 2.046843912647188e-19

R115_169 V115 V169 -138.1114905791811
L115_169 V115 V169 9.287721494647042e-11
C115_169 V115 V169 4.195595738437434e-20

R115_170 V115 V170 -474.70257601780014
L115_170 V115 V170 -4.301799319923804e-12
C115_170 V115 V170 -1.4994763269413575e-19

R115_171 V115 V171 -109.42246705617038
L115_171 V115 V171 1.1079866446698795e-10
C115_171 V115 V171 -2.0463648219199313e-19

R115_172 V115 V172 -161.4050045126615
L115_172 V115 V172 -1.8777396552725932e-12
C115_172 V115 V172 -2.0567489780208015e-19

R115_173 V115 V173 -195.8720985641223
L115_173 V115 V173 6.907350285561547e-11
C115_173 V115 V173 -9.110507269089883e-20

R115_174 V115 V174 195.01659281290785
L115_174 V115 V174 -2.9722896993776394e-12
C115_174 V115 V174 1.198508234360541e-19

R115_175 V115 V175 78.50403066584587
L115_175 V115 V175 -7.284130063271003e-13
C115_175 V115 V175 -5.436213188467146e-19

R115_176 V115 V176 540.2806482894482
L115_176 V115 V176 3.2171433411358053e-11
C115_176 V115 V176 -2.5978171991021378e-20

R115_177 V115 V177 142.48670088142566
L115_177 V115 V177 3.2656455484672753e-12
C115_177 V115 V177 2.56106144618787e-20

R115_178 V115 V178 518.8361644567211
L115_178 V115 V178 1.4293351646976808e-12
C115_178 V115 V178 7.206332006087241e-20

R115_179 V115 V179 611.202210069753
L115_179 V115 V179 1.1230755985608428e-12
C115_179 V115 V179 6.447660693285585e-19

R115_180 V115 V180 669.659852748203
L115_180 V115 V180 1.2329528256738458e-12
C115_180 V115 V180 1.5825875981270312e-19

R115_181 V115 V181 -511.99364965898536
L115_181 V115 V181 -7.537690443068102e-12
C115_181 V115 V181 3.2147619557860407e-19

R115_182 V115 V182 -129.88417123993554
L115_182 V115 V182 -8.511985208046201e-13
C115_182 V115 V182 -2.429327859581691e-19

R115_183 V115 V183 -133.70641821720548
L115_183 V115 V183 8.165756567331111e-13
C115_183 V115 V183 6.1743999017980715e-21

R115_184 V115 V184 -2116.766228323433
L115_184 V115 V184 3.715931525845313e-12
C115_184 V115 V184 9.046856172490996e-20

R115_185 V115 V185 -193.77106969797885
L115_185 V115 V185 -1.0159648410771918e-10
C115_185 V115 V185 -2.0864698012114807e-19

R115_186 V115 V186 -5677.52219028669
L115_186 V115 V186 1.0725323031690221e-11
C115_186 V115 V186 2.6894267990323826e-19

R115_187 V115 V187 584.3981425463761
L115_187 V115 V187 -5.382196370771949e-13
C115_187 V115 V187 -5.479013766786095e-19

R115_188 V115 V188 -778.0975844723912
L115_188 V115 V188 -1.5587476586776083e-12
C115_188 V115 V188 -1.1604267145080583e-19

R115_189 V115 V189 214.5732191082226
L115_189 V115 V189 -3.6030312148687817e-12
C115_189 V115 V189 -2.5394019352520474e-19

R115_190 V115 V190 157.82547242334368
L115_190 V115 V190 2.1756923364758536e-12
C115_190 V115 V190 1.6914208451781055e-19

R115_191 V115 V191 153.87600319738115
L115_191 V115 V191 -1.742373822213925e-12
C115_191 V115 V191 1.5225802550884783e-19

R115_192 V115 V192 914.7465136958224
L115_192 V115 V192 -1.394345475859106e-12
C115_192 V115 V192 -3.6076896697677273e-19

R115_193 V115 V193 512.4735122544131
L115_193 V115 V193 1.3819951523048863e-11
C115_193 V115 V193 8.807623817070768e-20

R115_194 V115 V194 -240.67597018940185
L115_194 V115 V194 -2.359901115160766e-12
C115_194 V115 V194 -8.554502582323178e-20

R115_195 V115 V195 -178.168962711619
L115_195 V115 V195 8.492567106207714e-13
C115_195 V115 V195 -8.646014843464676e-20

R115_196 V115 V196 446.7849070303413
L115_196 V115 V196 5.473858924615044e-13
C115_196 V115 V196 7.549530926806196e-19

R115_197 V115 V197 -226.0649999338486
L115_197 V115 V197 1.848388376631931e-12
C115_197 V115 V197 2.8473582217422523e-19

R115_198 V115 V198 -322.2106599529057
L115_198 V115 V198 -3.4274472153352325e-12
C115_198 V115 V198 -3.825517514739585e-20

R115_199 V115 V199 -349.4519054520155
L115_199 V115 V199 4.742919569781428e-12
C115_199 V115 V199 5.905579768917708e-20

R115_200 V115 V200 -299.6627088687777
L115_200 V115 V200 -1.3059420823803162e-11
C115_200 V115 V200 -7.482747268435066e-20

R116_116 V116 0 99.69209170924319
L116_116 V116 0 -2.2358492224976316e-13
C116_116 V116 0 -1.4408362623589724e-18

R116_117 V116 V117 797.8990494023354
L116_117 V116 V117 -2.3395777032101558e-12
C116_117 V116 V117 -1.7143000499176847e-19

R116_118 V116 V118 -460.2925974386202
L116_118 V116 V118 -4.50625745884852e-12
C116_118 V116 V118 6.376267183816276e-20

R116_119 V116 V119 -1567.3130305165644
L116_119 V116 V119 -3.3967572742086363e-12
C116_119 V116 V119 -6.603590466315348e-20

R116_120 V116 V120 59.77126651360031
L116_120 V116 V120 1.6206192959228815e-11
C116_120 V116 V120 -1.4725877322940901e-19

R116_121 V116 V121 -94.55849555237758
L116_121 V116 V121 -2.44352179755297e-10
C116_121 V116 V121 2.178667263700293e-19

R116_122 V116 V122 284.8713702157621
L116_122 V116 V122 -2.763080297653614e-12
C116_122 V116 V122 -2.2354937361416593e-19

R116_123 V116 V123 171.1436277284266
L116_123 V116 V123 -2.8357557424437544e-12
C116_123 V116 V123 -4.430943970865746e-19

R116_124 V116 V124 -257.91355444141135
L116_124 V116 V124 4.106063090672827e-13
C116_124 V116 V124 1.2075365679231727e-18

R116_125 V116 V125 4580.513831948226
L116_125 V116 V125 2.379224457669828e-12
C116_125 V116 V125 1.3623189416206272e-19

R116_126 V116 V126 212.60511572114854
L116_126 V116 V126 1.920046265801357e-12
C116_126 V116 V126 3.506889678244664e-20

R116_127 V116 V127 1085.5807552774952
L116_127 V116 V127 1.142652423113865e-12
C116_127 V116 V127 4.286357456297961e-19

R116_128 V116 V128 -104.4526729245216
L116_128 V116 V128 -1.1333589793770704e-12
C116_128 V116 V128 -3.055643836450237e-19

R116_129 V116 V129 99.60879455338427
L116_129 V116 V129 4.4221749134209775e-12
C116_129 V116 V129 -7.805257755586397e-20

R116_130 V116 V130 -189.4046206811627
L116_130 V116 V130 -4.239670814211447e-12
C116_130 V116 V130 4.0197357284298593e-20

R116_131 V116 V131 -251.2894854215218
L116_131 V116 V131 -2.467965424900627e-12
C116_131 V116 V131 -6.227031836363289e-20

R116_132 V116 V132 95.2895893166809
L116_132 V116 V132 -9.73375781382758e-13
C116_132 V116 V132 -5.339178143369284e-19

R116_133 V116 V133 -3177.648163248781
L116_133 V116 V133 -1.9827014868729317e-12
C116_133 V116 V133 -2.0619152709751658e-19

R116_134 V116 V134 505.94269664307205
L116_134 V116 V134 -3.3951479827400245e-12
C116_134 V116 V134 -1.9560316429930277e-19

R116_135 V116 V135 377.6881802754084
L116_135 V116 V135 -1.263081730878759e-12
C116_135 V116 V135 -5.689119902750049e-19

R116_136 V116 V136 -208.79956501953507
L116_136 V116 V136 8.427827468640757e-13
C116_136 V116 V136 7.14035073557715e-19

R116_137 V116 V137 -105.31782704429192
L116_137 V116 V137 -3.6138893692663884e-12
C116_137 V116 V137 3.5940124975719496e-20

R116_138 V116 V138 -784.7109684031944
L116_138 V116 V138 3.105070614453435e-12
C116_138 V116 V138 1.0052467367677003e-19

R116_139 V116 V139 -351.73487862823714
L116_139 V116 V139 9.471744995041057e-13
C116_139 V116 V139 7.237323542521071e-19

R116_140 V116 V140 951.8783899521401
L116_140 V116 V140 -1.1457167385808726e-12
C116_140 V116 V140 -6.057512262408828e-19

R116_141 V116 V141 -1811.2721210576167
L116_141 V116 V141 1.5821316880396798e-12
C116_141 V116 V141 2.0959955614590216e-19

R116_142 V116 V142 -1118.3801965609882
L116_142 V116 V142 7.0468901910940725e-12
C116_142 V116 V142 3.912040089717187e-20

R116_143 V116 V143 408.72917388572336
L116_143 V116 V143 -7.014869036180037e-12
C116_143 V116 V143 -1.464551760084833e-19

R116_144 V116 V144 114.68100646466975
L116_144 V116 V144 4.755998847208243e-12
C116_144 V116 V144 8.975334991633527e-20

R116_145 V116 V145 89.80849575223945
L116_145 V116 V145 2.213590128293085e-12
C116_145 V116 V145 -1.0286785890420777e-20

R116_146 V116 V146 92.66779696150722
L116_146 V116 V146 -3.473799433540524e-12
C116_146 V116 V146 -7.957395755587375e-20

R116_147 V116 V147 334.4565531849168
L116_147 V116 V147 1.1856821900569809e-11
C116_147 V116 V147 -2.1481280453415934e-19

R116_148 V116 V148 -113.28097144875302
L116_148 V116 V148 7.961181412921712e-13
C116_148 V116 V148 4.482832510243333e-19

R116_149 V116 V149 291.8415412878227
L116_149 V116 V149 -1.5963980508196078e-12
C116_149 V116 V149 2.9266492059721924e-20

R116_150 V116 V150 -160.56112702111326
L116_150 V116 V150 2.5588445926464123e-12
C116_150 V116 V150 1.4474678078108266e-19

R116_151 V116 V151 -1012.1488084109569
L116_151 V116 V151 -4.053068056766161e-10
C116_151 V116 V151 1.8416705407974684e-19

R116_152 V116 V152 -149.89580649021593
L116_152 V116 V152 -6.971496133822589e-13
C116_152 V116 V152 -1.8323706912719136e-19

R116_153 V116 V153 -85.9280512886229
L116_153 V116 V153 -1.382966187188756e-12
C116_153 V116 V153 -1.8196517305967806e-19

R116_154 V116 V154 -82.87668715572053
L116_154 V116 V154 -1.612886322093996e-12
C116_154 V116 V154 -3.9075406594208264e-20

R116_155 V116 V155 -96.44304729984096
L116_155 V116 V155 -7.201132605913823e-12
C116_155 V116 V155 1.7248679131515877e-19

R116_156 V116 V156 -405.4751556920796
L116_156 V116 V156 2.8255534587162677e-12
C116_156 V116 V156 -3.4872729142948105e-19

R116_157 V116 V157 -73.50700488808373
L116_157 V116 V157 1.2563818161764375e-12
C116_157 V116 V157 9.601897675351413e-20

R116_158 V116 V158 159.99657696484263
L116_158 V116 V158 1.0081214568920237e-11
C116_158 V116 V158 -2.066835266589646e-20

R116_159 V116 V159 672.666170553303
L116_159 V116 V159 -1.871285920689599e-12
C116_159 V116 V159 -3.173618748070748e-19

R116_160 V116 V160 65.51327536090385
L116_160 V116 V160 1.047531877786092e-12
C116_160 V116 V160 2.2803412123304985e-19

R116_161 V116 V161 124.33885030071005
L116_161 V116 V161 -5.9113853281901105e-12
C116_161 V116 V161 6.515646578590921e-20

R116_162 V116 V162 90.60871330304394
L116_162 V116 V162 3.807579141382991e-11
C116_162 V116 V162 -4.954187202469227e-20

R116_163 V116 V163 117.60362606618844
L116_163 V116 V163 2.2258813285893457e-12
C116_163 V116 V163 8.294468789603468e-20

R116_164 V116 V164 125.72542884895917
L116_164 V116 V164 -2.3575780685277142e-12
C116_164 V116 V164 -1.978563860739344e-19

R116_165 V116 V165 87.71963737904504
L116_165 V116 V165 1.5372278750132505e-12
C116_165 V116 V165 1.4962117476601e-19

R116_166 V116 V166 -125.58178359383479
L116_166 V116 V166 2.078414113850171e-12
C116_166 V116 V166 1.5818261130242403e-19

R116_167 V116 V167 -5980.127907881491
L116_167 V116 V167 6.009414701068814e-11
C116_167 V116 V167 3.6256832102344276e-20

R116_168 V116 V168 -75.81226542405481
L116_168 V116 V168 -1.6643027252328156e-12
C116_168 V116 V168 2.1953240544299885e-19

R116_169 V116 V169 -136.344065406599
L116_169 V116 V169 -4.493787336585429e-12
C116_169 V116 V169 -4.5004809224307463e-20

R116_170 V116 V170 -256.6232439975383
L116_170 V116 V170 -2.1308412305034925e-12
C116_170 V116 V170 3.676822506080552e-20

R116_171 V116 V171 -151.82965589161324
L116_171 V116 V171 -2.163021387975148e-12
C116_171 V116 V171 2.4299910388148398e-20

R116_172 V116 V172 -131.5722574462662
L116_172 V116 V172 9.501762910310367e-13
C116_172 V116 V172 -2.936481275957199e-22

R116_173 V116 V173 -149.41926128456302
L116_173 V116 V173 -2.5288337867718565e-12
C116_173 V116 V173 -1.7365383772189586e-19

R116_174 V116 V174 156.02997371384544
L116_174 V116 V174 -3.8710043381340756e-12
C116_174 V116 V174 -1.2941815804671255e-19

R116_175 V116 V175 755.5723619406916
L116_175 V116 V175 1.995742150830941e-12
C116_175 V116 V175 9.69734188383081e-20

R116_176 V116 V176 87.07870460238956
L116_176 V116 V176 -7.666969708048567e-13
C116_176 V116 V176 -5.671908558406928e-19

R116_177 V116 V177 157.91837869782057
L116_177 V116 V177 2.8559164747359418e-12
C116_177 V116 V177 1.2451684237073251e-19

R116_178 V116 V178 978.7629688620538
L116_178 V116 V178 1.979186214988018e-12
C116_178 V116 V178 -3.9822356543070545e-20

R116_179 V116 V179 -639.9437363424378
L116_179 V116 V179 3.065110470895366e-12
C116_179 V116 V179 -1.4882655050639011e-19

R116_180 V116 V180 85.91615934821878
L116_180 V116 V180 2.398003035864765e-12
C116_180 V116 V180 4.038492445084058e-19

R116_181 V116 V181 -1378.757163226593
L116_181 V116 V181 9.939280196266208e-12
C116_181 V116 V181 2.1337240175648958e-19

R116_182 V116 V182 -131.88358168297495
L116_182 V116 V182 -6.211432316199867e-12
C116_182 V116 V182 9.079015032171577e-20

R116_183 V116 V183 270.96485483237075
L116_183 V116 V183 -3.2869988138000356e-11
C116_183 V116 V183 1.0666754454696298e-19

R116_184 V116 V184 -76.82952333604786
L116_184 V116 V184 1.1008775788947673e-12
C116_184 V116 V184 -6.728386834189803e-20

R116_185 V116 V185 -149.14872450139285
L116_185 V116 V185 2.5087038900488525e-11
C116_185 V116 V185 -1.9838743584644032e-19

R116_186 V116 V186 767.4136757067331
L116_186 V116 V186 2.555858227206136e-12
C116_186 V116 V186 8.747441802637214e-20

R116_187 V116 V187 431.1375619319829
L116_187 V116 V187 2.039571937757332e-12
C116_187 V116 V187 1.386707145536977e-19

R116_188 V116 V188 -207.383103061902
L116_188 V116 V188 -6.009216514730026e-13
C116_188 V116 V188 -1.4396353021063623e-19

R116_189 V116 V189 254.29716644832948
L116_189 V116 V189 -6.918336937489457e-12
C116_189 V116 V189 -5.08801512676449e-20

R116_190 V116 V190 224.96275900278317
L116_190 V116 V190 8.717390721948859e-12
C116_190 V116 V190 -2.4026556616859968e-20

R116_191 V116 V191 -226.38370179337093
L116_191 V116 V191 -1.5400131152390642e-12
C116_191 V116 V191 -2.4680288898144554e-19

R116_192 V116 V192 87.29293562204343
L116_192 V116 V192 1.354319120774373e-12
C116_192 V116 V192 2.270059333565757e-19

R116_193 V116 V193 209.23695859651644
L116_193 V116 V193 -2.1239527869763522e-11
C116_193 V116 V193 2.473814710326809e-20

R116_194 V116 V194 -255.3476546439585
L116_194 V116 V194 -7.153971740676247e-12
C116_194 V116 V194 1.7242281569486917e-20

R116_195 V116 V195 749.2680119766856
L116_195 V116 V195 1.0474113655589941e-12
C116_195 V116 V195 5.1476900482264285e-19

R116_196 V116 V196 -167.16017483205772
L116_196 V116 V196 -1.6107379172360853e-12
C116_196 V116 V196 -6.49552196809086e-19

R116_197 V116 V197 -223.13881368331528
L116_197 V116 V197 8.604368696922886e-12
C116_197 V116 V197 7.321295533568129e-20

R116_198 V116 V198 -342.29235031554146
L116_198 V116 V198 -4.0483172340659667e-11
C116_198 V116 V198 1.1904805441336903e-19

R116_199 V116 V199 1656.0851864763056
L116_199 V116 V199 -1.3300283783809806e-11
C116_199 V116 V199 -7.712092028736937e-20

R116_200 V116 V200 -172.24979032273384
L116_200 V116 V200 3.809014098938385e-12
C116_200 V116 V200 1.8085813431052168e-19

R117_117 V117 0 94.95053668596104
L117_117 V117 0 -2.6204464272475574e-13
C117_117 V117 0 -1.875372641869164e-18

R117_118 V117 V118 -120.98051382020412
L117_118 V117 V118 -1.7665212116661966e-12
C117_118 V117 V118 -2.2626521631941997e-19

R117_119 V117 V119 2401.873220160977
L117_119 V117 V119 1.2415523264532495e-11
C117_119 V117 V119 -2.5654784323190172e-20

R117_120 V117 V120 235.11584645267428
L117_120 V117 V120 2.914906726208221e-10
C117_120 V117 V120 -1.8688774857541252e-19

R117_121 V117 V121 162.5750422412361
L117_121 V117 V121 1.2093446290412414e-11
C117_121 V117 V121 1.8486434967332167e-19

R117_122 V117 V122 349.9328215280831
L117_122 V117 V122 3.775932033013099e-12
C117_122 V117 V122 1.6642474343494021e-19

R117_123 V117 V123 -542.5542231618613
L117_123 V117 V123 2.5253234746755586e-12
C117_123 V117 V123 2.5933271347485227e-19

R117_124 V117 V124 -228.6758818173678
L117_124 V117 V124 1.7516014560593108e-12
C117_124 V117 V124 4.66637842300442e-19

R117_125 V117 V125 122.33326027963334
L117_125 V117 V125 1.5145109590513357e-12
C117_125 V117 V125 2.7066367576715807e-19

R117_126 V117 V126 151.53753629027838
L117_126 V117 V126 1.508540625189435e-12
C117_126 V117 V126 1.9919089145849405e-19

R117_127 V117 V127 539.9947727001996
L117_127 V117 V127 -2.507299144336649e-10
C117_127 V117 V127 1.6521937852757033e-20

R117_128 V117 V128 -611.2458732762287
L117_128 V117 V128 -6.000238160789157e-12
C117_128 V117 V128 2.312392615714562e-20

R117_129 V117 V129 -87.29074381262572
L117_129 V117 V129 2.6922387340828857e-12
C117_129 V117 V129 2.2703616751117484e-19

R117_130 V117 V130 -135.53119013748534
L117_130 V117 V130 -1.211183424605581e-12
C117_130 V117 V130 -3.484273516103082e-19

R117_131 V117 V131 -428.8089209051522
L117_131 V117 V131 -3.74778889025388e-12
C117_131 V117 V131 -1.8011625748568606e-19

R117_132 V117 V132 613.1369732959795
L117_132 V117 V132 -2.066207276526868e-12
C117_132 V117 V132 -4.354170292288384e-19

R117_133 V117 V133 -635.3129612803676
L117_133 V117 V133 -1.475766710932847e-12
C117_133 V117 V133 -3.1976722781597865e-19

R117_134 V117 V134 194.45197316950075
L117_134 V117 V134 2.7169244740556383e-12
C117_134 V117 V134 2.0718655308363985e-19

R117_135 V117 V135 511.86376036505
L117_135 V117 V135 1.4401737658498327e-11
C117_135 V117 V135 7.461182732134429e-20

R117_136 V117 V136 -15973.81623712701
L117_136 V117 V136 4.337245186062889e-12
C117_136 V117 V136 2.5073634189115248e-19

R117_137 V117 V137 88.5814842767331
L117_137 V117 V137 -2.7413747576530605e-12
C117_137 V117 V137 -2.8311617338922735e-19

R117_138 V117 V138 2243.2554111157547
L117_138 V117 V138 3.768995877622342e-12
C117_138 V117 V138 2.5392814934881097e-20

R117_139 V117 V139 260.48370898877215
L117_139 V117 V139 -2.2009203753383464e-11
C117_139 V117 V139 -9.555959795133848e-20

R117_140 V117 V140 137.10665879037015
L117_140 V117 V140 2.159422282099739e-11
C117_140 V117 V140 -1.733552836336431e-19

R117_141 V117 V141 -2137.8459705305545
L117_141 V117 V141 1.1124137551098515e-12
C117_141 V117 V141 4.1621356682818066e-19

R117_142 V117 V142 -140.21215735696265
L117_142 V117 V142 -2.1379505216226754e-12
C117_142 V117 V142 -1.0079090673989497e-19

R117_143 V117 V143 -115.27732501900549
L117_143 V117 V143 1.1027323627420935e-11
C117_143 V117 V143 1.110591240193855e-19

R117_144 V117 V144 -96.33852872462256
L117_144 V117 V144 -9.928482897198604e-12
C117_144 V117 V144 8.734968543955741e-20

R117_145 V117 V145 -51.59259034290573
L117_145 V117 V145 1.715709724306761e-11
C117_145 V117 V145 2.7956940941995464e-19

R117_146 V117 V146 -114.59327013494027
L117_146 V117 V146 1.078815332108024e-11
C117_146 V117 V146 -3.58412772925263e-20

R117_147 V117 V147 -312.2716756869933
L117_147 V117 V147 5.524667768156689e-12
C117_147 V117 V147 1.7109636575386736e-19

R117_148 V117 V148 -1000.0906272979644
L117_148 V117 V148 1.9501232053737053e-12
C117_148 V117 V148 2.0346227206051655e-19

R117_149 V117 V149 102.27374301736592
L117_149 V117 V149 -9.781544066793592e-13
C117_149 V117 V149 -6.176731607678222e-19

R117_150 V117 V150 54.94981319134944
L117_150 V117 V150 2.9816374895443643e-12
C117_150 V117 V150 3.5570491344606085e-19

R117_151 V117 V151 78.60578160343283
L117_151 V117 V151 2.766123501446312e-11
C117_151 V117 V151 -1.2338132514001104e-19

R117_152 V117 V152 113.99828176934363
L117_152 V117 V152 -8.236243604625782e-12
C117_152 V117 V152 -5.756052126700215e-20

R117_153 V117 V153 71.49517149354737
L117_153 V117 V153 -1.9602311313180547e-11
C117_153 V117 V153 -7.950269120365234e-20

R117_154 V117 V154 119.90488917574052
L117_154 V117 V154 -1.020324843336408e-11
C117_154 V117 V154 -2.521320811013046e-19

R117_155 V117 V155 -173.20361012600145
L117_155 V117 V155 -1.864874871071498e-12
C117_155 V117 V155 -1.4295632439561967e-19

R117_156 V117 V156 315.62032452689334
L117_156 V117 V156 -1.06173028803769e-11
C117_156 V117 V156 -2.2978555285459997e-19

R117_157 V117 V157 -441.0927274912766
L117_157 V117 V157 1.069810768370292e-12
C117_157 V117 V157 4.982120221625627e-19

R117_158 V117 V158 -63.66131607239683
L117_158 V117 V158 -4.462107132054094e-12
C117_158 V117 V158 2.8510311391483617e-20

R117_159 V117 V159 -158.4015937910424
L117_159 V117 V159 -3.062442125932523e-11
C117_159 V117 V159 -1.1006971036268593e-20

R117_160 V117 V160 -85.2066071265328
L117_160 V117 V160 -3.50001728505018e-12
C117_160 V117 V160 -6.175943228884959e-21

R117_161 V117 V161 -140.1823184781824
L117_161 V117 V161 6.747206772910405e-12
C117_161 V117 V161 5.0006428644445967e-20

R117_162 V117 V162 -252.91515541133276
L117_162 V117 V162 -3.348492154579905e-12
C117_162 V117 V162 -1.5670993045816453e-19

R117_163 V117 V163 182.96739849809305
L117_163 V117 V163 3.1048397900568163e-12
C117_163 V117 V163 5.004449018492805e-20

R117_164 V117 V164 157.0819235660429
L117_164 V117 V164 3.0427388212519676e-12
C117_164 V117 V164 -3.4466525677464695e-20

R117_165 V117 V165 -314.9528112775114
L117_165 V117 V165 -1.6792882539424747e-12
C117_165 V117 V165 -3.2514894064778776e-19

R117_166 V117 V166 42.27839632888198
L117_166 V117 V166 2.8458542784919822e-12
C117_166 V117 V166 7.508346400257529e-20

R117_167 V117 V167 339.86303196577336
L117_167 V117 V167 4.803358875460764e-12
C117_167 V117 V167 7.081106613807939e-20

R117_168 V117 V168 -2708.137399446352
L117_168 V117 V168 5.754685520595958e-12
C117_168 V117 V168 2.0238214925610777e-19

R117_169 V117 V169 245.113059141401
L117_169 V117 V169 5.740763130598324e-12
C117_169 V117 V169 2.7800302996500846e-19

R117_170 V117 V170 -61.90608505638803
L117_170 V117 V170 -4.430626605945006e-12
C117_170 V117 V170 -2.950413274141595e-20

R117_171 V117 V171 -106.09584413698781
L117_171 V117 V171 -1.8831827475757675e-12
C117_171 V117 V171 -1.1851405695811165e-19

R117_172 V117 V172 -123.98685417418477
L117_172 V117 V172 -6.507215768507953e-12
C117_172 V117 V172 -8.648985633177852e-20

R117_173 V117 V173 -315.189516008218
L117_173 V117 V173 4.5507559312741826e-10
C117_173 V117 V173 -2.076707482872025e-19

R117_174 V117 V174 -91.85254216785474
L117_174 V117 V174 -2.605972661238316e-12
C117_174 V117 V174 7.171000819270684e-20

R117_175 V117 V175 196.9661965738292
L117_175 V117 V175 -2.6011961840484492e-12
C117_175 V117 V175 -2.001735356683374e-19

R117_176 V117 V176 147.0851733198033
L117_176 V117 V176 -1.6582886385789961e-12
C117_176 V117 V176 -2.993629308452336e-19

R117_177 V117 V177 -2944.3501543567736
L117_177 V117 V177 7.882535960164399e-11
C117_177 V117 V177 6.541419434438806e-21

R117_178 V117 V178 71.387218542963
L117_178 V117 V178 1.973906611685081e-12
C117_178 V117 V178 6.50063172633091e-20

R117_179 V117 V179 2232.0850031941836
L117_179 V117 V179 1.340154523035957e-12
C117_179 V117 V179 3.0421238013486166e-19

R117_180 V117 V180 268.9740944443577
L117_180 V117 V180 1.2242833025282069e-12
C117_180 V117 V180 2.842652737430191e-19

R117_181 V117 V181 -661.3156513461518
L117_181 V117 V181 2.524785522309504e-12
C117_181 V117 V181 3.577088042308278e-19

R117_182 V117 V182 -1408.185803725434
L117_182 V117 V182 -1.7278816507361623e-12
C117_182 V117 V182 -1.6670425505304274e-19

R117_183 V117 V183 -461.5734720353584
L117_183 V117 V183 2.7409088038462513e-12
C117_183 V117 V183 9.811187332650257e-20

R117_184 V117 V184 -154.51886745814122
L117_184 V117 V184 3.3291919479977534e-12
C117_184 V117 V184 4.186155313832075e-20

R117_185 V117 V185 584.1150725879576
L117_185 V117 V185 -5.274329419885652e-11
C117_185 V117 V185 -2.6320451952437533e-19

R117_186 V117 V186 -179.01409792434217
L117_186 V117 V186 5.6869574980738405e-12
C117_186 V117 V186 1.2431724571574492e-19

R117_187 V117 V187 1144.1597051517056
L117_187 V117 V187 -1.6680107934514629e-12
C117_187 V117 V187 -2.8628902779341343e-19

R117_188 V117 V188 766.0703391685436
L117_188 V117 V188 -1.0765240560803097e-12
C117_188 V117 V188 -2.1472768709857052e-19

R117_189 V117 V189 177.90785271935368
L117_189 V117 V189 -2.6565037410326876e-12
C117_189 V117 V189 -2.5353583647341067e-19

R117_190 V117 V190 426.11354760882904
L117_190 V117 V190 1.0441938766443967e-11
C117_190 V117 V190 1.353396068612398e-19

R117_191 V117 V191 325.3579149952638
L117_191 V117 V191 -2.2668227058590024e-12
C117_191 V117 V191 -1.3442208718127251e-19

R117_192 V117 V192 227.1321869823274
L117_192 V117 V192 1.0641636360205345e-11
C117_192 V117 V192 -6.176899763141025e-20

R117_193 V117 V193 -200.68652929328087
L117_193 V117 V193 -3.3424040119781626e-11
C117_193 V117 V193 1.9028456515518198e-19

R117_194 V117 V194 4212.812953390001
L117_194 V117 V194 -8.16800870691905e-12
C117_194 V117 V194 8.39135944622605e-20

R117_195 V117 V195 -479.15186806628003
L117_195 V117 V195 1.1545193872448288e-12
C117_195 V117 V195 3.4329714695274053e-19

R117_196 V117 V196 -602.2697772610214
L117_196 V117 V196 2.495729103191215e-12
C117_196 V117 V196 1.211493175724259e-19

R117_197 V117 V197 -302.5161635058547
L117_197 V117 V197 1.3682193680523247e-12
C117_197 V117 V197 2.5134806741133884e-19

R117_198 V117 V198 494.4238656226361
L117_198 V117 V198 1.250342754125611e-09
C117_198 V117 V198 -5.200913805694407e-21

R117_199 V117 V199 2919.657112109281
L117_199 V117 V199 4.5971996194428395e-12
C117_199 V117 V199 6.569637284125332e-20

R117_200 V117 V200 -204.57637672331606
L117_200 V117 V200 3.765528670057607e-12
C117_200 V117 V200 9.393502385671223e-20

R118_118 V118 0 23.99203492807731
L118_118 V118 0 -4.0431864441041886e-13
C118_118 V118 0 -2.0511284333824578e-18

R118_119 V118 V119 -434.8627501025832
L118_119 V118 V119 6.696174880344536e-12
C118_119 V118 V119 -1.6259750771164168e-19

R118_120 V118 V120 388.35823609008844
L118_120 V118 V120 -1.0987268654672557e-11
C118_120 V118 V120 -4.674117723742965e-19

R118_121 V118 V121 -164.68156364040965
L118_121 V118 V121 -3.091474045157526e-12
C118_121 V118 V121 -8.864699754356275e-20

R118_122 V118 V122 76.03405322244873
L118_122 V118 V122 1.3135656890020055e-12
C118_122 V118 V122 2.634720482544306e-19

R118_123 V118 V123 -318.3420329483613
L118_123 V118 V123 1.595328524837855e-12
C118_123 V118 V123 5.537932409241164e-19

R118_124 V118 V124 -202.92571787215763
L118_124 V118 V124 1.939277464079429e-12
C118_124 V118 V124 6.32857096987706e-19

R118_125 V118 V125 766.8288281959486
L118_125 V118 V125 1.4076570356624368e-11
C118_125 V118 V125 -6.131732189580659e-20

R118_126 V118 V126 24.601380901825934
L118_126 V118 V126 6.237372424324681e-13
C118_126 V118 V126 5.108143297520749e-19

R118_127 V118 V127 67.68855176265026
L118_127 V118 V127 -1.3218796718467347e-11
C118_127 V118 V127 -1.1635012983700165e-19

R118_128 V118 V128 95.07793366052785
L118_128 V118 V128 -9.673969166500231e-12
C118_128 V118 V128 4.041846273303243e-20

R118_129 V118 V129 104.1222948908626
L118_129 V118 V129 1.4435740029651492e-12
C118_129 V118 V129 5.3824852038565845e-19

R118_130 V118 V130 -35.47659499271873
L118_130 V118 V130 -7.509071635682529e-13
C118_130 V118 V130 -4.553615670020298e-19

R118_131 V118 V131 -62.43231072566773
L118_131 V118 V131 -2.3213702555135934e-12
C118_131 V118 V131 -2.665824935795538e-19

R118_132 V118 V132 -60.36334457130039
L118_132 V118 V132 -1.4895699897598698e-12
C118_132 V118 V132 -6.120642458677047e-19

R118_133 V118 V133 -8323.629357787944
L118_133 V118 V133 -1.994268042088834e-12
C118_133 V118 V133 -4.1041565300849443e-19

R118_134 V118 V134 -71.10150991861806
L118_134 V118 V134 8.107266720962155e-12
C118_134 V118 V134 2.232144713297513e-20

R118_135 V118 V135 -104.33932369262295
L118_135 V118 V135 7.370629528721617e-12
C118_135 V118 V135 4.607868898250223e-19

R118_136 V118 V136 -58.77686057890217
L118_136 V118 V136 1.2217842152106129e-11
C118_136 V118 V136 5.364977461408145e-19

R118_137 V118 V137 -94.8754110508394
L118_137 V118 V137 -2.5341305530147907e-12
C118_137 V118 V137 -1.736754612420041e-19

R118_138 V118 V138 39.204425327935226
L118_138 V118 V138 1.4421842878625304e-12
C118_138 V118 V138 2.657431079934646e-19

R118_139 V118 V139 37.5709812631267
L118_139 V118 V139 -3.44792532249134e-12
C118_139 V118 V139 -7.25218457966854e-19

R118_140 V118 V140 24.97013748577904
L118_140 V118 V140 2.1912992204010193e-12
C118_140 V118 V140 -5.043994626129089e-19

R118_141 V118 V141 -111.30173068810296
L118_141 V118 V141 1.256427959490342e-12
C118_141 V118 V141 6.31815102463109e-19

R118_142 V118 V142 79.32816202882442
L118_142 V118 V142 2.0507010274951154e-11
C118_142 V118 V142 -5.639705102206669e-20

R118_143 V118 V143 -88.5097842227741
L118_143 V118 V143 1.893530913497661e-12
C118_143 V118 V143 3.389522984769928e-19

R118_144 V118 V144 -111.37821249102062
L118_144 V118 V144 -1.4195102721596403e-11
C118_144 V118 V144 9.727311489271302e-20

R118_145 V118 V145 76.28915808062094
L118_145 V118 V145 2.5957887459916103e-12
C118_145 V118 V145 1.351033893363598e-19

R118_146 V118 V146 -31.054617965908598
L118_146 V118 V146 -1.4590194105751257e-12
C118_146 V118 V146 -1.6581261423222606e-19

R118_147 V118 V147 -162.6554339128499
L118_147 V118 V147 5.6898746777659906e-11
C118_147 V118 V147 5.55393913765414e-19

R118_148 V118 V148 -63.210116010039606
L118_148 V118 V148 3.1132109496269076e-12
C118_148 V118 V148 4.0383921125785373e-19

R118_149 V118 V149 256.38522005954525
L118_149 V118 V149 -5.347051517267176e-13
C118_149 V118 V149 -1.026098437728513e-18

R118_150 V118 V150 -38.86319251671797
L118_150 V118 V150 -1.1344308298136127e-11
C118_150 V118 V150 4.2916468813275456e-19

R118_151 V118 V151 168.70320203072
L118_151 V118 V151 -4.103209679802029e-12
C118_151 V118 V151 -3.752062339531253e-19

R118_152 V118 V152 58.168442195870966
L118_152 V118 V152 -7.073515399020481e-12
C118_152 V118 V152 -8.44350933509164e-20

R118_153 V118 V153 -181.07465940147733
L118_153 V118 V153 9.099893270382856e-12
C118_153 V118 V153 1.0607516841549106e-19

R118_154 V118 V154 31.974300770100104
L118_154 V118 V154 1.8250671021945788e-12
C118_154 V118 V154 -2.0602612944990197e-19

R118_155 V118 V155 82.69745801506967
L118_155 V118 V155 -1.1771543830102424e-12
C118_155 V118 V155 -4.630133797729309e-19

R118_156 V118 V156 -133.03250626018638
L118_156 V118 V156 -4.7558858492293454e-11
C118_156 V118 V156 -3.483727020527029e-19

R118_157 V118 V157 -142.12313114741121
L118_157 V118 V157 5.511027773742628e-13
C118_157 V118 V157 1.0092225072839882e-18

R118_158 V118 V158 -541.9853257766207
L118_158 V118 V158 -3.3758878343974406e-12
C118_158 V118 V158 -9.837158083356964e-20

R118_159 V118 V159 -45.69816008651433
L118_159 V118 V159 2.290773187977185e-12
C118_159 V118 V159 3.2587632540819733e-19

R118_160 V118 V160 -75.18252175583622
L118_160 V118 V160 -7.801187985000974e-12
C118_160 V118 V160 1.0453182440713491e-19

R118_161 V118 V161 60.89788884433703
L118_161 V118 V161 -3.66780669666035e-12
C118_161 V118 V161 -2.655151796347062e-19

R118_162 V118 V162 -148.05066349634896
L118_162 V118 V162 -1.4964625621443935e-12
C118_162 V118 V162 -1.088306086684895e-19

R118_163 V118 V163 65.6994859610821
L118_163 V118 V163 1.829932975907584e-12
C118_163 V118 V163 5.0065479595042945e-20

R118_164 V118 V164 56.31211421511232
L118_164 V118 V164 2.343086223621721e-12
C118_164 V118 V164 -1.2521695230457558e-19

R118_165 V118 V165 -150.37943203141668
L118_165 V118 V165 -1.2243978592974427e-12
C118_165 V118 V165 -3.3050706688680986e-19

R118_166 V118 V166 -137.26568224330597
L118_166 V118 V166 3.668286224366562e-12
C118_166 V118 V166 1.732112922239646e-19

R118_167 V118 V167 710.096257957403
L118_167 V118 V167 -5.216386919386961e-12
C118_167 V118 V167 -1.2436046870320893e-19

R118_168 V118 V168 147.6141909135144
L118_168 V118 V168 -2.9314191434169497e-12
C118_168 V118 V168 7.437333551744545e-21

R118_169 V118 V169 -44.74506560232859
L118_169 V118 V169 4.8102656512732e-12
C118_169 V118 V169 4.046230795372397e-19

R118_170 V118 V170 -810.9296310803448
L118_170 V118 V170 -1.645767526315247e-11
C118_170 V118 V170 -2.795743401147237e-19

R118_171 V118 V171 -74.17031180579079
L118_171 V118 V171 -1.1307854351872596e-12
C118_171 V118 V171 -1.6832176674382886e-19

R118_172 V118 V172 -61.76743627571806
L118_172 V118 V172 -6.375328878323846e-12
C118_172 V118 V172 -4.835213866619812e-20

R118_173 V118 V173 56.600088099326015
L118_173 V118 V173 4.0549483439954354e-12
C118_173 V118 V173 -3.3815795335037425e-20

R118_174 V118 V174 159.92708723772154
L118_174 V118 V174 8.024393684333955e-12
C118_174 V118 V174 2.7486856186993165e-19

R118_175 V118 V175 28441.85871086849
L118_175 V118 V175 5.82758235154158e-11
C118_175 V118 V175 -2.269457267004002e-19

R118_176 V118 V176 222.03724787543538
L118_176 V118 V176 2.6915116530724798e-11
C118_176 V118 V176 -1.9636427923169285e-19

R118_177 V118 V177 152.74845519489614
L118_177 V118 V177 2.8337685696114934e-12
C118_177 V118 V177 -7.046062964065989e-20

R118_178 V118 V178 395.13929526121893
L118_178 V118 V178 6.928348078959887e-12
C118_178 V118 V178 1.67699522510557e-19

R118_179 V118 V179 99.1939760820785
L118_179 V118 V179 1.0443180135345992e-12
C118_179 V118 V179 5.323121573516701e-19

R118_180 V118 V180 94.99875127503476
L118_180 V118 V180 1.1727399950358148e-12
C118_180 V118 V180 4.227994402078547e-19

R118_181 V118 V181 -69.69281086185848
L118_181 V118 V181 -2.5737498102707276e-12
C118_181 V118 V181 4.361744535020006e-21

R118_182 V118 V182 -60.43911787594817
L118_182 V118 V182 -1.1553433953966253e-12
C118_182 V118 V182 -2.739720327744498e-19

R118_183 V118 V183 -254.69445373345405
L118_183 V118 V183 2.0461048349513013e-12
C118_183 V118 V183 9.164627332909957e-20

R118_184 V118 V184 -184.42428856232405
L118_184 V118 V184 6.107354990604395e-12
C118_184 V118 V184 -3.9259019288965153e-20

R118_185 V118 V185 779.2999198044566
L118_185 V118 V185 -3.8357150588738455e-12
C118_185 V118 V185 2.4604009121026015e-21

R118_186 V118 V186 -231.15250127499826
L118_186 V118 V186 4.9000542856372385e-12
C118_186 V118 V186 3.7240173877239566e-20

R118_187 V118 V187 -4401.384447817808
L118_187 V118 V187 -9.833296014458788e-13
C118_187 V118 V187 -5.560757306237457e-19

R118_188 V118 V188 328.24234342946346
L118_188 V118 V188 -7.630198280930168e-13
C118_188 V118 V188 -3.9260188639697686e-19

R118_189 V118 V189 167.45613365737103
L118_189 V118 V189 3.981956693396293e-12
C118_189 V118 V189 -5.448845475900356e-20

R118_190 V118 V190 216.16416067082105
L118_190 V118 V190 5.6837873653735754e-12
C118_190 V118 V190 2.1355694632158127e-19

R118_191 V118 V191 603.671488897229
L118_191 V118 V191 -1.548238082312097e-12
C118_191 V118 V191 9.68063915057573e-21

R118_192 V118 V192 224.6152063407979
L118_192 V118 V192 4.254528760347018e-12
C118_192 V118 V192 1.4885114551790647e-19

R118_193 V118 V193 582.9542216825594
L118_193 V118 V193 4.658421757927821e-12
C118_193 V118 V193 1.700157824585811e-19

R118_194 V118 V194 -204.82976678315032
L118_194 V118 V194 2.372505815373224e-12
C118_194 V118 V194 3.532947333677039e-19

R118_195 V118 V195 -377.7193141636257
L118_195 V118 V195 9.492713760594082e-13
C118_195 V118 V195 2.2160622117572517e-19

R118_196 V118 V196 -163.94074476601878
L118_196 V118 V196 1.2611018606133226e-12
C118_196 V118 V196 9.9279298145681e-20

R118_197 V118 V197 -1250.684527651365
L118_197 V118 V197 4.144230870431852e-12
C118_197 V118 V197 -1.8159842754239532e-20

R118_198 V118 V198 -110.41060469811937
L118_198 V118 V198 -5.4230919093041045e-12
C118_198 V118 V198 -5.998740230201884e-20

R118_199 V118 V199 -265.7291359998227
L118_199 V118 V199 3.5619893926653757e-12
C118_199 V118 V199 1.0507788518217023e-19

R118_200 V118 V200 179.61508475492155
L118_200 V118 V200 2.729977748202559e-11
C118_200 V118 V200 -6.237585487220082e-20

R119_119 V119 0 134.59781974527624
L119_119 V119 0 -2.678218216055853e-12
C119_119 V119 0 -5.706269024773246e-19

R119_120 V119 V120 4415.07852299903
L119_120 V119 V120 -2.4559634139757828e-11
C119_120 V119 V120 -2.875068449239369e-19

R119_121 V119 V121 195.64009480159163
L119_121 V119 V121 9.775174408019087e-12
C119_121 V119 V121 -6.000919277050829e-20

R119_122 V119 V122 528.7367393790648
L119_122 V119 V122 -1.0436594507191098e-11
C119_122 V119 V122 -1.0057244682095396e-19

R119_123 V119 V123 48.88179301232105
L119_123 V119 V123 1.43449263355825e-12
C119_123 V119 V123 1.7179266501854357e-19

R119_124 V119 V124 -2269.970881461351
L119_124 V119 V124 1.8735188867272356e-12
C119_124 V119 V124 5.552521701760723e-19

R119_125 V119 V125 -707.5074756340431
L119_125 V119 V125 -1.1785454769901514e-11
C119_125 V119 V125 -6.512340041637363e-20

R119_126 V119 V126 381.2803674425721
L119_126 V119 V126 -1.613506127466463e-10
C119_126 V119 V126 1.0900169222533499e-19

R119_127 V119 V127 39.12016038514459
L119_127 V119 V127 9.648486678622816e-13
C119_127 V119 V127 1.062160055025047e-19

R119_128 V119 V128 205.02045266644095
L119_128 V119 V128 -3.871726533625571e-12
C119_128 V119 V128 -1.30505279419626e-19

R119_129 V119 V129 -11197.235107046608
L119_129 V119 V129 -9.937836081202842e-12
C119_129 V119 V129 8.241059532243871e-20

R119_130 V119 V130 -411.55175544620266
L119_130 V119 V130 5.3683367023376286e-11
C119_130 V119 V130 -1.1978296383862723e-20

R119_131 V119 V131 -29.8334769180011
L119_131 V119 V131 -1.0824120003143892e-12
C119_131 V119 V131 -3.925298078986988e-20

R119_132 V119 V132 -83.3898269755207
L119_132 V119 V132 -3.3344080184820658e-12
C119_132 V119 V132 -2.307532914834622e-19

R119_133 V119 V133 -525.7189740820044
L119_133 V119 V133 1.7183669452761933e-11
C119_133 V119 V133 1.3601788946993482e-20

R119_134 V119 V134 -130.6880301645049
L119_134 V119 V134 -3.1443342299758486e-12
C119_134 V119 V134 -2.1421654098508852e-19

R119_135 V119 V135 103.45921480320897
L119_135 V119 V135 7.888605527236808e-12
C119_135 V119 V135 -6.220101700890956e-20

R119_136 V119 V136 -118.62201780791248
L119_136 V119 V136 3.5315478623221976e-12
C119_136 V119 V136 4.606646010871135e-19

R119_137 V119 V137 -2105.7393477489727
L119_137 V119 V137 3.806164557297926e-12
C119_137 V119 V137 1.0552185713170285e-19

R119_138 V119 V138 102.06363402892713
L119_138 V119 V138 2.5541794945280828e-12
C119_138 V119 V138 2.2850695064284654e-19

R119_139 V119 V139 -509.86792816506886
L119_139 V119 V139 -1.2950077160968968e-11
C119_139 V119 V139 -5.75144813265305e-20

R119_140 V119 V140 56.12700498466673
L119_140 V119 V140 -6.866732256906088e-12
C119_140 V119 V140 -4.853276868943855e-19

R119_141 V119 V141 444.86238016625526
L119_141 V119 V141 -7.506423449167307e-12
C119_141 V119 V141 -9.872782587168938e-20

R119_142 V119 V142 88.95386329920126
L119_142 V119 V142 2.670074519166417e-12
C119_142 V119 V142 1.747745697467488e-20

R119_143 V119 V143 -160.33313242197195
L119_143 V119 V143 -8.598695670561359e-12
C119_143 V119 V143 7.166683029119285e-20

R119_144 V119 V144 -586.3534334328808
L119_144 V119 V144 5.78657249274083e-11
C119_144 V119 V144 2.3714897990921246e-20

R119_145 V119 V145 501.5411862158441
L119_145 V119 V145 -3.7872604267267e-12
C119_145 V119 V145 -1.0240389138650803e-19

R119_146 V119 V146 -51.818562732816694
L119_146 V119 V146 -1.6359368065321346e-12
C119_146 V119 V146 -9.298900081762394e-20

R119_147 V119 V147 59.21241020081025
L119_147 V119 V147 2.5440818194825785e-12
C119_147 V119 V147 5.035960931125083e-20

R119_148 V119 V148 -102.70888092652905
L119_148 V119 V148 5.4546706288172424e-12
C119_148 V119 V148 3.1206115669291415e-19

R119_149 V119 V149 -180.08414767594456
L119_149 V119 V149 3.0558536697587052e-12
C119_149 V119 V149 7.805083002196316e-20

R119_150 V119 V150 -109.09463421205253
L119_150 V119 V150 -1.1063790827377225e-11
C119_150 V119 V150 -4.061548299431677e-20

R119_151 V119 V151 -6294.20541852833
L119_151 V119 V151 1.4346256001109612e-11
C119_151 V119 V151 -2.944993844942299e-20

R119_152 V119 V152 189.3026037184486
L119_152 V119 V152 -3.704028568603184e-12
C119_152 V119 V152 -1.1247262078681289e-19

R119_153 V119 V153 -335.96121747968965
L119_153 V119 V153 -1.8418986854223753e-11
C119_153 V119 V153 1.416743975376429e-19

R119_154 V119 V154 76.46320351782144
L119_154 V119 V154 5.018374312532243e-12
C119_154 V119 V154 1.4052683519375398e-19

R119_155 V119 V155 -181.0048133715767
L119_155 V119 V155 -4.716397892704256e-12
C119_155 V119 V155 7.047841524878703e-21

R119_156 V119 V156 3438.9294168025654
L119_156 V119 V156 6.36207014319283e-12
C119_156 V119 V156 -1.7699684733697155e-19

R119_157 V119 V157 110.92331530007561
L119_157 V119 V157 1.9430369066265375e-11
C119_157 V119 V157 6.921311778853726e-20

R119_158 V119 V158 1819.5238397364355
L119_158 V119 V158 4.962726689218338e-12
C119_158 V119 V158 -4.2912983909817486e-20

R119_159 V119 V159 -170.6446395681789
L119_159 V119 V159 -2.6274458106613194e-12
C119_159 V119 V159 -1.4381338469311335e-20

R119_160 V119 V160 -457.70513188655923
L119_160 V119 V160 4.1116218445561e-12
C119_160 V119 V160 1.9394668498618665e-19

R119_161 V119 V161 339.7809446512448
L119_161 V119 V161 -4.882345588491903e-12
C119_161 V119 V161 -2.3971725396928337e-19

R119_162 V119 V162 -149.2252217778271
L119_162 V119 V162 -7.586662415002417e-12
C119_162 V119 V162 -2.5402959963466533e-20

R119_163 V119 V163 345.48310632588755
L119_163 V119 V163 2.4682880376309016e-12
C119_163 V119 V163 6.882186415068624e-20

R119_164 V119 V164 1366.2209053741544
L119_164 V119 V164 -6.548554933983512e-12
C119_164 V119 V164 -1.3815068350677415e-19

R119_165 V119 V165 -112.57162485310903
L119_165 V119 V165 6.525092591177488e-12
C119_165 V119 V165 9.07144717316148e-20

R119_166 V119 V166 1325.4702721200472
L119_166 V119 V166 2.939153345312839e-11
C119_166 V119 V166 3.548842465560423e-20

R119_167 V119 V167 -141.5658916540471
L119_167 V119 V167 -3.251232369533188e-12
C119_167 V119 V167 -1.3568191150264582e-19

R119_168 V119 V168 923.6922611904465
L119_168 V119 V168 -5.580521525872694e-12
C119_168 V119 V168 -1.1356249932765827e-19

R119_169 V119 V169 -207.2021609042837
L119_169 V119 V169 -2.0091803615670468e-11
C119_169 V119 V169 2.420652784403991e-19

R119_170 V119 V170 -549.8189603181424
L119_170 V119 V170 -1.487338698672592e-11
C119_170 V119 V170 3.027684124788692e-21

R119_171 V119 V171 69.27606768873129
L119_171 V119 V171 2.5997625308468834e-12
C119_171 V119 V171 1.1491674960876192e-19

R119_172 V119 V172 -521.2759997065469
L119_172 V119 V172 2.7947037224629574e-12
C119_172 V119 V172 1.4574862506148721e-19

R119_173 V119 V173 87.63077561947044
L119_173 V119 V173 2.961413516224812e-11
C119_173 V119 V173 -9.438088493864332e-20

R119_174 V119 V174 -3872.850023603735
L119_174 V119 V174 9.454396615659557e-12
C119_174 V119 V174 9.702388970049107e-20

R119_175 V119 V175 -155.8185138201455
L119_175 V119 V175 2.6077401383539687e-12
C119_175 V119 V175 6.6141464590914514e-21

R119_176 V119 V176 366.7895090174251
L119_176 V119 V176 -6.259753839193353e-12
C119_176 V119 V176 -1.4493420086873092e-19

R119_177 V119 V177 -331.6275290026896
L119_177 V119 V177 3.7447830630692716e-11
C119_177 V119 V177 -2.575294649430618e-20

R119_178 V119 V178 161.25201625532188
L119_178 V119 V178 9.650277084732784e-12
C119_178 V119 V178 -3.649136403161618e-20

R119_179 V119 V179 -64.95630963661218
L119_179 V119 V179 -1.269534379433346e-12
C119_179 V119 V179 -7.587832356138793e-21

R119_180 V119 V180 337.06283978348523
L119_180 V119 V180 7.602209905946987e-11
C119_180 V119 V180 1.120569117370074e-19

R119_181 V119 V181 -235.15714193990857
L119_181 V119 V181 -2.0566126308380632e-11
C119_181 V119 V181 -9.95323645009249e-20

R119_182 V119 V182 -196.37542094157067
L119_182 V119 V182 1.8236823425660724e-09
C119_182 V119 V182 1.606404655134829e-20

R119_183 V119 V183 63.638820580193396
L119_183 V119 V183 3.077472397213478e-12
C119_183 V119 V183 3.6973475416565174e-20

R119_184 V119 V184 -283.48429965746595
L119_184 V119 V184 6.375326647367323e-11
C119_184 V119 V184 -4.821818177352955e-20

R119_185 V119 V185 226.97334721597107
L119_185 V119 V185 -1.5449422730720847e-11
C119_185 V119 V185 7.023934871428001e-20

R119_186 V119 V186 -188.92698755755853
L119_186 V119 V186 1.4208824831352386e-10
C119_186 V119 V186 -4.087533206071999e-20

R119_187 V119 V187 283.1010992273317
L119_187 V119 V187 2.6099851801830773e-12
C119_187 V119 V187 -9.231273688979807e-20

R119_188 V119 V188 482.97941566356644
L119_188 V119 V188 -3.288584347034212e-12
C119_188 V119 V188 -1.0964355932923192e-19

R119_189 V119 V189 -599.4187269315188
L119_189 V119 V189 8.813055218394918e-12
C119_189 V119 V189 1.2008626089968079e-19

R119_190 V119 V190 335.37671958213735
L119_190 V119 V190 -1.1850918974090353e-10
C119_190 V119 V190 -1.9056162050416785e-20

R119_191 V119 V191 -79.15485454846606
L119_191 V119 V191 -4.319072667934736e-12
C119_191 V119 V191 5.686252212063088e-20

R119_192 V119 V192 583.4324691831679
L119_192 V119 V192 2.0163087033194e-12
C119_192 V119 V192 2.816895841696022e-19

R119_193 V119 V193 -631.3704498618783
L119_193 V119 V193 1.3616340256311678e-11
C119_193 V119 V193 2.5651599786632496e-20

R119_194 V119 V194 -1285.6181072434276
L119_194 V119 V194 5.176661267861481e-12
C119_194 V119 V194 2.7326674510943653e-19

R119_195 V119 V195 99.56699419728173
L119_195 V119 V195 4.244197430138111e-12
C119_195 V119 V195 2.2858654413902144e-20

R119_196 V119 V196 -237.61551463738033
L119_196 V119 V196 -1.5870387637111673e-12
C119_196 V119 V196 -4.0023846686075285e-19

R119_197 V119 V197 304.2610935254141
L119_197 V119 V197 -1.1882060165764155e-11
C119_197 V119 V197 -1.7588966803522063e-19

R119_198 V119 V198 -252.79241695786487
L119_198 V119 V198 -6.706513381912201e-11
C119_198 V119 V198 -9.898389018336826e-22

R119_199 V119 V199 439.9642932037876
L119_199 V119 V199 -1.3889266387488832e-11
C119_199 V119 V199 1.1355878636646155e-20

R119_200 V119 V200 264.24926070280094
L119_200 V119 V200 9.45568278630026e-12
C119_200 V119 V200 -1.9317845717687898e-20

R120_120 V120 0 -287.98501970209173
L120_120 V120 0 -8.026206915843401e-13
C120_120 V120 0 -2.0924330270315952e-18

R120_121 V120 V121 251.21239118080425
L120_121 V120 V121 -1.0284287773292869e-11
C120_121 V120 V121 -8.721710276190118e-20

R120_122 V120 V122 -417.171977473045
L120_122 V120 V122 -1.0507516112665835e-11
C120_122 V120 V122 -5.964948093889584e-20

R120_123 V120 V123 -401.1537773200347
L120_123 V120 V123 5.01516073921291e-12
C120_123 V120 V123 2.6739587690040426e-19

R120_124 V120 V124 44.611967687013795
L120_124 V120 V124 5.875516126771628e-13
C120_124 V120 V124 1.2107511000249364e-18

R120_125 V120 V125 -169.92079308830492
L120_125 V120 V125 -5.688597595022996e-12
C120_125 V120 V125 -4.8980407553404233e-20

R120_126 V120 V126 -284.50125106636915
L120_126 V120 V126 4.2654032153217875e-12
C120_126 V120 V126 3.2423482596481934e-19

R120_127 V120 V127 -291.44397994881325
L120_127 V120 V127 -2.5031107770715418e-11
C120_127 V120 V127 2.310276743294197e-19

R120_128 V120 V128 37.141476170885944
L120_128 V120 V128 3.7671297530664355e-12
C120_128 V120 V128 -1.9363503238412746e-19

R120_129 V120 V129 318.57652691288564
L120_129 V120 V129 4.33557424627076e-12
C120_129 V120 V129 2.9931460556108227e-19

R120_130 V120 V130 255.13901872539535
L120_130 V120 V130 -4.891704475927992e-12
C120_130 V120 V130 -2.6071768009343496e-19

R120_131 V120 V131 387.5636387010112
L120_131 V120 V131 -4.896705842909274e-12
C120_131 V120 V131 -4.037436730509492e-19

R120_132 V120 V132 -24.225458611434934
L120_132 V120 V132 -8.984614603792285e-13
C120_132 V120 V132 -4.530843164060774e-19

R120_133 V120 V133 -331.00503946514357
L120_133 V120 V133 -4.001360009520896e-12
C120_133 V120 V133 -2.350379571794706e-19

R120_134 V120 V134 -103.50795050282854
L120_134 V120 V134 -4.8766970768631394e-12
C120_134 V120 V134 -2.136469851065986e-19

R120_135 V120 V135 -218.67769666946896
L120_135 V120 V135 3.799053000144629e-10
C120_135 V120 V135 3.688587884988785e-21

R120_136 V120 V136 160.47737946284133
L120_136 V120 V136 1.3549039904547127e-12
C120_136 V120 V136 8.667642660548259e-19

R120_137 V120 V137 2614.5755612167095
L120_137 V120 V137 4.133064242772495e-12
C120_137 V120 V137 9.112086203017173e-20

R120_138 V120 V138 116.52422883491882
L120_138 V120 V138 1.653012914238265e-12
C120_138 V120 V138 3.813578181332243e-19

R120_139 V120 V139 133.77588853893997
L120_139 V120 V139 8.827460953541063e-12
C120_139 V120 V139 3.3715049142640607e-20

R120_140 V120 V140 178.88240319283878
L120_140 V120 V140 -1.4486514588019628e-12
C120_140 V120 V140 -1.0249917343684466e-18

R120_141 V120 V141 625.910268109867
L120_141 V120 V141 4.6870984711657376e-12
C120_141 V120 V141 2.1837054117376534e-19

R120_142 V120 V142 91.2098267511169
L120_142 V120 V142 8.879048910805515e-12
C120_142 V120 V142 -2.7397404200007207e-20

R120_143 V120 V143 -529.5985372966314
L120_143 V120 V143 6.117680709674099e-12
C120_143 V120 V143 9.475337251714902e-20

R120_144 V120 V144 -130.2208053445389
L120_144 V120 V144 7.754137908219354e-12
C120_144 V120 V144 1.8697045453816622e-19

R120_145 V120 V145 1027.7176781841738
L120_145 V120 V145 -5.090681011816913e-12
C120_145 V120 V145 -6.911744572783209e-20

R120_146 V120 V146 -51.89994870792391
L120_146 V120 V146 -2.1474297391087998e-12
C120_146 V120 V146 -1.5098516594759297e-19

R120_147 V120 V147 -364.8131679899939
L120_147 V120 V147 1.0091359768976576e-10
C120_147 V120 V147 1.8916026441790188e-19

R120_148 V120 V148 62.28748831033579
L120_148 V120 V148 1.0686889423586062e-12
C120_148 V120 V148 5.619692683140166e-19

R120_149 V120 V149 -192.61457928145816
L120_149 V120 V149 -2.6420803041923244e-12
C120_149 V120 V149 -3.739324723936707e-19

R120_150 V120 V150 -161.36744906026044
L120_150 V120 V150 3.6687845046053725e-10
C120_150 V120 V150 1.814134011033379e-19

R120_151 V120 V151 511.3827138050111
L120_151 V120 V151 -5.031232297566539e-12
C120_151 V120 V151 -1.5234049995083254e-19

R120_152 V120 V152 206.56394300699478
L120_152 V120 V152 -3.3817586576203072e-12
C120_152 V120 V152 -1.6590349900050904e-19

R120_153 V120 V153 -1867.1698191822638
L120_153 V120 V153 -1.2811923179130834e-10
C120_153 V120 V153 1.44747771015473e-19

R120_154 V120 V154 78.9746414828208
L120_154 V120 V154 8.696886417756426e-12
C120_154 V120 V154 3.335514152381638e-20

R120_155 V120 V155 152.9905340787993
L120_155 V120 V155 -5.870576554971898e-12
C120_155 V120 V155 -1.0525477245390972e-19

R120_156 V120 V156 -74.67505506257312
L120_156 V120 V156 -2.517295327304491e-12
C120_156 V120 V156 -4.786318350511303e-19

R120_157 V120 V157 99.47452855391492
L120_157 V120 V157 1.5104974405736356e-12
C120_157 V120 V157 5.75861053424286e-19

R120_158 V120 V158 328.1338953921208
L120_158 V120 V158 5.232954742510529e-12
C120_158 V120 V158 -6.956994448877979e-20

R120_159 V120 V159 -190.00442364703815
L120_159 V120 V159 5.49693279532081e-12
C120_159 V120 V159 8.666099507094223e-20

R120_160 V120 V160 -133.98953714313305
L120_160 V120 V160 -5.658573418052143e-12
C120_160 V120 V160 2.8239460239823557e-19

R120_161 V120 V161 264.6913631796152
L120_161 V120 V161 -3.5482306598078544e-12
C120_161 V120 V161 -3.400341001174249e-19

R120_162 V120 V162 -142.47149869029474
L120_162 V120 V162 -2.63218377872768e-12
C120_162 V120 V162 -9.560934304756338e-20

R120_163 V120 V163 -453.41373560769773
L120_163 V120 V163 -1.4714621917623683e-11
C120_163 V120 V163 7.56508584165644e-20

R120_164 V120 V164 154.1932523659537
L120_164 V120 V164 1.833095305165182e-12
C120_164 V120 V164 -1.9200515309819018e-19

R120_165 V120 V165 -113.12270192770747
L120_165 V120 V165 -5.973468711115061e-12
C120_165 V120 V165 -6.088934969505105e-20

R120_166 V120 V166 -1535.176318998699
L120_166 V120 V166 -2.5906758092545368e-11
C120_166 V120 V166 1.304645643344855e-19

R120_167 V120 V167 248.17412551085062
L120_167 V120 V167 3.3793441017492055e-11
C120_167 V120 V167 -1.538770782790118e-19

R120_168 V120 V168 -170.60809643983683
L120_168 V120 V168 -1.8420319037635666e-12
C120_168 V120 V168 -1.040136100475478e-19

R120_169 V120 V169 -291.663021381793
L120_169 V120 V169 5.074559508435477e-12
C120_169 V120 V169 4.723725823420786e-19

R120_170 V120 V170 669.2289497583614
L120_170 V120 V170 3.24364629981356e-11
C120_170 V120 V170 -1.0916533791864826e-19

R120_171 V120 V171 2057.5496448922263
L120_171 V120 V171 -5.921513174028825e-12
C120_171 V120 V171 -4.362594353517977e-20

R120_172 V120 V172 69.06248158015947
L120_172 V120 V172 1.8930200159673096e-12
C120_172 V120 V172 1.3401420629478541e-19

R120_173 V120 V173 73.2655013413279
L120_173 V120 V173 2.5294798473045123e-11
C120_173 V120 V173 -1.8125260548183154e-19

R120_174 V120 V174 -445.07590307760256
L120_174 V120 V174 1.1641731959956997e-11
C120_174 V120 V174 2.40047798943285e-19

R120_175 V120 V175 -722.8487481398572
L120_175 V120 V175 9.936007632315134e-11
C120_175 V120 V175 1.793801127477256e-20

R120_176 V120 V176 -278.58383323478193
L120_176 V120 V176 3.3700484061674603e-12
C120_176 V120 V176 -3.4772431603171406e-19

R120_177 V120 V177 -416.9591124182737
L120_177 V120 V177 1.0455694838186067e-11
C120_177 V120 V177 -6.336973282446433e-20

R120_178 V120 V178 151.93644829574785
L120_178 V120 V178 4.230187383379824e-12
C120_178 V120 V178 2.0799701989672374e-20

R120_179 V120 V179 148.54723291253995
L120_179 V120 V179 2.338463410451644e-12
C120_179 V120 V179 2.1340252652198316e-19

R120_180 V120 V180 -34.0786546349378
L120_180 V120 V180 -1.4987317852854285e-12
C120_180 V120 V180 3.573152995396892e-19

R120_181 V120 V181 -206.84495339166563
L120_181 V120 V181 -1.0832432384583953e-11
C120_181 V120 V181 -5.186977840255327e-20

R120_182 V120 V182 -605.7756579799221
L120_182 V120 V182 -3.2976019609305592e-12
C120_182 V120 V182 -9.390609487849511e-20

R120_183 V120 V183 -130.07368289719747
L120_183 V120 V183 9.521496291944535e-12
C120_183 V120 V183 1.067723758098481e-19

R120_184 V120 V184 45.25464060075585
L120_184 V120 V184 1.4809579956633445e-12
C120_184 V120 V184 -3.692803383733959e-20

R120_185 V120 V185 142.80357858996726
L120_185 V120 V185 -6.957313241167015e-12
C120_185 V120 V185 7.080212683531543e-20

R120_186 V120 V186 -160.54543405375148
L120_186 V120 V186 2.0029459610227228e-11
C120_186 V120 V186 -2.8258401625900306e-20

R120_187 V120 V187 -311.38544223090554
L120_187 V120 V187 -3.2629697985071127e-12
C120_187 V120 V187 -2.746761463408877e-19

R120_188 V120 V188 76.48463324230512
L120_188 V120 V188 -1.8066844445371083e-12
C120_188 V120 V188 -4.062019804363146e-19

R120_189 V120 V189 -482.20773744429874
L120_189 V120 V189 4.4805311637678194e-12
C120_189 V120 V189 8.41839736266843e-20

R120_190 V120 V190 294.9929655817299
L120_190 V120 V190 2.925664882487377e-11
C120_190 V120 V190 7.945904810074762e-20

R120_191 V120 V191 112.50498552248996
L120_191 V120 V191 -3.6312017986205672e-12
C120_191 V120 V191 -1.0563427384759461e-19

R120_192 V120 V192 -53.84267051931931
L120_192 V120 V192 5.622314436704256e-12
C120_192 V120 V192 4.747284708529732e-19

R120_193 V120 V193 -174.50783446411106
L120_193 V120 V193 1.1686264721102345e-11
C120_193 V120 V193 1.098901389357753e-19

R120_194 V120 V194 8528.165092634097
L120_194 V120 V194 3.1710547029360596e-12
C120_194 V120 V194 4.832730501971635e-19

R120_195 V120 V195 -218.61292165517594
L120_195 V120 V195 2.0916814261487893e-12
C120_195 V120 V195 4.213658508831158e-19

R120_196 V120 V196 95.88675536364477
L120_196 V120 V196 1.4526889056146819e-11
C120_196 V120 V196 -5.904404406476021e-19

R120_197 V120 V197 226.64962526091767
L120_197 V120 V197 -1.9103462763800823e-10
C120_197 V120 V197 -1.9159422971419157e-19

R120_198 V120 V198 -349.2766826725864
L120_198 V120 V198 -4.692957124269867e-11
C120_198 V120 V198 1.9601002563878006e-20

R120_199 V120 V199 -433.0506378196735
L120_199 V120 V199 7.137756574871449e-12
C120_199 V120 V199 3.352811758852515e-20

R120_200 V120 V200 118.448749265581
L120_200 V120 V200 -1.0845938019052867e-11
C120_200 V120 V200 -3.290675505428235e-20

R121_121 V121 0 43.937787848273175
L121_121 V121 0 2.380663050854197e-13
C121_121 V121 0 5.274388537952023e-19

R121_122 V121 V122 231.49407965278408
L121_122 V121 V122 4.2568640939007806e-12
C121_122 V121 V122 1.713543605004454e-19

R121_123 V121 V123 427.79823741740046
L121_123 V121 V123 1.0824649789012481e-11
C121_123 V121 V123 -9.632402014408262e-21

R121_124 V121 V124 294.3613722197445
L121_124 V121 V124 8.80088610478415e-12
C121_124 V121 V124 -2.0686149104467035e-19

R121_125 V121 V125 -178.4790648490026
L121_125 V121 V125 6.8289266900146365e-12
C121_125 V121 V125 5.746424099953544e-20

R121_126 V121 V126 119.55200105057334
L121_126 V121 V126 5.84326675407169e-12
C121_126 V121 V126 -1.2100985522745112e-19

R121_127 V121 V127 1575.7558625888037
L121_127 V121 V127 2.8438418290516693e-11
C121_127 V121 V127 3.3563827691806556e-20

R121_128 V121 V128 826.3143353875834
L121_128 V121 V128 5.930933593706169e-11
C121_128 V121 V128 6.202843181676089e-20

R121_129 V121 V129 37.68347874024031
L121_129 V121 V129 8.055904864999274e-13
C121_129 V121 V129 5.375489593112434e-19

R121_130 V121 V130 -205.17831999294503
L121_130 V121 V130 -2.6238907545369916e-12
C121_130 V121 V130 -6.240568493343471e-20

R121_131 V121 V131 -347.1555305802897
L121_131 V121 V131 -1.1640716414119572e-11
C121_131 V121 V131 2.6267869928088293e-20

R121_132 V121 V132 -190.5145562002929
L121_132 V121 V132 -4.37028088636423e-12
C121_132 V121 V132 1.0374764054711479e-19

R121_133 V121 V133 -1306.1773852661443
L121_133 V121 V133 -6.420353609922354e-12
C121_133 V121 V133 -1.1691724888622184e-19

R121_134 V121 V134 -182.36325952694816
L121_134 V121 V134 1.7707146728960648e-12
C121_134 V121 V134 3.71975695315285e-19

R121_135 V121 V135 -128.29157765401536
L121_135 V121 V135 -5.454148857827207e-12
C121_135 V121 V135 -7.982693487366558e-20

R121_136 V121 V136 -144.5461588403588
L121_136 V121 V136 -7.324743150606005e-11
C121_136 V121 V136 -9.28968417945158e-20

R121_137 V121 V137 -41.39565073979019
L121_137 V121 V137 -6.5965878670766646e-12
C121_137 V121 V137 3.41393534503683e-20

R121_138 V121 V138 270.8978548003579
L121_138 V121 V138 -3.660197168569405e-12
C121_138 V121 V138 -2.8520892444581264e-19

R121_139 V121 V139 104.04828499872782
L121_139 V121 V139 4.071359891229254e-11
C121_139 V121 V139 9.860036276369877e-21

R121_140 V121 V140 111.48274102042782
L121_140 V121 V140 5.615610637868259e-12
C121_140 V121 V140 1.997399832435072e-19

R121_141 V121 V141 -302.0538204477498
L121_141 V121 V141 -3.647422324879239e-12
C121_141 V121 V141 -1.0435399336685502e-19

R121_142 V121 V142 115.74898217959422
L121_142 V121 V142 -2.0748228202013272e-12
C121_142 V121 V142 -1.3589164038417536e-19

R121_143 V121 V143 125.82529610970526
L121_143 V121 V143 1.738961083738128e-12
C121_143 V121 V143 1.6862215511681814e-19

R121_144 V121 V144 107.37580210818716
L121_144 V121 V144 6.950962634602816e-12
C121_144 V121 V144 -1.0641884452454512e-19

R121_145 V121 V145 33.24142225941899
L121_145 V121 V145 -4.756742311393547e-12
C121_145 V121 V145 -1.830703546093829e-19

R121_146 V121 V146 95.17620751354065
L121_146 V121 V146 1.2829049199381116e-12
C121_146 V121 V146 2.004837575418037e-19

R121_147 V121 V147 -373.7371944666227
L121_147 V121 V147 -2.6827362831370494e-12
C121_147 V121 V147 -2.336979509157413e-19

R121_148 V121 V148 -186.5776193211169
L121_148 V121 V148 -5.095828220196982e-12
C121_148 V121 V148 -2.0605006514384036e-19

R121_149 V121 V149 438.31308484403587
L121_149 V121 V149 -2.0313636562941898e-12
C121_149 V121 V149 -2.483908471967547e-19

R121_150 V121 V150 -35.14403047825555
L121_150 V121 V150 -2.892462438511351e-12
C121_150 V121 V150 8.252353029483033e-20

R121_151 V121 V151 -60.91301645820915
L121_151 V121 V151 -1.4420191190562897e-12
C121_151 V121 V151 -1.3527001166259562e-19

R121_152 V121 V152 -210.52843001305718
L121_152 V121 V152 -7.981459965571359e-12
C121_152 V121 V152 1.2052809265304292e-19

R121_153 V121 V153 -37.69667832904565
L121_153 V121 V153 2.658566628042542e-12
C121_153 V121 V153 4.655686888198639e-19

R121_154 V121 V154 -74.95561564076431
L121_154 V121 V154 -6.020525636218436e-12
C121_154 V121 V154 -1.2145202046313563e-19

R121_155 V121 V155 122.99637256498568
L121_155 V121 V155 8.596235492140192e-12
C121_155 V121 V155 5.132921747825391e-20

R121_156 V121 V156 -91.51677580320525
L121_156 V121 V156 -1.2697464189160976e-11
C121_156 V121 V156 1.3954384823412775e-19

R121_157 V121 V157 -46.83217170831814
L121_157 V121 V157 1.4314490411347572e-12
C121_157 V121 V157 4.860991278841473e-19

R121_158 V121 V158 48.55838922140286
L121_158 V121 V158 1.2630505808403445e-11
C121_158 V121 V158 7.891525867534082e-20

R121_159 V121 V159 181.80970669446907
L121_159 V121 V159 1.6827125698045746e-12
C121_159 V121 V159 1.037983718191383e-19

R121_160 V121 V160 81.65550016732877
L121_160 V121 V160 2.174701494402369e-12
C121_160 V121 V160 -5.797200451157904e-20

R121_161 V121 V161 45.950285482716254
L121_161 V121 V161 -3.2085768462642995e-12
C121_161 V121 V161 -5.705740295073707e-19

R121_162 V121 V162 53.7607297986633
L121_162 V121 V162 4.4961361634578696e-12
C121_162 V121 V162 1.0746539514818416e-19

R121_163 V121 V163 92.85374328161693
L121_163 V121 V163 1.8640020110545763e-12
C121_163 V121 V163 2.322770691031519e-19

R121_164 V121 V164 77.2207034887411
L121_164 V121 V164 4.654011007978532e-12
C121_164 V121 V164 2.3154698112240266e-20

R121_165 V121 V165 74.98212814997127
L121_165 V121 V165 -9.679460192364418e-13
C121_165 V121 V165 -2.78043286902149e-19

R121_166 V121 V166 -33.43954425930501
L121_166 V121 V166 -1.347505918513658e-12
C121_166 V121 V166 -2.82690630001198e-19

R121_167 V121 V167 -109.39124865061011
L121_167 V121 V167 -1.6940951245180999e-12
C121_167 V121 V167 -2.1049368673180238e-19

R121_168 V121 V168 -409.47007930989247
L121_168 V121 V168 -1.898925929403022e-12
C121_168 V121 V168 -2.0882162897178062e-19

R121_169 V121 V169 -49.04762792411186
L121_169 V121 V169 4.619008160710852e-12
C121_169 V121 V169 3.132743543525045e-19

R121_170 V121 V170 907.0224418009869
L121_170 V121 V170 -5.618344362508622e-10
C121_170 V121 V170 -9.579795497875465e-20

R121_171 V121 V171 -177.61225235971526
L121_171 V121 V171 -1.2643057413850905e-12
C121_171 V121 V171 -3.401425787746488e-19

R121_172 V121 V172 -131.6888953467394
L121_172 V121 V172 -3.2184550759465814e-12
C121_172 V121 V172 -6.07414969953781e-20

R121_173 V121 V173 1116.082253499077
L121_173 V121 V173 1.0885787874837453e-12
C121_173 V121 V173 3.301545162784417e-19

R121_174 V121 V174 47.06967331553235
L121_174 V121 V174 1.0737558616956671e-12
C121_174 V121 V174 5.464548689410421e-19

R121_175 V121 V175 206.39915702404278
L121_175 V121 V175 1.1923649184300061e-12
C121_175 V121 V175 3.3802448702931036e-19

R121_176 V121 V176 267.99803734578944
L121_176 V121 V176 9.487452710284155e-13
C121_176 V121 V176 4.413417316161995e-19

R121_177 V121 V177 124.88839516179557
L121_177 V121 V177 -1.3462376840324243e-12
C121_177 V121 V177 -4.119589305539804e-19

R121_178 V121 V178 -231.24398481721423
L121_178 V121 V178 1.984556463214059e-11
C121_178 V121 V178 -2.6801648215976824e-20

R121_179 V121 V179 152.00345971700867
L121_179 V121 V179 2.2412995947247505e-12
C121_179 V121 V179 1.7447097714837397e-19

R121_180 V121 V180 172.33010336031387
L121_180 V121 V180 1.3161872904761105e-11
C121_180 V121 V180 -7.599596933042012e-20

R121_181 V121 V181 -321.9094831810569
L121_181 V121 V181 3.0826420494446595e-12
C121_181 V121 V181 -2.756650357545385e-19

R121_182 V121 V182 -64.64586400305323
L121_182 V121 V182 -1.0858488482542551e-12
C121_182 V121 V182 -2.1638928533376169e-19

R121_183 V121 V183 -144.9539211111082
L121_183 V121 V183 -8.915286869757188e-12
C121_183 V121 V183 2.497009509508789e-20

R121_184 V121 V184 -244.90619246319233
L121_184 V121 V184 -2.3525380519252593e-12
C121_184 V121 V184 -3.986709421607072e-20

R121_185 V121 V185 -130.86386278368693
L121_185 V121 V185 -1.0530285845407705e-11
C121_185 V121 V185 4.482686815030285e-19

R121_186 V121 V186 477.479920887969
L121_186 V121 V186 -1.3106169141926252e-12
C121_186 V121 V186 -2.3046355740133415e-19

R121_187 V121 V187 522.9462534095362
L121_187 V121 V187 -1.3949006110089173e-12
C121_187 V121 V187 -2.1339465559146727e-19

R121_188 V121 V188 -12403.319016906866
L121_188 V121 V188 -1.4514426435083237e-12
C121_188 V121 V188 -2.588107073268545e-19

R121_189 V121 V189 256.30215823442273
L121_189 V121 V189 -9.410329350763716e-12
C121_189 V121 V189 -1.704318860396782e-19

R121_190 V121 V190 112.04500942566776
L121_190 V121 V190 1.441457173452031e-12
C121_190 V121 V190 1.8353981522783813e-19

R121_191 V121 V191 316.370407587649
L121_191 V121 V191 -1.0429422213585617e-11
C121_191 V121 V191 -2.5064473443698397e-19

R121_192 V121 V192 241.5488702793144
L121_192 V121 V192 2.0951622579935974e-12
C121_192 V121 V192 -1.4459564365356703e-21

R121_193 V121 V193 127.16742748885281
L121_193 V121 V193 1.6788159769027188e-12
C121_193 V121 V193 2.1574586138682691e-19

R121_194 V121 V194 -132.07127341941074
L121_194 V121 V194 1.7302059456275148e-12
C121_194 V121 V194 2.9789586386144403e-19

R121_195 V121 V195 -206.24101481140335
L121_195 V121 V195 1.618985705673058e-12
C121_195 V121 V195 3.6496925550282257e-19

R121_196 V121 V196 -199.15560489458449
L121_196 V121 V196 1.0827487868689261e-12
C121_196 V121 V196 5.005600176862948e-19

R121_197 V121 V197 -147.43618159609616
L121_197 V121 V197 -5.4548189272755934e-12
C121_197 V121 V197 -2.1917244539265016e-19

R121_198 V121 V198 -96.08876311100967
L121_198 V121 V198 -1.6408896504031812e-12
C121_198 V121 V198 -1.0583075970319996e-19

R121_199 V121 V199 -229.32400061406156
L121_199 V121 V199 1.202310747585205e-11
C121_199 V121 V199 2.90459195040128e-19

R121_200 V121 V200 823.1528698659021
L121_200 V121 V200 -1.7507119049606769e-12
C121_200 V121 V200 -1.5476268753852972e-19

R122_122 V122 0 -88.17599684084665
L122_122 V122 0 1.1365242625419064e-12
C122_122 V122 0 1.0277955140941896e-18

R122_123 V122 V123 -429.69868639646904
L122_123 V122 V123 2.935671884174619e-12
C122_123 V122 V123 2.0433835929728863e-19

R122_124 V122 V124 15787.310523006361
L122_124 V122 V124 1.4013599317475774e-12
C122_124 V122 V124 4.46747167571085e-19

R122_125 V122 V125 -2059.400641257443
L122_125 V122 V125 -7.588208415505053e-12
C122_125 V122 V125 -1.1877473654626571e-19

R122_126 V122 V126 -83.37654944081615
L122_126 V122 V126 -8.334154777060773e-11
C122_126 V122 V126 1.2598660783072813e-19

R122_127 V122 V127 -278.88231073065117
L122_127 V122 V127 -5.002474111467864e-12
C122_127 V122 V127 -5.3570964406342444e-20

R122_128 V122 V128 -879.2996631095962
L122_128 V122 V128 -2.768614728820541e-12
C122_128 V122 V128 -1.993198778592045e-19

R122_129 V122 V129 -175.79179657794478
L122_129 V122 V129 -1.699840330938615e-12
C122_129 V122 V129 -3.283292927594943e-19

R122_130 V122 V130 91.96923055327142
L122_130 V122 V130 9.093127747927858e-13
C122_130 V122 V130 5.432251601991124e-19

R122_131 V122 V131 172.8750941780872
L122_131 V122 V131 -6.04593270658406e-12
C122_131 V122 V131 -1.7004671003662183e-19

R122_132 V122 V132 228.4677634404944
L122_132 V122 V132 -4.235279788756337e-12
C122_132 V122 V132 -1.7045582704832706e-19

R122_133 V122 V133 654.384371030648
L122_133 V122 V133 1.6356398523461421e-12
C122_133 V122 V133 3.375490550831024e-19

R122_134 V122 V134 626.2919581973973
L122_134 V122 V134 -1.304188771157547e-12
C122_134 V122 V134 -6.963893739778709e-19

R122_135 V122 V135 11272.662982329983
L122_135 V122 V135 2.005981446256755e-12
C122_135 V122 V135 2.409968377153716e-19

R122_136 V122 V136 262.47822782165997
L122_136 V122 V136 1.9168204214236924e-12
C122_136 V122 V136 3.0585330066162334e-19

R122_137 V122 V137 259.18061445909825
L122_137 V122 V137 1.8653668169674098e-12
C122_137 V122 V137 3.042953775668557e-19

R122_138 V122 V138 -166.91431278713773
L122_138 V122 V138 6.159378963976597e-12
C122_138 V122 V138 3.1637861731005437e-19

R122_139 V122 V139 -213.43678108682806
L122_139 V122 V139 -3.672742440400413e-12
C122_139 V122 V139 -5.462137352691902e-20

R122_140 V122 V140 -97.36366466160034
L122_140 V122 V140 -2.1589260061321505e-12
C122_140 V122 V140 -2.0510840791413935e-19

R122_141 V122 V141 515.3579061251484
L122_141 V122 V141 -1.2122840841797678e-12
C122_141 V122 V141 -5.578025260796332e-19

R122_142 V122 V142 -2795.399558264719
L122_142 V122 V142 3.642703572016237e-12
C122_142 V122 V142 9.744701620485813e-20

R122_143 V122 V143 324.5423848717341
L122_143 V122 V143 -4.614261122388074e-12
C122_143 V122 V143 -2.330367181660986e-19

R122_144 V122 V144 453.99303663101387
L122_144 V122 V144 7.933335980564779e-11
C122_144 V122 V144 -1.0587457096553517e-19

R122_145 V122 V145 -309.42453450723735
L122_145 V122 V145 -2.16624860795501e-12
C122_145 V122 V145 -2.472744200757664e-19

R122_146 V122 V146 424.46267916517326
L122_146 V122 V146 -2.2067517136774103e-12
C122_146 V122 V146 -3.6490242833064777e-20

R122_147 V122 V147 -2563.2411458584993
L122_147 V122 V147 6.335514528588378e-12
C122_147 V122 V147 1.7714405783150394e-19

R122_148 V122 V148 234.4194280571187
L122_148 V122 V148 5.864223560637429e-12
C122_148 V122 V148 1.6169119756402708e-19

R122_149 V122 V149 -197.85131457361612
L122_149 V122 V149 7.288828898997626e-13
C122_149 V122 V149 8.478932113425723e-19

R122_150 V122 V150 142.27219079063312
L122_150 V122 V150 2.0379670461364457e-12
C122_150 V122 V150 -4.386462931052933e-19

R122_151 V122 V151 -505.1830482492112
L122_151 V122 V151 -9.909392742526407e-12
C122_151 V122 V151 5.104710366267099e-20

R122_152 V122 V152 -284.05391585338066
L122_152 V122 V152 -2.9474604418912077e-12
C122_152 V122 V152 -7.724713024139388e-20

R122_153 V122 V153 257.28423245460914
L122_153 V122 V153 5.458815248749549e-12
C122_153 V122 V153 1.1628702111906108e-19

R122_154 V122 V154 -369.577893606976
L122_154 V122 V154 -8.497943076825412e-12
C122_154 V122 V154 4.1966031302896777e-19

R122_155 V122 V155 1025.941817226096
L122_155 V122 V155 7.662085094032912e-12
C122_155 V122 V155 1.180431210059157e-19

R122_156 V122 V156 606.2398334769267
L122_156 V122 V156 5.062901709538007e-12
C122_156 V122 V156 -2.6893846063137773e-20

R122_157 V122 V157 127.58597001094057
L122_157 V122 V157 -9.527349543489438e-13
C122_157 V122 V157 -7.044025989830864e-19

R122_158 V122 V158 -1487.725626406315
L122_158 V122 V158 -4.675726077529092e-12
C122_158 V122 V158 -1.576802270402983e-19

R122_159 V122 V159 232.39918704020727
L122_159 V122 V159 2.874203511998999e-12
C122_159 V122 V159 9.984477495475212e-20

R122_160 V122 V160 451.42084470922777
L122_160 V122 V160 2.179332044971617e-12
C122_160 V122 V160 2.273666027999001e-19

R122_161 V122 V161 -146.0975812590009
L122_161 V122 V161 -1.982863542124246e-12
C122_161 V122 V161 -2.0195178450519144e-19

R122_162 V122 V162 -152.04325473480282
L122_162 V122 V162 3.035872731352159e-12
C122_162 V122 V162 9.899381141579742e-20

R122_163 V122 V163 -158.6195367602816
L122_163 V122 V163 -1.3893294019690147e-12
C122_163 V122 V163 -2.752351725811411e-19

R122_164 V122 V164 -147.23314363286522
L122_164 V122 V164 -1.8944945059073226e-12
C122_164 V122 V164 -1.7213182857800484e-19

R122_165 V122 V165 -366.1963960293727
L122_165 V122 V165 9.743944865443681e-13
C122_165 V122 V165 5.615653616510262e-19

R122_166 V122 V166 237.3381013470067
L122_166 V122 V166 2.5523099323527624e-12
C122_166 V122 V166 6.698313938361826e-21

R122_167 V122 V167 -703.4491249236494
L122_167 V122 V167 -9.212406569192936e-12
C122_167 V122 V167 -6.740860432380941e-20

R122_168 V122 V168 -451.46115687955563
L122_168 V122 V168 -2.7284223914371575e-12
C122_168 V122 V168 -1.8866686171487766e-19

R122_169 V122 V169 105.41558356625366
L122_169 V122 V169 4.4836857679181395e-12
C122_169 V122 V169 5.071628146005189e-20

R122_170 V122 V170 108.12215731192964
L122_170 V122 V170 -2.530453015732274e-12
C122_170 V122 V170 2.0142219233085172e-19

R122_171 V122 V171 164.69997396875507
L122_171 V122 V171 1.0177668082055194e-12
C122_171 V122 V171 4.516198910446386e-19

R122_172 V122 V172 141.35682077922394
L122_172 V122 V172 1.0514532746534566e-12
C122_172 V122 V172 3.271871851372907e-19

R122_173 V122 V173 -392.21131333027296
L122_173 V122 V173 -1.318993547580777e-12
C122_173 V122 V173 -2.263454251780492e-19

R122_174 V122 V174 -118.25517543664682
L122_174 V122 V174 1.6029744339571932e-11
C122_174 V122 V174 -1.5067986685960197e-19

R122_175 V122 V175 7647.162172159376
L122_175 V122 V175 -1.1957170303410868e-11
C122_175 V122 V175 -4.537879559042051e-20

R122_176 V122 V176 -614.4182924659175
L122_176 V122 V176 -6.127463675471086e-12
C122_176 V122 V176 -9.725345357210665e-20

R122_177 V122 V177 -192.25527928631587
L122_177 V122 V177 6.4955200191612235e-12
C122_177 V122 V177 1.529915396738771e-19

R122_178 V122 V178 -156.25458815013118
L122_178 V122 V178 1.0771442905884978e-11
C122_178 V122 V178 -2.397634098605847e-19

R122_179 V122 V179 -555.1552226772667
L122_179 V122 V179 -1.5809880124878613e-12
C122_179 V122 V179 -2.8859329439645236e-19

R122_180 V122 V180 -186.83638449182206
L122_180 V122 V180 -1.3098587999138613e-12
C122_180 V122 V180 -1.4558953728871697e-19

R122_181 V122 V181 223.56527727790655
L122_181 V122 V181 5.513590143078429e-12
C122_181 V122 V181 -1.6991697747158539e-19

R122_182 V122 V182 81.74209071503579
L122_182 V122 V182 2.2290571406162254e-12
C122_182 V122 V182 2.841100316810017e-19

R122_183 V122 V183 -1024.2744210905446
L122_183 V122 V183 1.064886522190552e-10
C122_183 V122 V183 -6.866540845623124e-20

R122_184 V122 V184 369.2902114815752
L122_184 V122 V184 2.4622702933686077e-12
C122_184 V122 V184 -1.4083554190379825e-20

R122_185 V122 V185 288.6531298415593
L122_185 V122 V185 -4.125587114351588e-12
C122_185 V122 V185 -7.265951675744572e-21

R122_186 V122 V186 467.10057276704765
L122_186 V122 V186 2.6929870008355022e-12
C122_186 V122 V186 8.057713559889379e-20

R122_187 V122 V187 -1044.602667062426
L122_187 V122 V187 2.4088289125626324e-12
C122_187 V122 V187 1.6415034737294418e-19

R122_188 V122 V188 -40898.10991619363
L122_188 V122 V188 3.127567758761643e-11
C122_188 V122 V188 7.944762822980076e-20

R122_189 V122 V189 -208.55631167050205
L122_189 V122 V189 2.8452773890083944e-12
C122_189 V122 V189 3.5646406559357915e-19

R122_190 V122 V190 -126.93153054730361
L122_190 V122 V190 -6.126001521381506e-12
C122_190 V122 V190 -3.1806531353367915e-19

R122_191 V122 V191 901.8215922772617
L122_191 V122 V191 3.1106792567890164e-12
C122_191 V122 V191 3.278389560114673e-19

R122_192 V122 V192 -449.0061889365538
L122_192 V122 V192 3.664548804084631e-12
C122_192 V122 V192 3.9538421904747185e-19

R122_193 V122 V193 -387.4779065451841
L122_193 V122 V193 -1.5488947569429944e-11
C122_193 V122 V193 -1.4539797398517226e-19

R122_194 V122 V194 166.74354531499807
L122_194 V122 V194 -8.066012986318289e-12
C122_194 V122 V194 1.1638442211297882e-19

R122_195 V122 V195 2686.7660634871722
L122_195 V122 V195 -1.900236599915916e-12
C122_195 V122 V195 -4.537636606422727e-19

R122_196 V122 V196 548.3866035692347
L122_196 V122 V196 -1.446967401637986e-12
C122_196 V122 V196 -6.931976575366394e-19

R122_197 V122 V197 257.51128815668676
L122_197 V122 V197 -1.6386089285941424e-12
C122_197 V122 V197 -3.0698045859518995e-19

R122_198 V122 V198 174.17106983897935
L122_198 V122 V198 9.06544720847832e-12
C122_198 V122 V198 1.149353387139843e-19

R122_199 V122 V199 19802.860193315457
L122_199 V122 V199 -2.6534647244452334e-12
C122_199 V122 V199 -2.643548750550339e-19

R122_200 V122 V200 -714.7023931755563
L122_200 V122 V200 -8.42489174171459e-12
C122_200 V122 V200 -1.1482822517778715e-19

R123_123 V123 0 1173.0256810396882
L123_123 V123 0 8.291830157994561e-13
C123_123 V123 0 1.0152372460463267e-18

R123_124 V123 V124 -328.10689692948364
L123_124 V123 V124 -8.007137438383591e-11
C123_124 V123 V124 1.4095874493703688e-19

R123_125 V123 V125 1142.0608061148687
L123_125 V123 V125 -1.4132611495067991e-11
C123_125 V123 V125 7.704485107485742e-20

R123_126 V123 V126 -2896.960899562341
L123_126 V123 V126 -1.0833705745415497e-12
C123_126 V123 V126 -4.404703366557534e-19

R123_127 V123 V127 -75.07685780205459
L123_127 V123 V127 7.841033311034981e-13
C123_127 V123 V127 9.314582760238175e-19

R123_128 V123 V128 1454.333925422716
L123_128 V123 V128 -3.2470357775937963e-12
C123_128 V123 V128 -3.2008316551670136e-19

R123_129 V123 V129 -186.61907667901565
L123_129 V123 V129 -2.7717263173472766e-12
C123_129 V123 V129 -2.872667509263836e-19

R123_130 V123 V130 354.5839319044821
L123_130 V123 V130 3.0101680209129454e-12
C123_130 V123 V130 8.080219273163007e-20

R123_131 V123 V131 44.49130819517425
L123_131 V123 V131 7.862216403782498e-13
C123_131 V123 V131 3.7056752027414064e-19

R123_132 V123 V132 162.5862915905314
L123_132 V123 V132 1.0576862918777189e-12
C123_132 V123 V132 5.135706254291714e-19

R123_133 V123 V133 291.25933398313197
L123_133 V123 V133 2.9419145278987245e-12
C123_133 V123 V133 8.044115939159352e-20

R123_134 V123 V134 269.9926691740634
L123_134 V123 V134 3.5658045614934507e-12
C123_134 V123 V134 1.7472481233698144e-19

R123_135 V123 V135 -101.02776875654389
L123_135 V123 V135 -4.00369892862563e-13
C123_135 V123 V135 -1.5965186499371538e-18

R123_136 V123 V136 330.04959415967375
L123_136 V123 V136 4.022834940694747e-12
C123_136 V123 V136 1.0617119690281558e-19

R123_137 V123 V137 317.12329133087826
L123_137 V123 V137 5.0654642979635716e-12
C123_137 V123 V137 8.129516120124646e-20

R123_138 V123 V138 -215.09808343855957
L123_138 V123 V138 -1.3379504144419269e-12
C123_138 V123 V138 -3.418923010715733e-19

R123_139 V123 V139 144.36526227720321
L123_139 V123 V139 3.2243633204927633e-13
C123_139 V123 V139 1.859604931109001e-18

R123_140 V123 V140 -154.12882216210855
L123_140 V123 V140 -1.5366529632999479e-12
C123_140 V123 V140 -2.843794589874518e-19

R123_141 V123 V141 -334.9167360891883
L123_141 V123 V141 -1.3732602913351439e-12
C123_141 V123 V141 -2.196940628392638e-19

R123_142 V123 V142 -165.8971695956556
L123_142 V123 V142 -3.457953611190861e-11
C123_142 V123 V142 5.695105569607117e-20

R123_143 V123 V143 1034.4438313146811
L123_143 V123 V143 -9.579040956786666e-13
C123_143 V123 V143 -3.2382499883383443e-19

R123_144 V123 V144 -646.9164390537608
L123_144 V123 V144 -7.486525427989309e-11
C123_144 V123 V144 1.3520121356745858e-19

R123_145 V123 V145 -237.61031056000184
L123_145 V123 V145 -3.961016002086043e-12
C123_145 V123 V145 -9.270571036283308e-20

R123_146 V123 V146 259.24886164886726
L123_146 V123 V146 2.311541849521873e-12
C123_146 V123 V146 1.6721117152783692e-19

R123_147 V123 V147 -79.39277049878602
L123_147 V123 V147 -8.489791459567787e-13
C123_147 V123 V147 -1.0043579060996142e-18

R123_148 V123 V148 236.48690470817795
L123_148 V123 V148 3.0796649880093444e-12
C123_148 V123 V148 3.001243738226839e-20

R123_149 V123 V149 1120.2795501904782
L123_149 V123 V149 7.08020582084751e-13
C123_149 V123 V149 5.359457085800808e-19

R123_150 V123 V150 123.70866648411932
L123_150 V123 V150 -4.3007195206454657e-11
C123_150 V123 V150 -6.973882751945357e-20

R123_151 V123 V151 -271.3491579648497
L123_151 V123 V151 1.6047673769992678e-12
C123_151 V123 V151 4.788414024560976e-19

R123_152 V123 V152 -746.8129632980496
L123_152 V123 V152 -2.8885040470444344e-12
C123_152 V123 V152 -9.902032762055591e-20

R123_153 V123 V153 126.86712548644395
L123_153 V123 V153 -1.473698267897519e-11
C123_153 V123 V153 -2.7587011700559534e-19

R123_154 V123 V154 1017.2383619230433
L123_154 V123 V154 -7.869630845507263e-12
C123_154 V123 V154 -1.3845219213604682e-19

R123_155 V123 V155 45.146210060166815
L123_155 V123 V155 4.785684047173358e-13
C123_155 V123 V155 6.547494201184481e-19

R123_156 V123 V156 520.3985793701685
L123_156 V123 V156 4.512681108074892e-12
C123_156 V123 V156 -9.735570320368964e-20

R123_157 V123 V157 407.776672234061
L123_157 V123 V157 -1.0836771909225311e-12
C123_157 V123 V157 -3.0892621119337005e-19

R123_158 V123 V158 -133.84352477308943
L123_158 V123 V158 4.739607259867028e-12
C123_158 V123 V158 1.68341543074816e-19

R123_159 V123 V159 -233.57814556643856
L123_159 V123 V159 -5.100669328845152e-13
C123_159 V123 V159 -7.569503925580286e-19

R123_160 V123 V160 -1091.1714852262683
L123_160 V123 V160 1.7455880118808792e-11
C123_160 V123 V160 1.473967566135057e-19

R123_161 V123 V161 -135.50248291168677
L123_161 V123 V161 2.750394731133797e-12
C123_161 V123 V161 3.2385396583821603e-19

R123_162 V123 V162 -201.494471600086
L123_162 V123 V162 2.1153358430260227e-12
C123_162 V123 V162 1.8758282299243074e-19

R123_163 V123 V163 -83.71313491908944
L123_163 V123 V163 5.8216562340884696e-12
C123_163 V123 V163 4.0680065136604667e-19

R123_164 V123 V164 -122.67373365121497
L123_164 V123 V164 -4.657734069324825e-12
C123_164 V123 V164 7.030809782803032e-20

R123_165 V123 V165 -402.23311512834374
L123_165 V123 V165 9.213340189402056e-12
C123_165 V123 V165 -9.857848309344782e-20

R123_166 V123 V166 141.5900967811482
L123_166 V123 V166 -5.063303576450817e-12
C123_166 V123 V166 -9.435443764195965e-20

R123_167 V123 V167 121.28768285930008
L123_167 V123 V167 1.2143615412896284e-12
C123_167 V123 V167 7.62073136108574e-20

R123_168 V123 V168 360.903109207421
L123_168 V123 V168 2.572916117089782e-12
C123_168 V123 V168 1.30000199861518e-19

R123_169 V123 V169 138.516854446933
L123_169 V123 V169 -1.8673242670684173e-12
C123_169 V123 V169 -4.5538383824393e-19

R123_170 V123 V170 274.1545173695413
L123_170 V123 V170 1.1633849796421249e-11
C123_170 V123 V170 3.746893624341129e-20

R123_171 V123 V171 -2245.333717372241
L123_171 V123 V171 -1.2327049514970523e-12
C123_171 V123 V171 -2.9630378306150096e-19

R123_172 V123 V172 190.5568413306984
L123_172 V123 V172 -1.8361200748441277e-11
C123_172 V123 V172 -1.5930851797393294e-19

R123_173 V123 V173 -304.65609147276285
L123_173 V123 V173 2.441608301165492e-12
C123_173 V123 V173 3.259004860395215e-19

R123_174 V123 V174 -174.26371507819314
L123_174 V123 V174 2.4838551832534134e-11
C123_174 V123 V174 -1.9859113919822811e-19

R123_175 V123 V175 -293.33210852127274
L123_175 V123 V175 8.473978932429126e-13
C123_175 V123 V175 7.5480567635605785e-19

R123_176 V123 V176 -270.9727941467733
L123_176 V123 V176 -6.420749251028381e-12
C123_176 V123 V176 -1.0039869809529388e-19

R123_177 V123 V177 -309.46578686556217
L123_177 V123 V177 -5.9806066496835085e-12
C123_177 V123 V177 2.9053198938927376e-21

R123_178 V123 V178 -172.1674288746916
L123_178 V123 V178 -1.710477035239353e-12
C123_178 V123 V178 4.260041690960134e-20

R123_179 V123 V179 84.73181552375125
L123_179 V123 V179 2.75639632642595e-11
C123_179 V123 V179 -6.270788920315527e-19

R123_180 V123 V180 -214.62831921477064
L123_180 V123 V180 -2.8852632222250498e-12
C123_180 V123 V180 1.9299767682093986e-20

R123_181 V123 V181 292.52645362862506
L123_181 V123 V181 3.369135802213458e-12
C123_181 V123 V181 -3.193504351126417e-20

R123_182 V123 V182 97.2497664050225
L123_182 V123 V182 1.1432597683731423e-12
C123_182 V123 V182 1.5277294932653132e-19

R123_183 V123 V183 -102.13029249360085
L123_183 V123 V183 -5.984205870928213e-13
C123_183 V123 V183 3.3594636072433895e-20

R123_184 V123 V184 238.61976690989047
L123_184 V123 V184 -4.958609408150114e-12
C123_184 V123 V184 -1.180586177318652e-19

R123_185 V123 V185 461.8433275589135
L123_185 V123 V185 1.200305540755275e-11
C123_185 V123 V185 3.80485216749017e-20

R123_186 V123 V186 307.630930600765
L123_186 V123 V186 -7.056218165791582e-12
C123_186 V123 V186 -2.3651779524096723e-19

R123_187 V123 V187 -232.120784002702
L123_187 V123 V187 4.96980078086439e-13
C123_187 V123 V187 7.640088767850334e-19

R123_188 V123 V188 931.8231115468759
L123_188 V123 V188 1.5060728224557682e-12
C123_188 V123 V188 1.7196888694671886e-19

R123_189 V123 V189 -389.4778544778607
L123_189 V123 V189 -2.7419415543641173e-12
C123_189 V123 V189 -1.4058429376835456e-19

R123_190 V123 V190 -123.14946017901144
L123_190 V123 V190 -2.55977016303799e-12
C123_190 V123 V190 2.3655676879784266e-20

R123_191 V123 V191 133.24783939732723
L123_191 V123 V191 2.8238050748855416e-12
C123_191 V123 V191 -6.628807924889533e-19

R123_192 V123 V192 -299.164295021215
L123_192 V123 V192 3.837223034423892e-12
C123_192 V123 V192 -1.2232887196023086e-20

R123_193 V123 V193 -635.3416308283261
L123_193 V123 V193 1.1120235732981872e-11
C123_193 V123 V193 -2.0492124561962135e-20

R123_194 V123 V194 227.64585037207868
L123_194 V123 V194 -6.931062982257116e-12
C123_194 V123 V194 -3.297798911766984e-19

R123_195 V123 V195 -236.26144671665736
L123_195 V123 V195 -1.9121358387209545e-12
C123_195 V123 V195 8.683882579747367e-19

R123_196 V123 V196 895.9824346303246
L123_196 V123 V196 -8.772247506742238e-13
C123_196 V123 V196 -4.711470169682211e-19

R123_197 V123 V197 694.6095893605964
L123_197 V123 V197 8.696815266828068e-12
C123_197 V123 V197 1.1585356977400726e-19

R123_198 V123 V198 200.20330508941
L123_198 V123 V198 2.6046300447582025e-12
C123_198 V123 V198 7.756818101813544e-20

R123_199 V123 V199 -617.4792570445886
L123_199 V123 V199 1.2333002560865923e-11
C123_199 V123 V199 4.4348432316552505e-21

R123_200 V123 V200 -44774.44000774768
L123_200 V123 V200 2.228075479645521e-12
C123_200 V123 V200 3.1636072175881455e-19

R124_124 V124 0 213.69836208241745
L124_124 V124 0 1.4917858347427606e-13
C124_124 V124 0 4.388732848424843e-18

R124_125 V124 V125 250.80645289875795
L124_125 V124 V125 -3.1462994891351686e-12
C124_125 V124 V125 -4.494302218425818e-20

R124_126 V124 V126 363.38003135809777
L124_126 V124 V126 -7.573423178368114e-13
C124_126 V124 V126 -5.801698328260505e-19

R124_127 V124 V127 216.96431472871362
L124_127 V124 V127 -7.477928619145972e-13
C124_127 V124 V127 -9.275041456921709e-19

R124_128 V124 V128 -74.57240579907165
L124_128 V124 V128 6.016944315292908e-13
C124_128 V124 V128 9.014661189870308e-19

R124_129 V124 V129 -123.56867077793754
L124_129 V124 V129 -2.9749641902204368e-12
C124_129 V124 V129 -2.8466049542072883e-19

R124_130 V124 V130 -1196.5483478545443
L124_130 V124 V130 2.4844465642071917e-12
C124_130 V124 V130 2.1173942257438553e-19

R124_131 V124 V131 -695.7926467770855
L124_131 V124 V131 9.412465067298133e-13
C124_131 V124 V131 7.123819527499662e-19

R124_132 V124 V132 38.440545820836796
L124_132 V124 V132 4.430533408671797e-13
C124_132 V124 V132 1.3380643317786716e-18

R124_133 V124 V133 263.2657422380934
L124_133 V124 V133 1.4604172202822963e-12
C124_133 V124 V133 5.110734884116912e-19

R124_134 V124 V134 202.46667431205753
L124_134 V124 V134 1.1155234341532842e-12
C124_134 V124 V134 8.075123378489081e-19

R124_135 V124 V135 2063.3393400480254
L124_135 V124 V135 1.1807913629294574e-12
C124_135 V124 V135 7.303179860177907e-19

R124_136 V124 V136 -154.58313901650942
L124_136 V124 V136 -3.1215650747718056e-13
C124_136 V124 V136 -2.4091785694727296e-18

R124_137 V124 V137 313.18447566483326
L124_137 V124 V137 -3.35900850108005e-12
C124_137 V124 V137 -2.2343139657785413e-19

R124_138 V124 V138 -246.1445303701071
L124_138 V124 V138 -7.492180255422746e-13
C124_138 V124 V138 -8.053501016779712e-19

R124_139 V124 V139 -1431.7630739539868
L124_139 V124 V139 -6.645591950062594e-13
C124_139 V124 V139 -1.0380887007036749e-18

R124_140 V124 V140 6407.475032909364
L124_140 V124 V140 3.721498186815365e-13
C124_140 V124 V140 2.4019302738674857e-18

R124_141 V124 V141 -537.5168661959276
L124_141 V124 V141 -1.2238027424228498e-12
C124_141 V124 V141 -3.9804579827579445e-19

R124_142 V124 V142 -173.53876873677618
L124_142 V124 V142 -2.683588378390118e-12
C124_142 V124 V142 -8.263456046208291e-20

R124_143 V124 V143 -628.3055083457256
L124_143 V124 V143 -6.457097037572161e-12
C124_143 V124 V143 1.116208181208952e-19

R124_144 V124 V144 291.4072128347537
L124_144 V124 V144 -2.9051240404732764e-12
C124_144 V124 V144 -3.226332810476642e-19

R124_145 V124 V145 -240.99829362009862
L124_145 V124 V145 9.232809734302506e-12
C124_145 V124 V145 1.3175726824101205e-19

R124_146 V124 V146 230.49246220082225
L124_146 V124 V146 7.64221943797459e-13
C124_146 V124 V146 3.744323032403909e-19

R124_147 V124 V147 1964.9230163589357
L124_147 V124 V147 -1.2128930257627929e-11
C124_147 V124 V147 5.4273246878592974e-21

R124_148 V124 V148 -71.55561399984069
L124_148 V124 V148 -3.1702531079897464e-13
C124_148 V124 V148 -1.4766365752914137e-18

R124_149 V124 V149 -1602.8733073356589
L124_149 V124 V149 1.0253894121762519e-12
C124_149 V124 V149 2.543965262309552e-19

R124_150 V124 V150 157.73466113461976
L124_150 V124 V150 -1.850974443089571e-12
C124_150 V124 V150 -2.643130912867978e-19

R124_151 V124 V151 -587.8122480897066
L124_151 V124 V151 2.074528821274599e-12
C124_151 V124 V151 -5.666047529306068e-20

R124_152 V124 V152 -575.8862613929256
L124_152 V124 V152 4.393810083160056e-13
C124_152 V124 V152 5.11659424499912e-19

R124_153 V124 V153 140.73216608322195
L124_153 V124 V153 1.5109366514004557e-12
C124_153 V124 V153 -3.7274231882032295e-22

R124_154 V124 V154 807.4311514186954
L124_154 V124 V154 1.59924003569415e-12
C124_154 V124 V154 -1.547436172624336e-19

R124_155 V124 V155 168.3457827778365
L124_155 V124 V155 2.8944003558383907e-12
C124_155 V124 V155 -1.143346265870789e-19

R124_156 V124 V156 65.40518080595187
L124_156 V124 V156 8.988612581653447e-12
C124_156 V124 V156 1.1518795797815124e-18

R124_157 V124 V157 386.01337278722053
L124_157 V124 V157 -6.177948620412232e-13
C124_157 V124 V157 -6.853572908963276e-19

R124_158 V124 V158 -116.20837193805671
L124_158 V124 V158 -2.7048861672549e-12
C124_158 V124 V158 1.5529110668730264e-19

R124_159 V124 V159 -593.6149728346186
L124_159 V124 V159 3.771625809710025e-12
C124_159 V124 V159 2.986981984139421e-19

R124_160 V124 V160 513.5701197599877
L124_160 V124 V160 -9.2023349003527e-13
C124_160 V124 V160 -8.72593000468045e-19

R124_161 V124 V161 -123.0170351465051
L124_161 V124 V161 1.0106548123872775e-12
C124_161 V124 V161 4.349254807833766e-19

R124_162 V124 V162 -214.3703094359976
L124_162 V124 V162 1.6236206238687579e-12
C124_162 V124 V162 1.7403485588937478e-19

R124_163 V124 V163 -251.49054303504147
L124_163 V124 V163 -3.0960883240374047e-12
C124_163 V124 V163 -1.8385282486764091e-19

R124_164 V124 V164 -60.515991470948606
L124_164 V124 V164 -5.223073024555545e-12
C124_164 V124 V164 6.305810900299703e-19

R124_165 V124 V165 -334.5600018651627
L124_165 V124 V165 -1.7570371465339714e-12
C124_165 V124 V165 -2.485121793639644e-19

R124_166 V124 V166 135.0604883076366
L124_166 V124 V166 -2.288213743229001e-12
C124_166 V124 V166 -3.7594364393336194e-19

R124_167 V124 V167 -325.331341775851
L124_167 V124 V167 4.7494278378390765e-12
C124_167 V124 V167 2.0570159978220834e-19

R124_168 V124 V168 82.59020047503795
L124_168 V124 V168 5.305188365558124e-13
C124_168 V124 V168 1.4889973014555294e-20

R124_169 V124 V169 138.87758188434293
L124_169 V124 V169 -2.029891625817349e-12
C124_169 V124 V169 -6.57458608458953e-19

R124_170 V124 V170 386.1075310264798
L124_170 V124 V170 2.2245962668728765e-12
C124_170 V124 V170 6.101861651090856e-20

R124_171 V124 V171 205.3193229964359
L124_171 V124 V171 1.3168465384563198e-12
C124_171 V124 V171 -7.740732091930717e-20

R124_172 V124 V172 -434.87007233721175
L124_172 V124 V172 -4.863887430277557e-13
C124_172 V124 V172 -3.3734603381971145e-19

R124_173 V124 V173 -214.70743099301836
L124_173 V124 V173 1.2776933489130167e-12
C124_173 V124 V173 5.539720138959462e-19

R124_174 V124 V174 -208.2253313722528
L124_174 V124 V174 5.085432522924561e-11
C124_174 V124 V174 -1.0638763400028655e-19

R124_175 V124 V175 -2048.582467462767
L124_175 V124 V175 -1.3299536046310063e-12
C124_175 V124 V175 -1.726339070872814e-19

R124_176 V124 V176 -204.8596623157787
L124_176 V124 V176 7.24391365293345e-13
C124_176 V124 V176 1.2395510694774414e-18

R124_177 V124 V177 -248.79953837009123
L124_177 V124 V177 -3.1207511367737018e-12
C124_177 V124 V177 -1.0451426712843019e-19

R124_178 V124 V178 -159.50106197589477
L124_178 V124 V178 -1.2439417090005898e-12
C124_178 V124 V178 4.011054488176109e-20

R124_179 V124 V179 -354.1145409113282
L124_179 V124 V179 -1.5291397835481478e-12
C124_179 V124 V179 -9.310630324575542e-21

R124_180 V124 V180 71.86705696979256
L124_180 V124 V180 2.7475814749383638e-11
C124_180 V124 V180 -9.928157797748537e-19

R124_181 V124 V181 254.666329858325
L124_181 V124 V181 1.1755138343886279e-11
C124_181 V124 V181 -1.226457371585421e-19

R124_182 V124 V182 117.98686226039706
L124_182 V124 V182 2.1164947555908066e-12
C124_182 V124 V182 -6.022094752626424e-20

R124_183 V124 V183 344.31038644144513
L124_183 V124 V183 -7.695648580723188e-12
C124_183 V124 V183 -2.8248675895453805e-19

R124_184 V124 V184 -125.13983412727927
L124_184 V124 V184 -5.371019034549141e-13
C124_184 V124 V184 1.4829401760907483e-19

R124_185 V124 V185 797.6611371148143
L124_185 V124 V185 9.297757182790159e-12
C124_185 V124 V185 1.3831842001777397e-19

R124_186 V124 V186 234.38768256301248
L124_186 V124 V186 -1.461806953338124e-12
C124_186 V124 V186 -4.689768270165445e-20

R124_187 V124 V187 800.7756638959432
L124_187 V124 V187 -3.5407529514941264e-12
C124_187 V124 V187 1.5222242726289842e-19

R124_188 V124 V188 -131.70336663129942
L124_188 V124 V188 2.774328276417087e-13
C124_188 V124 V188 7.3853212623763e-19

R124_189 V124 V189 -462.5217231515907
L124_189 V124 V189 -1.9794600897335223e-12
C124_189 V124 V189 -1.7568201265125684e-19

R124_190 V124 V190 -116.77518712705722
L124_190 V124 V190 -5.032351225658785e-12
C124_190 V124 V190 6.4754935881181665e-21

R124_191 V124 V191 -214.95971823629955
L124_191 V124 V191 6.980798656552843e-13
C124_191 V124 V191 3.975542750498897e-19

R124_192 V124 V192 124.24695528620515
L124_192 V124 V192 -5.899057839777478e-13
C124_192 V124 V192 -1.1099960233243298e-18

R124_193 V124 V193 4827.864307832282
L124_193 V124 V193 1.4757274778231983e-11
C124_193 V124 V193 -1.5294872865903376e-19

R124_194 V124 V194 260.17119871953474
L124_194 V124 V194 -1.4404213032038438e-12
C124_194 V124 V194 -7.706579349524545e-19

R124_195 V124 V195 348.8891597096866
L124_195 V124 V195 -5.156828514915358e-13
C124_195 V124 V195 -1.1678895393880069e-18

R124_196 V124 V196 -201.080202822712
L124_196 V124 V196 7.256492691893013e-13
C124_196 V124 V196 1.9468605127276467e-18

R124_197 V124 V197 781.5435067812128
L124_197 V124 V197 3.079401077401126e-12
C124_197 V124 V197 2.762975881259263e-19

R124_198 V124 V198 235.38059389900843
L124_198 V124 V198 6.919733287239535e-12
C124_198 V124 V198 -2.0043991961873175e-19

R124_199 V124 V199 -4349.988464744284
L124_199 V124 V199 3.81895103214918e-12
C124_199 V124 V199 1.5031854248582969e-19

R124_200 V124 V200 -414.70938100218785
L124_200 V124 V200 -1.7679412156530464e-11
C124_200 V124 V200 -2.0710594838829107e-19

R125_125 V125 0 130.42535773388454
L125_125 V125 0 3.174618691196873e-13
C125_125 V125 0 7.627461154096558e-19

R125_126 V125 V126 -631.6012399585692
L125_126 V125 V126 -2.683860979671313e-12
C125_126 V125 V126 -1.709892111638959e-20

R125_127 V125 V127 1119.2369188138107
L125_127 V125 V127 -7.704665699241091e-12
C125_127 V125 V127 -1.0384740548050761e-19

R125_128 V125 V128 209.19930285973257
L125_128 V125 V128 1.90450705544364e-11
C125_128 V125 V128 -6.588565387960844e-20

R125_129 V125 V129 75.66571728005991
L125_129 V125 V129 3.2727987228141058e-12
C125_129 V125 V129 7.627107885327746e-20

R125_130 V125 V130 251.4672553170567
L125_130 V125 V130 1.7418438363023145e-12
C125_130 V125 V130 1.937511754855552e-19

R125_131 V125 V131 -6454.968434200925
L125_131 V125 V131 8.335295136133007e-12
C125_131 V125 V131 3.892226408001457e-20

R125_132 V125 V132 -193.37877898802506
L125_132 V125 V132 3.3326485468970043e-12
C125_132 V125 V132 1.563145353280969e-19

R125_133 V125 V133 170.8452314191989
L125_133 V125 V133 1.4229050655254676e-12
C125_133 V125 V133 2.3409132360627925e-19

R125_134 V125 V134 -161.80499700482085
L125_134 V125 V134 -3.570337005752639e-12
C125_134 V125 V134 -2.343338312483115e-19

R125_135 V125 V135 -248.0772210807293
L125_135 V125 V135 1.0850759538895364e-11
C125_135 V125 V135 1.4553764747205206e-19

R125_136 V125 V136 -306.2445050462428
L125_136 V125 V136 -6.3819202558204565e-12
C125_136 V125 V136 3.058876381470436e-20

R125_137 V125 V137 -55.42887875066135
L125_137 V125 V137 1.1479642673430551e-11
C125_137 V125 V137 1.63442114629187e-19

R125_138 V125 V138 851.1248024123643
L125_138 V125 V138 -8.361672104772276e-12
C125_138 V125 V138 1.2844233558018528e-19

R125_139 V125 V139 609.0002166793635
L125_139 V125 V139 -4.753883275789214e-12
C125_139 V125 V139 -2.0283180008013482e-19

R125_140 V125 V140 -3708.2273095473493
L125_140 V125 V140 2.8791924252230453e-11
C125_140 V125 V140 -8.161338538634293e-20

R125_141 V125 V141 9162.563864535923
L125_141 V125 V141 -1.4702319320898016e-12
C125_141 V125 V141 -3.6172217988806024e-19

R125_142 V125 V142 85.43873271345304
L125_142 V125 V142 2.000225697790268e-12
C125_142 V125 V142 4.92162417125163e-20

R125_143 V125 V143 135.63858048927418
L125_143 V125 V143 6.37682115575771e-12
C125_143 V125 V143 5.1171273613633134e-21

R125_144 V125 V144 93.49022707034615
L125_144 V125 V144 9.185429170399856e-12
C125_144 V125 V144 -6.233669697580413e-20

R125_145 V125 V145 48.857072689066634
L125_145 V125 V145 -2.8701885439464563e-12
C125_145 V125 V145 -1.32767150927827e-19

R125_146 V125 V146 234.1476630648501
L125_146 V125 V146 -6.9850408359596075e-12
C125_146 V125 V146 -3.007346483699164e-20

R125_147 V125 V147 475.9398749405932
L125_147 V125 V147 -6.4435062102917195e-12
C125_147 V125 V147 1.0482409411692327e-19

R125_148 V125 V148 -278.7687668902672
L125_148 V125 V148 -2.5207200937647617e-12
C125_148 V125 V148 2.0405599785008182e-20

R125_149 V125 V149 -199.11238434698802
L125_149 V125 V149 1.2492315461007096e-12
C125_149 V125 V149 2.7177233831408193e-19

R125_150 V125 V150 -39.8034273135319
L125_150 V125 V150 -2.129093748008344e-12
C125_150 V125 V150 -1.8970558026016563e-19

R125_151 V125 V151 -69.24335378933588
L125_151 V125 V151 -3.4469605377640746e-12
C125_151 V125 V151 -5.296462810748648e-20

R125_152 V125 V152 -178.29147789488954
L125_152 V125 V152 7.462781134821325e-11
C125_152 V125 V152 6.787189861988866e-21

R125_153 V125 V153 -52.22621312189822
L125_153 V125 V153 4.244669579304735e-12
C125_153 V125 V153 1.2495146941602082e-19

R125_154 V125 V154 -406.5936603972365
L125_154 V125 V154 3.5809903241655402e-12
C125_154 V125 V154 1.8386424102055026e-19

R125_155 V125 V155 77.30293405758198
L125_155 V125 V155 3.668344690859189e-12
C125_155 V125 V155 -4.3498922474330876e-20

R125_156 V125 V156 -217.90183097985937
L125_156 V125 V156 8.0421038826978e-12
C125_156 V125 V156 3.77428967824037e-20

R125_157 V125 V157 -774.0354537242349
L125_157 V125 V157 -1.469266517928895e-12
C125_157 V125 V157 -1.8616237916633194e-19

R125_158 V125 V158 63.32826647174015
L125_158 V125 V158 4.377344774639348e-12
C125_158 V125 V158 -8.18207505587918e-20

R125_159 V125 V159 580.6362685377426
L125_159 V125 V159 2.2419582192791042e-12
C125_159 V125 V159 1.5969108398023697e-19

R125_160 V125 V160 86.88873549554071
L125_160 V125 V160 2.2447860254568104e-12
C125_160 V125 V160 7.917769932509925e-20

R125_161 V125 V161 144.3315786453133
L125_161 V125 V161 9.791847511798338e-10
C125_161 V125 V161 -2.5661939555419647e-20

R125_162 V125 V162 372.199933874075
L125_162 V125 V162 8.661421281978898e-12
C125_162 V125 V162 9.100324959654152e-20

R125_163 V125 V163 -357.6747453694856
L125_163 V125 V163 -9.438100534561796e-12
C125_163 V125 V163 -2.4350080170967302e-20

R125_164 V125 V164 -191.71105493035665
L125_164 V125 V164 -5.084173672292991e-12
C125_164 V125 V164 -9.010515988304495e-21

R125_165 V125 V165 1646.5059147568654
L125_165 V125 V165 -1.5509346480231375e-12
C125_165 V125 V165 -1.2475873249740863e-19

R125_166 V125 V166 -45.525357761918166
L125_166 V125 V166 -2.6509276377467718e-12
C125_166 V125 V166 -4.702903198557277e-22

R125_167 V125 V167 -271.40171678376964
L125_167 V125 V167 -2.669834207368508e-12
C125_167 V125 V167 -1.089900928580692e-19

R125_168 V125 V168 296.52794014400763
L125_168 V125 V168 -2.3089153348711662e-12
C125_168 V125 V168 -1.947626554839432e-19

R125_169 V125 V169 -143.82242492861266
L125_169 V125 V169 1.4064301360139524e-12
C125_169 V125 V169 1.6310457292094227e-19

R125_170 V125 V170 81.79123165026706
L125_170 V125 V170 4.536425553858443e-11
C125_170 V125 V170 -5.041370594911126e-20

R125_171 V125 V171 139.92424045152566
L125_171 V125 V171 3.811170011421336e-12
C125_171 V125 V171 8.983337600868146e-20

R125_172 V125 V172 180.28934563589098
L125_172 V125 V172 4.1381905708305086e-12
C125_172 V125 V172 1.1021030855589798e-19

R125_173 V125 V173 605.1269356445566
L125_173 V125 V173 -7.104032669806783e-12
C125_173 V125 V173 5.3689218165215704e-20

R125_174 V125 V174 74.15262646905964
L125_174 V125 V174 1.3005159802803277e-12
C125_174 V125 V174 4.0048845572650824e-20

R125_175 V125 V175 -354.1879193858368
L125_175 V125 V175 1.6228293775743768e-12
C125_175 V125 V175 7.860056262433185e-20

R125_176 V125 V176 -222.1549834832975
L125_176 V125 V176 1.157528029542827e-12
C125_176 V125 V176 1.5453348796255487e-19

R125_177 V125 V177 267.8286508336474
L125_177 V125 V177 4.567229330926015e-12
C125_177 V125 V177 4.3792919232363946e-20

R125_178 V125 V178 -71.95768027337215
L125_178 V125 V178 -2.930456173049973e-12
C125_178 V125 V178 8.384144956544665e-21

R125_179 V125 V179 1009.5432838211734
L125_179 V125 V179 -2.0303241765396713e-12
C125_179 V125 V179 -7.578369489110887e-20

R125_180 V125 V180 -206.01580603901067
L125_180 V125 V180 -1.481597049370843e-12
C125_180 V125 V180 -7.914922163158749e-20

R125_181 V125 V181 -725.700235704626
L125_181 V125 V181 -1.3125883797189675e-12
C125_181 V125 V181 -4.1931517643877873e-19

R125_182 V125 V182 -690.5760499296133
L125_182 V125 V182 3.654738228582832e-11
C125_182 V125 V182 2.974036216748703e-20

R125_183 V125 V183 -6570.7987184152025
L125_183 V125 V183 -4.71615972433767e-12
C125_183 V125 V183 -5.604807455000408e-20

R125_184 V125 V184 165.0791206425087
L125_184 V125 V184 -3.422362905194733e-12
C125_184 V125 V184 -6.939314190333096e-20

R125_185 V125 V185 -172.74116522404896
L125_185 V125 V185 -3.970354764230022e-12
C125_185 V125 V185 1.9806000558027176e-19

R125_186 V125 V186 120.10710108043162
L125_186 V125 V186 -9.178354628122804e-12
C125_186 V125 V186 -1.1128046942881831e-19

R125_187 V125 V187 1552.8629188194152
L125_187 V125 V187 4.0048428770184885e-12
C125_187 V125 V187 3.691259346064299e-20

R125_188 V125 V188 592.0649730180626
L125_188 V125 V188 2.2619132752100686e-12
C125_188 V125 V188 3.292666072126166e-20

R125_189 V125 V189 381.79061114012876
L125_189 V125 V189 8.210979953724943e-13
C125_189 V125 V189 2.848512694100661e-19

R125_190 V125 V190 -259.86332454549466
L125_190 V125 V190 -1.3389872359465674e-11
C125_190 V125 V190 -5.862430972437251e-20

R125_191 V125 V191 -222.08080816258519
L125_191 V125 V191 3.402648036566372e-12
C125_191 V125 V191 1.8761051256932252e-19

R125_192 V125 V192 -157.97178408080475
L125_192 V125 V192 3.9112803549176954e-12
C125_192 V125 V192 2.270226073263588e-19

R125_193 V125 V193 287.35353940162025
L125_193 V125 V193 -2.4456172564410764e-12
C125_193 V125 V193 -8.077291035914398e-20

R125_194 V125 V194 -305.48275419050765
L125_194 V125 V194 1.5470012341109943e-12
C125_194 V125 V194 1.2700568425223177e-19

R125_195 V125 V195 744.8889958529676
L125_195 V125 V195 -2.4232349716743737e-12
C125_195 V125 V195 -2.814120520290566e-19

R125_196 V125 V196 7220.916432416433
L125_196 V125 V196 -1.0562346693450815e-09
C125_196 V125 V196 -1.900686213865251e-19

R125_197 V125 V197 -2790.197825418248
L125_197 V125 V197 -3.018752746881281e-12
C125_197 V125 V197 -1.9736995371871038e-19

R125_198 V125 V198 -2525.307814144508
L125_198 V125 V198 -3.036543386562224e-11
C125_198 V125 V198 -8.63834698962008e-22

R125_199 V125 V199 449.8294414446449
L125_199 V125 V199 -2.1174924122861003e-11
C125_199 V125 V199 -3.788451241024555e-20

R125_200 V125 V200 104.71396753558436
L125_200 V125 V200 -3.1816062431696357e-12
C125_200 V125 V200 -1.0532872683553594e-19

R126_126 V126 0 -27.90938939417277
L126_126 V126 0 3.048707856491897e-13
C126_126 V126 0 9.324571360536544e-19

R126_127 V126 V127 -73.38886962179411
L126_127 V126 V127 -4.8440579991936664e-11
C126_127 V126 V127 8.654503044470706e-20

R126_128 V126 V128 -119.9859851789935
L126_128 V126 V128 3.318159822367305e-12
C126_128 V126 V128 -5.434299596359985e-22

R126_129 V126 V129 -91.02500048465234
L126_129 V126 V129 -2.2296882689685303e-12
C126_129 V126 V129 -2.0318787742501067e-19

R126_130 V126 V130 37.38991582021018
L126_130 V126 V130 8.322305635631647e-13
C126_130 V126 V130 4.104393669105163e-19

R126_131 V126 V131 60.541101655700224
L126_131 V126 V131 1.48615920943658e-12
C126_131 V126 V131 2.5842483822092925e-19

R126_132 V126 V132 64.28939819622462
L126_132 V126 V132 1.0350654866538334e-12
C126_132 V126 V132 5.466082703558279e-19

R126_133 V126 V133 819.0675351066909
L126_133 V126 V133 2.1737878981892243e-12
C126_133 V126 V133 2.5159253066891575e-19

R126_134 V126 V134 70.73029781938882
L126_134 V126 V134 2.5427783843361005e-12
C126_134 V126 V134 2.413372051978869e-19

R126_135 V126 V135 120.29250624862556
L126_135 V126 V135 -2.2493024629436466e-12
C126_135 V126 V135 -4.441966679447569e-19

R126_136 V126 V136 65.01227715064725
L126_136 V126 V136 -1.589414294593517e-12
C126_136 V126 V136 -4.1592635350183845e-19

R126_137 V126 V137 89.81874811000175
L126_137 V126 V137 4.8025108916481294e-12
C126_137 V126 V137 5.2713943854690816e-20

R126_138 V126 V138 -41.03779255003136
L126_138 V126 V138 -8.850945018050064e-13
C126_138 V126 V138 -4.2095222747040605e-19

R126_139 V126 V139 -42.41664197469623
L126_139 V126 V139 2.2738648840090536e-12
C126_139 V126 V139 5.390647560123812e-19

R126_140 V126 V140 -27.055479495313833
L126_140 V126 V140 8.729963847574689e-12
C126_140 V126 V140 3.3003556694898103e-19

R126_141 V126 V141 129.5144375606766
L126_141 V126 V141 -1.496027207799672e-12
C126_141 V126 V141 -3.6345421177786945e-19

R126_142 V126 V142 -76.7630575613894
L126_142 V126 V142 1.5501989539064158e-09
C126_142 V126 V142 5.0059302229409307e-20

R126_143 V126 V143 113.81609130910667
L126_143 V126 V143 -2.5057798511315594e-12
C126_143 V126 V143 -1.0665640186947628e-19

R126_144 V126 V144 114.16871848876187
L126_144 V126 V144 5.609767071257998e-11
C126_144 V126 V144 -4.9889536115383504e-20

R126_145 V126 V145 -68.8471508728378
L126_145 V126 V145 -3.4310506715485436e-12
C126_145 V126 V145 -6.006570751190389e-20

R126_146 V126 V146 36.47433034973691
L126_146 V126 V146 1.1008707180891806e-12
C126_146 V126 V146 1.2258590488299175e-19

R126_147 V126 V147 176.94824029234505
L126_147 V126 V147 -2.7105562236887365e-12
C126_147 V126 V147 -5.516909073333361e-19

R126_148 V126 V148 89.16489807909747
L126_148 V126 V148 -1.3041419544710704e-12
C126_148 V126 V148 -3.266507634409444e-19

R126_149 V126 V149 -313.9969712751657
L126_149 V126 V149 7.508997902036232e-13
C126_149 V126 V149 4.720600309285279e-19

R126_150 V126 V150 34.708503347958235
L126_150 V126 V150 -5.253299274075648e-12
C126_150 V126 V150 -1.344411818531728e-19

R126_151 V126 V151 -141.34212207706756
L126_151 V126 V151 3.934521805260942e-12
C126_151 V126 V151 2.497810106066554e-19

R126_152 V126 V152 -64.57264348599811
L126_152 V126 V152 2.639194919840272e-12
C126_152 V126 V152 9.03544909454152e-20

R126_153 V126 V153 118.773706518443
L126_153 V126 V153 1.6235975812164192e-11
C126_153 V126 V153 -4.995719620478859e-20

R126_154 V126 V154 -37.93573140973488
L126_154 V126 V154 -3.234094715769925e-12
C126_154 V126 V154 5.234747484370986e-21

R126_155 V126 V155 -260.7056194261719
L126_155 V126 V155 9.725132901860293e-13
C126_155 V126 V155 2.7170692785453796e-19

R126_156 V126 V156 114.61376391870522
L126_156 V126 V156 5.7676878909558015e-12
C126_156 V126 V156 2.775119959795977e-19

R126_157 V126 V157 115.24523644729943
L126_157 V126 V157 -7.7352239993199e-13
C126_157 V126 V157 -3.658704231561969e-19

R126_158 V126 V158 -180.58021884843325
L126_158 V126 V158 3.778311962525612e-12
C126_158 V126 V158 1.5324129604336618e-19

R126_159 V126 V159 59.77279610919932
L126_159 V126 V159 -2.1682511378068493e-12
C126_159 V126 V159 -1.9591679194222217e-19

R126_160 V126 V160 70.69477506146289
L126_160 V126 V160 1.7873648518562703e-11
C126_160 V126 V160 -1.501787628792118e-19

R126_161 V126 V161 -53.93783044253598
L126_161 V126 V161 2.4692692727156224e-12
C126_161 V126 V161 1.836855072729302e-19

R126_162 V126 V162 254.70249278959736
L126_162 V126 V162 1.402390222280893e-12
C126_162 V126 V162 1.0214825731837621e-19

R126_163 V126 V163 -54.97487692635899
L126_163 V126 V163 -3.1887460813892673e-12
C126_163 V126 V163 1.241700045357745e-19

R126_164 V126 V164 -41.69865855247153
L126_164 V126 V164 -1.9998260363568418e-12
C126_164 V126 V164 1.4507829146401737e-19

R126_165 V126 V165 295.74101689917023
L126_165 V126 V165 -5.82096851340288e-11
C126_165 V126 V165 -1.0637242650584576e-19

R126_166 V126 V166 69.54582130408792
L126_166 V126 V166 -2.2264353111665025e-12
C126_166 V126 V166 -1.3823696897196829e-19

R126_167 V126 V167 -752.3068292033895
L126_167 V126 V167 3.6158117688405195e-12
C126_167 V126 V167 7.318077658728614e-20

R126_168 V126 V168 -273.16401109476806
L126_168 V126 V168 1.6661669865593707e-12
C126_168 V126 V168 -6.925426752366264e-21

R126_169 V126 V169 42.41461885579407
L126_169 V126 V169 -6.2825555867265624e-12
C126_169 V126 V169 -2.5736480051664237e-19

R126_170 V126 V170 -556.8466815178701
L126_170 V126 V170 3.0954688301752826e-12
C126_170 V126 V170 4.015994675826013e-20

R126_171 V126 V171 60.45368591171125
L126_171 V126 V171 1.9479631474330436e-12
C126_171 V126 V171 -1.3055414018556873e-19

R126_172 V126 V172 54.288033944089776
L126_172 V126 V172 -5.838095846620898e-12
C126_172 V126 V172 -1.2617852159659724e-19

R126_173 V126 V173 -58.441399062639796
L126_173 V126 V173 2.5540534297604527e-12
C126_173 V126 V173 3.234375655146597e-19

R126_174 V126 V174 -111.16920408930126
L126_174 V126 V174 -4.941972114824383e-12
C126_174 V126 V174 -9.763466372717502e-20

R126_175 V126 V175 -540.2176657345576
L126_175 V126 V175 7.1945817063127775e-12
C126_175 V126 V175 2.747466392150844e-19

R126_176 V126 V176 -170.72908456040236
L126_176 V126 V176 3.5821371747923966e-12
C126_176 V126 V176 2.721516533469447e-19

R126_177 V126 V177 -118.25356212936441
L126_177 V126 V177 -3.0670390062539698e-12
C126_177 V126 V177 -3.3030108475877094e-20

R126_178 V126 V178 -781.8851865693866
L126_178 V126 V178 -3.359311213476503e-12
C126_178 V126 V178 2.5908278166678496e-20

R126_179 V126 V179 -108.99313670168891
L126_179 V126 V179 -1.6643543509642143e-12
C126_179 V126 V179 -2.4303753092346455e-19

R126_180 V126 V180 -80.57370931040619
L126_180 V126 V180 -1.8264579517081594e-12
C126_180 V126 V180 -2.0138471082237468e-19

R126_181 V126 V181 65.78667338936901
L126_181 V126 V181 2.6447443085508216e-11
C126_181 V126 V181 -2.133033603827886e-19

R126_182 V126 V182 51.15386703960926
L126_182 V126 V182 1.5304762383650706e-12
C126_182 V126 V182 5.647034809761829e-20

R126_183 V126 V183 340.196164634479
L126_183 V126 V183 -2.243235140533117e-12
C126_183 V126 V183 -7.284453367540852e-20

R126_184 V126 V184 158.54121190123757
L126_184 V126 V184 -2.6700059148768012e-12
C126_184 V126 V184 -7.647742178321401e-20

R126_185 V126 V185 -3364.540484191202
L126_185 V126 V185 3.158222392317945e-12
C126_185 V126 V185 1.6795632912074435e-19

R126_186 V126 V186 208.7572142380074
L126_186 V126 V186 -2.0216756698936835e-12
C126_186 V126 V186 -1.424122414468794e-19

R126_187 V126 V187 2344.3294037424753
L126_187 V126 V187 1.368873802038258e-12
C126_187 V126 V187 2.838906993082656e-19

R126_188 V126 V188 -2389.1517328257273
L126_188 V126 V188 7.007095148797222e-13
C126_188 V126 V188 2.3231575794287634e-19

R126_189 V126 V189 -135.40642650746634
L126_189 V126 V189 -9.734337517566275e-12
C126_189 V126 V189 -4.858366046347388e-21

R126_190 V126 V190 -126.67329068943496
L126_190 V126 V190 2.130753612583755e-11
C126_190 V126 V190 4.3489401506467115e-20

R126_191 V126 V191 -607.4109744239415
L126_191 V126 V191 1.5949611655358128e-12
C126_191 V126 V191 -7.198074469282867e-20

R126_192 V126 V192 -166.75256437058988
L126_192 V126 V192 -2.307067123730741e-12
C126_192 V126 V192 -1.3637258784485167e-19

R126_193 V126 V193 -858.339104446528
L126_193 V126 V193 -5.138578158117977e-12
C126_193 V126 V193 -6.903959200911063e-20

R126_194 V126 V194 201.48637257147143
L126_194 V126 V194 -3.0154047289601237e-12
C126_194 V126 V194 -2.6910465807862e-19

R126_195 V126 V195 462.3228569769702
L126_195 V126 V195 -1.2139803334704216e-12
C126_195 V126 V195 9.107494072771592e-21

R126_196 V126 V196 224.4877877438602
L126_196 V126 V196 -1.5652389891023257e-11
C126_196 V126 V196 1.6414881944412775e-19

R126_197 V126 V197 664.8055173289183
L126_197 V126 V197 2.3241656734131778e-11
C126_197 V126 V197 1.6918237496633308e-20

R126_198 V126 V198 88.2921827502702
L126_198 V126 V198 -9.852116297498432e-12
C126_198 V126 V198 7.766785624780591e-22

R126_199 V126 V199 275.6506645546702
L126_199 V126 V199 2.314715054973522e-11
C126_199 V126 V199 1.1027615026475115e-19

R126_200 V126 V200 -366.2052850457733
L126_200 V126 V200 1.3089290728882135e-11
C126_200 V126 V200 9.494126453187816e-21

R127_127 V127 0 -39.617289994007564
L127_127 V127 0 6.337671901869269e-13
C127_127 V127 0 1.0802916851713056e-18

R127_128 V127 V128 -141.39186708655654
L127_128 V127 V128 1.2189600078691894e-12
C127_128 V127 V128 3.9869514531597026e-19

R127_129 V127 V129 -200.20349830795175
L127_129 V127 V129 -1.0174135409444482e-11
C127_129 V127 V129 -7.133211254409986e-20

R127_130 V127 V130 123.28858138803497
L127_130 V127 V130 3.5412873977494163e-12
C127_130 V127 V130 1.1023710375657782e-19

R127_131 V127 V131 27.134457284459362
L127_131 V127 V131 8.26630298916312e-13
C127_131 V127 V131 1.5513423930980918e-19

R127_132 V127 V132 72.79238364302462
L127_132 V127 V132 9.781405397228729e-11
C127_132 V127 V132 4.8985450758706025e-20

R127_133 V127 V133 9784.154298662463
L127_133 V127 V133 5.053259394220116e-12
C127_133 V127 V133 2.5347369144550956e-19

R127_134 V127 V134 98.860482253148
L127_134 V127 V134 2.9572598802158194e-11
C127_134 V127 V134 -6.288461241317846e-20

R127_135 V127 V135 287.24275309937144
L127_135 V127 V135 5.271889497860991e-13
C127_135 V127 V135 1.2965869714610014e-18

R127_136 V127 V136 66.5219258854988
L127_136 V127 V136 -1.1429710552120611e-12
C127_136 V127 V136 -7.510192830260386e-19

R127_137 V127 V137 133.0660068449556
L127_137 V127 V137 -2.0021137449075165e-11
C127_137 V127 V137 -2.357508176143692e-20

R127_138 V127 V138 -66.54572022316539
L127_138 V127 V138 -1.0330899635870809e-11
C127_138 V127 V138 7.586262755217055e-20

R127_139 V127 V139 -53.404682013479444
L127_139 V127 V139 -3.454536145280289e-13
C127_139 V127 V139 -1.5745564172155668e-18

R127_140 V127 V140 -30.722441022933193
L127_140 V127 V140 1.2349680807891217e-12
C127_140 V127 V140 9.430115177344545e-19

R127_141 V127 V141 368.38544770692636
L127_141 V127 V141 -1.4488852248786558e-11
C127_141 V127 V141 -2.050970359192253e-19

R127_142 V127 V142 -69.95138880550057
L127_142 V127 V142 -4.655504586593941e-12
C127_142 V127 V142 2.6585287545348927e-21

R127_143 V127 V143 197.52504094247823
L127_143 V127 V143 1.758426409878315e-12
C127_143 V127 V143 1.6026238771288912e-19

R127_144 V127 V144 194.84615806894953
L127_144 V127 V144 -1.0900434795167242e-11
C127_144 V127 V144 -2.582578715797602e-19

R127_145 V127 V145 -89.72641844596487
L127_145 V127 V145 2.07167056929442e-11
C127_145 V127 V145 4.3133431532433023e-20

R127_146 V127 V146 35.62951768489949
L127_146 V127 V146 2.2901273263044276e-12
C127_146 V127 V146 -4.123270594383672e-20

R127_147 V127 V147 -471.94626907229286
L127_147 V127 V147 1.4654623091249775e-12
C127_147 V127 V147 7.089619839904791e-19

R127_148 V127 V148 76.25291975339746
L127_148 V127 V148 -9.62390755688359e-13
C127_148 V127 V148 -4.958702077531859e-19

R127_149 V127 V149 186.38858760437336
L127_149 V127 V149 -9.833006445914326e-12
C127_149 V127 V149 7.473372341901863e-20

R127_150 V127 V150 66.06652231902179
L127_150 V127 V150 1.598142582294004e-11
C127_150 V127 V150 -2.362920916166292e-19

R127_151 V127 V151 109.45625325058701
L127_151 V127 V151 -4.390143645808968e-12
C127_151 V127 V151 -3.211896343040448e-19

R127_152 V127 V152 -107.46855294997165
L127_152 V127 V152 1.2376416935832138e-12
C127_152 V127 V152 2.410784907067242e-19

R127_153 V127 V153 176.56614476562527
L127_153 V127 V153 2.5032217445395386e-12
C127_153 V127 V153 1.6591173010515026e-19

R127_154 V127 V154 -47.584076724798344
L127_154 V127 V154 4.012727655281272e-11
C127_154 V127 V154 2.1324369167158424e-19

R127_155 V127 V155 -69.94069237600839
L127_155 V127 V155 -9.715743370107162e-13
C127_155 V127 V155 -3.8504228782656676e-19

R127_156 V127 V156 1487.826113942877
L127_156 V127 V156 -1.6666971037776474e-11
C127_156 V127 V156 4.728680701697354e-19

R127_157 V127 V157 -175.04602051484827
L127_157 V127 V157 -1.852950474734835e-12
C127_157 V127 V157 -3.1074273064033595e-19

R127_158 V127 V158 303.05783006126376
L127_158 V127 V158 -5.859364763747485e-12
C127_158 V127 V158 -5.724947890223885e-20

R127_159 V127 V159 252.10025558241324
L127_159 V127 V159 7.379901969519923e-13
C127_159 V127 V159 6.508617227084339e-19

R127_160 V127 V160 118.53373633458344
L127_160 V127 V160 -5.845807442584866e-12
C127_160 V127 V160 -3.554295876333978e-19

R127_161 V127 V161 -129.41766850375973
L127_161 V127 V161 -1.1223274079805306e-09
C127_161 V127 V161 -6.518055285196213e-20

R127_162 V127 V162 90.04948506755568
L127_162 V127 V162 1.645354962695755e-11
C127_162 V127 V162 -4.2325294681573357e-20

R127_163 V127 V163 -887.9574748878805
L127_163 V127 V163 -3.1489132565022136e-12
C127_163 V127 V163 -3.7686231277342654e-19

R127_164 V127 V164 -184.65334885588692
L127_164 V127 V164 -9.461798568933578e-12
C127_164 V127 V164 1.30078729244776e-19

R127_165 V127 V165 96.05012884483706
L127_165 V127 V165 4.540190197144583e-12
C127_165 V127 V165 1.6648859775572876e-19

R127_166 V127 V166 -228.680222936789
L127_166 V127 V166 -8.878253451591162e-12
C127_166 V127 V166 -6.804853005228374e-20

R127_167 V127 V167 64.3559369332534
L127_167 V127 V167 -9.712343782817491e-12
C127_167 V127 V167 -7.02699695117596e-20

R127_168 V127 V168 -193.75719965238315
L127_168 V127 V168 5.261397179990002e-12
C127_168 V127 V168 -1.2263405819087117e-19

R127_169 V127 V169 96.30837351360698
L127_169 V127 V169 2.2037243441958424e-12
C127_169 V127 V169 1.0643176997192898e-19

R127_170 V127 V170 834.6529996844494
L127_170 V127 V170 2.9284469551457863e-12
C127_170 V127 V170 8.663635136897274e-20

R127_171 V127 V171 -60.519970914402
L127_171 V127 V171 1.994441761101301e-12
C127_171 V127 V171 3.465555645993075e-19

R127_172 V127 V172 168.96934158000036
L127_172 V127 V172 -5.192867933495814e-12
C127_172 V127 V172 6.065685108881838e-20

R127_173 V127 V173 -67.17034439560638
L127_173 V127 V173 -2.1658312999578003e-12
C127_173 V127 V173 -1.2924142510265957e-19

R127_174 V127 V174 178.47281175662997
L127_174 V127 V174 -9.30593212536534e-12
C127_174 V127 V174 -1.5756502124629633e-20

R127_175 V127 V175 385.12856845235007
L127_175 V127 V175 -9.479984494267137e-13
C127_175 V127 V175 -4.983302765060716e-19

R127_176 V127 V176 -264.4498169076309
L127_176 V127 V176 1.9457476897986228e-12
C127_176 V127 V176 4.570480865316877e-19

R127_177 V127 V177 473.55805972536353
L127_177 V127 V177 -6.20380168322089e-11
C127_177 V127 V177 -1.0070070427083145e-21

R127_178 V127 V178 -143.43447078118587
L127_178 V127 V178 -5.853860489280328e-12
C127_178 V127 V178 -5.836854310237774e-20

R127_179 V127 V179 85.12733678809056
L127_179 V127 V179 2.184543571039977e-12
C127_179 V127 V179 2.176184880706395e-19

R127_180 V127 V180 -194.4248526333894
L127_180 V127 V180 -2.2590468185193016e-12
C127_180 V127 V180 -3.8485873937575954e-19

R127_181 V127 V181 136.95529315671055
L127_181 V127 V181 -2.8087093502097707e-11
C127_181 V127 V181 -5.175772051703554e-20

R127_182 V127 V182 230.8938322041279
L127_182 V127 V182 -7.897338869188694e-11
C127_182 V127 V182 -1.266433687361719e-20

R127_183 V127 V183 -99.66345440164037
L127_183 V127 V183 3.2976406413622566e-12
C127_183 V127 V183 -1.0822747490750702e-19

R127_184 V127 V184 222.8492671655604
L127_184 V127 V184 2.0013333922747986e-11
C127_184 V127 V184 1.0534640265366013e-19

R127_185 V127 V185 -184.83926557352743
L127_185 V127 V185 2.0670584692478553e-11
C127_185 V127 V185 3.1863581928332866e-20

R127_186 V127 V186 149.68739769425414
L127_186 V127 V186 3.5198464961556016e-11
C127_186 V127 V186 1.0832651030209691e-19

R127_187 V127 V187 -394.79590936013955
L127_187 V127 V187 -7.277454570103364e-13
C127_187 V127 V187 -3.1120932271160644e-19

R127_188 V127 V188 -389.3263822362544
L127_188 V127 V188 1.0835627664840672e-12
C127_188 V127 V188 1.6320629658843454e-19

R127_189 V127 V189 1851.7127480240124
L127_189 V127 V189 4.1450717070481435e-12
C127_189 V127 V189 1.4365558614082334e-19

R127_190 V127 V190 -4822.4428920872615
L127_190 V127 V190 -9.677092511694093e-11
C127_190 V127 V190 -1.0101940897404994e-19

R127_191 V127 V191 104.9750014218889
L127_191 V127 V191 1.0201526780132023e-12
C127_191 V127 V191 6.045286521174138e-19

R127_192 V127 V192 -424.0903950805357
L127_192 V127 V192 -9.790852786133973e-13
C127_192 V127 V192 -2.3369082074750337e-19

R127_193 V127 V193 444.1230020403174
L127_193 V127 V193 -4.8677837357661315e-12
C127_193 V127 V193 -1.0378220858806573e-19

R127_194 V127 V194 14667.229092710397
L127_194 V127 V194 -1.0207864377505456e-11
C127_194 V127 V194 -1.060227972967333e-20

R127_195 V127 V195 -105.87600579735144
L127_195 V127 V195 -8.839329014342164e-13
C127_195 V127 V195 -1.0599759275649912e-18

R127_196 V127 V196 160.01713153211162
L127_196 V127 V196 6.713525791682208e-13
C127_196 V127 V196 7.210582835623236e-19

R127_197 V127 V197 -292.2452507629897
L127_197 V127 V197 -4.98682961335473e-12
C127_197 V127 V197 -8.610259017668004e-20

R127_198 V127 V198 208.30929206279743
L127_198 V127 V198 -9.384637058175605e-12
C127_198 V127 V198 -6.79079610614696e-20

R127_199 V127 V199 639.8482078252437
L127_199 V127 V199 -1.558976725787775e-11
C127_199 V127 V199 9.371033502978435e-21

R127_200 V127 V200 -216.78641505445177
L127_200 V127 V200 -2.0598820694102716e-12
C127_200 V127 V200 -3.406114118809342e-19

R128_128 V128 0 -42.30896929870311
L128_128 V128 0 -3.8897769376117623e-13
C128_128 V128 0 -2.5872471691007567e-19

R128_129 V128 V129 -119.03670605425316
L128_129 V128 V129 -3.802625989809468e-12
C128_129 V128 V129 -9.810348478316107e-20

R128_130 V128 V130 323.7619305439349
L128_130 V128 V130 8.073555169782462e-12
C128_130 V128 V130 1.7606553268998883e-19

R128_131 V128 V131 110.00851486201562
L128_131 V128 V131 -2.1937901141401705e-12
C128_131 V128 V131 -1.4012427057087031e-19

R128_132 V128 V132 21.50039209961162
L128_132 V128 V132 1.6695503516108616e-12
C128_132 V128 V132 -9.859464173333738e-20

R128_133 V128 V133 732.4953624075465
L128_133 V128 V133 1.8914124700743583e-11
C128_133 V128 V133 9.457424272794125e-20

R128_134 V128 V134 76.7665958264411
L128_134 V128 V134 -3.492249900456881e-12
C128_134 V128 V134 -3.64736705262549e-19

R128_135 V128 V135 142.57990442315386
L128_135 V128 V135 -1.93579180603099e-12
C128_135 V128 V135 -4.822823179296237e-19

R128_136 V128 V136 83.8680557740475
L128_136 V128 V136 6.214309080925293e-13
C128_136 V128 V136 7.303675634371728e-19

R128_137 V128 V137 116.05165145483573
L128_137 V128 V137 2.4147275454485085e-12
C128_137 V128 V137 1.5610864970585538e-19

R128_138 V128 V138 -65.0258485482097
L128_138 V128 V138 4.175731550144282e-12
C128_138 V128 V138 1.9988837353359394e-19

R128_139 V128 V139 -54.525330496007044
L128_139 V128 V139 1.1658108369211365e-12
C128_139 V128 V139 7.430446425630889e-19

R128_140 V128 V140 -27.65934212769015
L128_140 V128 V140 -5.80388780085303e-13
C128_140 V128 V140 -6.691508099817352e-19

R128_141 V128 V141 501.1615944761167
L128_141 V128 V141 -2.7464631164199826e-11
C128_141 V128 V141 -2.424922143546338e-19

R128_142 V128 V142 -54.106860769917894
L128_142 V128 V142 3.4594987943865886e-11
C128_142 V128 V142 7.860272138816145e-20

R128_143 V128 V143 160.0049707546221
L128_143 V128 V143 -1.8610753936806025e-11
C128_143 V128 V143 -1.9006985973419678e-19

R128_144 V128 V144 199.9413647792908
L128_144 V128 V144 4.918269256713668e-12
C128_144 V128 V144 2.6221667297158126e-20

R128_145 V128 V145 -79.26527218672625
L128_145 V128 V145 -2.7279280098252906e-12
C128_145 V128 V145 -9.660152442059378e-20

R128_146 V128 V146 30.2520260402732
L128_146 V128 V146 -1.467016302277889e-11
C128_146 V128 V146 -7.67915706218763e-20

R128_147 V128 V147 238.2493286895974
L128_147 V128 V147 -1.0398461081561213e-11
C128_147 V128 V147 -2.8720041318085165e-19

R128_148 V128 V148 146.6404025670142
L128_148 V128 V148 8.488638282974419e-13
C128_148 V128 V148 3.3941652389552197e-19

R128_149 V128 V149 147.22241390184175
L128_149 V128 V149 6.738309294036644e-12
C128_149 V128 V149 3.558366464540604e-19

R128_150 V128 V150 63.0993326907888
L128_150 V128 V150 2.4956852983868814e-12
C128_150 V128 V150 -1.6961148289800317e-19

R128_151 V128 V151 -352.0760901888248
L128_151 V128 V151 -3.63380601853293e-12
C128_151 V128 V151 1.664964301210079e-19

R128_152 V128 V152 -304.9751261977915
L128_152 V128 V152 -9.78312958754449e-13
C128_152 V128 V152 -1.4687600032957255e-19

R128_153 V128 V153 149.73363906722267
L128_153 V128 V153 -2.3102665902516397e-11
C128_153 V128 V153 7.49814705336673e-21

R128_154 V128 V154 -43.5636865649256
L128_154 V128 V154 -2.0284723582799393e-12
C128_154 V128 V154 1.8375358658933058e-19

R128_155 V128 V155 -112.19197032630778
L128_155 V128 V155 4.129233810377706e-12
C128_155 V128 V155 2.7102092455401416e-19

R128_156 V128 V156 214.3442880869593
L128_156 V128 V156 1.5949575965073214e-11
C128_156 V128 V156 -2.5620241941926337e-19

R128_157 V128 V157 -120.30028892887701
L128_157 V128 V157 1.126033939625993e-11
C128_157 V128 V157 -2.189504843308975e-19

R128_158 V128 V158 3213.480929592215
L128_158 V128 V158 9.168306247542881e-12
C128_158 V128 V158 -3.2100381910407155e-20

R128_159 V128 V159 68.0828455765788
L128_159 V128 V159 -5.284163620491029e-12
C128_159 V128 V159 -2.5167173466896907e-19

R128_160 V128 V160 -432.58988075113916
L128_160 V128 V160 1.4439015396601876e-12
C128_160 V128 V160 3.656202477399354e-19

R128_161 V128 V161 -104.88952298975501
L128_161 V128 V161 -1.7067736538598052e-12
C128_161 V128 V161 -5.612217331504165e-20

R128_162 V128 V162 80.10419660241895
L128_162 V128 V162 -6.223357374734035e-11
C128_162 V128 V162 3.8575039040510355e-20

R128_163 V128 V163 -251.24460155384986
L128_163 V128 V163 1.4284542472220386e-11
C128_163 V128 V163 9.057936371265931e-20

R128_164 V128 V164 -337.2962360621308
L128_164 V128 V164 -5.447553997015347e-12
C128_164 V128 V164 -1.898641988879373e-19

R128_165 V128 V165 80.92341549721986
L128_165 V128 V165 3.0398686151139744e-12
C128_165 V128 V165 1.4831131566778378e-19

R128_166 V128 V166 -338.06495268270857
L128_166 V128 V166 9.596802216263082e-12
C128_166 V128 V166 2.750833597556619e-20

R128_167 V128 V167 -709.2003584512672
L128_167 V128 V167 -5.541516343303741e-12
C128_167 V128 V167 -8.001592919737698e-20

R128_168 V128 V168 82.44764219516954
L128_168 V128 V168 -2.117078192314731e-12
C128_168 V128 V168 -1.2099200697804149e-19

R128_169 V128 V169 90.62393628421925
L128_169 V128 V169 1.884194140717271e-12
C128_169 V128 V169 9.743590565814235e-20

R128_170 V128 V170 5905.100996970142
L128_170 V128 V170 -1.280107495589979e-11
C128_170 V128 V170 5.602387524153961e-20

R128_171 V128 V171 590.5544811928996
L128_171 V128 V171 -6.0311156053345824e-12
C128_171 V128 V171 6.438548932880685e-20

R128_172 V128 V172 -63.20905223353064
L128_172 V128 V172 1.5081631297160863e-12
C128_172 V128 V172 1.951090289016816e-19

R128_173 V128 V173 -51.55270287790765
L128_173 V128 V173 -1.9177124266063093e-12
C128_173 V128 V173 -9.196472673082381e-20

R128_174 V128 V174 144.75116832603842
L128_174 V128 V174 5.092433239326998e-12
C128_174 V128 V174 -7.742225296954156e-20

R128_175 V128 V175 1565.9092700932754
L128_175 V128 V175 1.5070220410275004e-12
C128_175 V128 V175 2.487020196551764e-19

R128_176 V128 V176 -369.0067341171463
L128_176 V128 V176 -1.8438879717148374e-12
C128_176 V128 V176 -2.89125805965931e-19

R128_177 V128 V177 512.9212566940295
L128_177 V128 V177 -1.1524722628613116e-11
C128_177 V128 V177 3.1691575341136347e-20

R128_178 V128 V178 -95.19245837403069
L128_178 V128 V178 -1.6755012821738738e-11
C128_178 V128 V178 -2.5017800710988155e-20

R128_179 V128 V179 -152.30673029343424
L128_179 V128 V179 -1.8455788441227737e-11
C128_179 V128 V179 -2.348085574495832e-19

R128_180 V128 V180 38.93857330361097
L128_180 V128 V180 1.479349079037677e-12
C128_180 V128 V180 1.7220025901121798e-19

R128_181 V128 V181 113.64421056001065
L128_181 V128 V181 1.892817928128103e-11
C128_181 V128 V181 -1.0362773995244071e-19

R128_182 V128 V182 278.05712223940714
L128_182 V128 V182 1.6362784248944135e-11
C128_182 V128 V182 1.1516145457690169e-19

R128_183 V128 V183 213.01982714154045
L128_183 V128 V183 1.0348991309687158e-11
C128_183 V128 V183 4.6646854481004053e-20

R128_184 V128 V184 -56.30230954091679
L128_184 V128 V184 3.754059417913909e-12
C128_184 V128 V184 -5.410043377989667e-20

R128_185 V128 V185 -116.88443089855942
L128_185 V128 V185 -1.8056039847227428e-10
C128_185 V128 V185 4.3557026472822043e-20

R128_186 V128 V186 128.3697505231128
L128_186 V128 V186 3.9523283492549056e-12
C128_186 V128 V186 -7.412567109230543e-20

R128_187 V128 V187 607.9705046773671
L128_187 V128 V187 1.8335010039349454e-12
C128_187 V128 V187 2.1563566687076005e-19

R128_188 V128 V188 -112.26814075108308
L128_188 V128 V188 -5.912657904608455e-13
C128_188 V128 V188 -1.3686353691818726e-19

R128_189 V128 V189 1186.5838140692015
L128_189 V128 V189 1.9021353784449205e-12
C128_189 V128 V189 1.7205216268258918e-19

R128_190 V128 V190 -664.1581296168922
L128_190 V128 V190 -1.047092125318409e-11
C128_190 V128 V190 -9.46160271923848e-20

R128_191 V128 V191 -325.2919195712474
L128_191 V128 V191 -1.5826275371105259e-12
C128_191 V128 V191 -1.5768501443473062e-19

R128_192 V128 V192 89.0135634161017
L128_192 V128 V192 8.017602958087715e-13
C128_192 V128 V192 4.103492439376356e-19

R128_193 V128 V193 163.3248908123778
L128_193 V128 V193 -1.3592965003254304e-11
C128_193 V128 V193 -2.7193649557686495e-20

R128_194 V128 V194 -11565.982347908935
L128_194 V128 V194 2.153183477672629e-12
C128_194 V128 V194 1.4748181118375005e-19

R128_195 V128 V195 994.9125486286285
L128_195 V128 V195 1.2504461753737992e-12
C128_195 V128 V195 3.172776017537849e-19

R128_196 V128 V196 -145.94758047935943
L128_196 V128 V196 -8.571150297231895e-13
C128_196 V128 V196 -7.929637604258085e-19

R128_197 V128 V197 -164.86394884323283
L128_197 V128 V197 -2.5479160792201346e-12
C128_197 V128 V197 -1.6419261816049867e-19

R128_198 V128 V198 181.15558775859256
L128_198 V128 V198 -1.3790794903579367e-11
C128_198 V128 V198 8.537261499445897e-20

R128_199 V128 V199 199.61753694507198
L128_199 V128 V199 -4.405217068304744e-12
C128_199 V128 V199 -1.1718967472827853e-19

R128_200 V128 V200 -123.8343383837336
L128_200 V128 V200 7.458170761497646e-12
C128_200 V128 V200 1.2505909193278322e-19

R129_129 V129 0 -31.226098970376533
L129_129 V129 0 1.403758828071282e-11
C129_129 V129 0 2.0532242810925286e-18

R129_130 V129 V130 192.5527119181372
L129_130 V129 V130 1.10511046992676e-12
C129_130 V129 V130 4.474512957954117e-19

R129_131 V129 V131 118.08294767395206
L129_131 V129 V131 3.650649127948115e-12
C129_131 V129 V131 1.9970256403819642e-19

R129_132 V129 V132 61.36433600606519
L129_132 V129 V132 1.6324001416661829e-12
C129_132 V129 V132 3.4703071382698534e-19

R129_133 V129 V133 -2046.5770357298081
L129_133 V129 V133 9.201392943593404e-13
C129_133 V129 V133 8.663012730426648e-19

R129_134 V129 V134 83.09964899412509
L129_134 V129 V134 -1.3470285892802225e-12
C129_134 V129 V134 -4.952567853572031e-19

R129_135 V129 V135 103.72077687555014
L129_135 V129 V135 3.4777252399357473e-12
C129_135 V129 V135 -1.8322682290010068e-20

R129_136 V129 V136 95.15080707962763
L129_136 V129 V136 4.806767283753097e-12
C129_136 V129 V136 -1.9447615159831736e-19

R129_137 V129 V137 27.388242639692667
L129_137 V129 V137 9.554929014015776e-13
C129_137 V129 V137 2.7416230954053897e-19

R129_138 V129 V138 -118.43448965098271
L129_138 V129 V138 4.316132822094952e-12
C129_138 V129 V138 2.010046143576764e-19

R129_139 V129 V139 -77.66796371910529
L129_139 V129 V139 -1.784875282539067e-11
C129_139 V129 V139 2.2919139419330926e-19

R129_140 V129 V140 -68.23507733725042
L129_140 V129 V140 -2.3275249757425164e-12
C129_140 V129 V140 1.311112832778709e-19

R129_141 V129 V141 316.05194295189926
L129_141 V129 V141 -9.10678328188867e-13
C129_141 V129 V141 -7.426051626946016e-19

R129_142 V129 V142 -54.38581298263327
L129_142 V129 V142 2.2116253886357478e-12
C129_142 V129 V142 1.7952711475657912e-19

R129_143 V129 V143 -100.7992716274945
L129_143 V129 V143 -1.2997809799009459e-12
C129_143 V129 V143 -3.5933767469957465e-19

R129_144 V129 V144 -67.84504189432302
L129_144 V129 V144 -3.540860485282794e-12
C129_144 V129 V144 -5.510934498634505e-20

R129_145 V129 V145 -21.882405339344185
L129_145 V129 V145 -2.4335123164674098e-12
C129_145 V129 V145 -7.224623242146168e-21

R129_146 V129 V146 -130.83451074050603
L129_146 V129 V146 -1.0642664596752928e-12
C129_146 V129 V146 -1.1113787857267702e-19

R129_147 V129 V147 -842.9979635047276
L129_147 V129 V147 3.863363048763033e-12
C129_147 V129 V147 -8.707383726588459e-20

R129_148 V129 V148 105.29023454459667
L129_148 V129 V148 4.536071011236062e-11
C129_148 V129 V148 -1.2553366054253956e-19

R129_149 V129 V149 341.29553324378105
L129_149 V129 V149 5.853723077928293e-13
C129_149 V129 V149 1.0817078974983746e-18

R129_150 V129 V150 21.27425271390403
L129_150 V129 V150 1.4817755110867666e-12
C129_150 V129 V150 -6.091926745613767e-19

R129_151 V129 V151 41.39771356160393
L129_151 V129 V151 1.5831948157684224e-12
C129_151 V129 V151 3.098962728640945e-19

R129_152 V129 V152 183.8663847363587
L129_152 V129 V152 4.653858642759235e-12
C129_152 V129 V152 -1.5338614333858786e-20

R129_153 V129 V153 26.19378723575137
L129_153 V129 V153 2.230785381794963e-11
C129_153 V129 V153 -3.321105734912716e-19

R129_154 V129 V154 88.57017424221985
L129_154 V129 V154 4.546935557289747e-12
C129_154 V129 V154 4.735825977381773e-19

R129_155 V129 V155 -63.51424237951768
L129_155 V129 V155 3.248566052137119e-12
C129_155 V129 V155 2.6585528579235545e-19

R129_156 V129 V156 58.558976123061896
L129_156 V129 V156 4.807784894545119e-12
C129_156 V129 V156 1.8300657113184153e-19

R129_157 V129 V157 46.631627990452245
L129_157 V129 V157 -6.854413567927402e-13
C129_157 V129 V157 -1.117157427674632e-18

R129_158 V129 V158 -33.3020460061661
L129_158 V129 V158 -1.4341206417768545e-11
C129_158 V129 V158 -1.789263896296378e-20

R129_159 V129 V159 -393.3426454249712
L129_159 V129 V159 -1.7004912399898424e-12
C129_159 V129 V159 -1.6569428275963945e-19

R129_160 V129 V160 -54.32148202833177
L129_160 V129 V160 -3.849582610958036e-12
C129_160 V129 V160 4.9250697763583513e-20

R129_161 V129 V161 -34.562417686002995
L129_161 V129 V161 1.763292459470342e-11
C129_161 V129 V161 3.2617132243070227e-19

R129_162 V129 V162 -49.54132079426101
L129_162 V129 V162 -8.260564388311641e-11
C129_162 V129 V162 2.894853433928355e-20

R129_163 V129 V163 -86.82909864272976
L129_163 V129 V163 -1.5925985705199192e-12
C129_163 V129 V163 -3.2005239234723685e-19

R129_164 V129 V164 -84.25442659970363
L129_164 V129 V164 -2.1272992371998756e-12
C129_164 V129 V164 -2.4889816397608006e-20

R129_165 V129 V165 -77.55304693735042
L129_165 V129 V165 7.70070421991549e-13
C129_165 V129 V165 7.743760113883371e-19

R129_166 V129 V166 22.62237778017814
L129_166 V129 V166 1.835178415463302e-12
C129_166 V129 V166 1.9647702670871465e-20

R129_167 V129 V167 81.49081525241884
L129_167 V129 V167 2.2958409216527153e-12
C129_167 V129 V167 1.2442184777673571e-19

R129_168 V129 V168 3027.7415204915296
L129_168 V129 V168 2.17332288759735e-12
C129_168 V129 V168 -1.6342162302859342e-20

R129_169 V129 V169 36.59698003140952
L129_169 V129 V169 -2.2180894242980637e-12
C129_169 V129 V169 -5.36713466972277e-19

R129_170 V129 V170 -153.02880313560337
L129_170 V129 V170 4.741608307299829e-12
C129_170 V129 V170 3.326541333028163e-19

R129_171 V129 V171 1153.0340521129424
L129_171 V129 V171 1.0000803646690545e-12
C129_171 V129 V171 5.15038409620405e-19

R129_172 V129 V172 188.75687727952814
L129_172 V129 V172 2.0622930665725315e-12
C129_172 V129 V172 2.2709825659780445e-19

R129_173 V129 V173 -184.75256767194904
L129_173 V129 V173 -2.9556829238910366e-12
C129_173 V129 V173 -1.7999457190499379e-19

R129_174 V129 V174 -32.94914380358924
L129_174 V129 V174 -1.2084645138210634e-12
C129_174 V129 V174 -6.36899901116051e-19

R129_175 V129 V175 -391.30901456106903
L129_175 V129 V175 -1.909536458712503e-12
C129_175 V129 V175 -4.3700825465759553e-20

R129_176 V129 V176 -521.0381295321517
L129_176 V129 V176 -1.331114318513669e-12
C129_176 V129 V176 -5.2432864124159676e-20

R129_177 V129 V177 -99.8909247710029
L129_177 V129 V177 -9.836559194034119e-12
C129_177 V129 V177 1.7487666730977449e-19

R129_178 V129 V178 107.69549041137486
L129_178 V129 V178 -4.1149168647657885e-12
C129_178 V129 V178 -1.190175541145031e-19

R129_179 V129 V179 -146.95872468680744
L129_179 V129 V179 -1.581563610362292e-12
C129_179 V129 V179 -5.798738400716945e-19

R129_180 V129 V180 -423.98975451921694
L129_180 V129 V180 -3.0770385352847226e-12
C129_180 V129 V180 -3.6467141906676966e-19

R129_181 V129 V181 145.3007891646088
L129_181 V129 V181 4.466847017988523e-12
C129_181 V129 V181 1.9366271669652621e-19

R129_182 V129 V182 50.80578720631301
L129_182 V129 V182 6.937776601713079e-13
C129_182 V129 V182 4.435950920452062e-19

R129_183 V129 V183 140.56914787630666
L129_183 V129 V183 -9.575107795491021e-12
C129_183 V129 V183 -1.2649785488482132e-19

R129_184 V129 V184 1233.3171923148032
L129_184 V129 V184 5.899022054596831e-12
C129_184 V129 V184 3.9622275536923935e-20

R129_185 V129 V185 120.31732373685814
L129_185 V129 V185 2.5110724207871004e-12
C129_185 V129 V185 -1.610895485082649e-19

R129_186 V129 V186 -250.1176129570563
L129_186 V129 V186 2.124425896700164e-11
C129_186 V129 V186 2.4510394160472188e-20

R129_187 V129 V187 -309.78846934912184
L129_187 V129 V187 1.4338482587961021e-12
C129_187 V129 V187 5.566636990536738e-19

R129_188 V129 V188 -240.8615325038713
L129_188 V129 V188 1.3370387805286428e-12
C129_188 V129 V188 4.731580920862528e-19

R129_189 V129 V189 -189.00578241653272
L129_189 V129 V189 -2.710297990987892e-12
C129_189 V129 V189 2.3601045480344714e-19

R129_190 V129 V190 -107.13052518071385
L129_190 V129 V190 -2.0012734231938127e-12
C129_190 V129 V190 -3.526695139525287e-19

R129_191 V129 V191 -488.47320690146483
L129_191 V129 V191 1.6440095921839924e-12
C129_191 V129 V191 3.176195843730836e-19

R129_192 V129 V192 -1132.0659338767248
L129_192 V129 V192 -8.678764132246426e-09
C129_192 V129 V192 2.9457981901522147e-20

R129_193 V129 V193 -116.93960135528903
L129_193 V129 V193 1.5119210619032584e-11
C129_193 V129 V193 -2.638734657428076e-19

R129_194 V129 V194 101.84033736770361
L129_194 V129 V194 -3.5468743644150793e-12
C129_194 V129 V194 -3.912322819919456e-19

R129_195 V129 V195 196.204149799429
L129_195 V129 V195 -8.978956014844171e-13
C129_195 V129 V195 -6.845097678657338e-19

R129_196 V129 V196 153.09867465850795
L129_196 V129 V196 -7.378555900803359e-13
C129_196 V129 V196 -5.939689030171146e-19

R129_197 V129 V197 152.78124978045844
L129_197 V129 V197 -1.602080462421045e-12
C129_197 V129 V197 -1.755212542425578e-19

R129_198 V129 V198 71.61708500417231
L129_198 V129 V198 4.113988724800647e-12
C129_198 V129 V198 9.477401453124949e-20

R129_199 V129 V199 168.28759207665271
L129_199 V129 V199 -2.0007021092312728e-12
C129_199 V129 V199 -3.566429882010264e-19

R129_200 V129 V200 -141.1446920481126
L129_200 V129 V200 7.252878086582667e-12
C129_200 V129 V200 6.159426853372786e-20

R130_130 V130 0 47.1689897640078
L130_130 V130 0 -2.573503743126028e-13
C130_130 V130 0 -2.1535756917174188e-18

R130_131 V130 V131 -83.96351183843589
L130_131 V130 V131 -2.8052252324430804e-12
C130_131 V130 V131 -9.567622052518941e-20

R130_132 V130 V132 -106.3775398460143
L130_132 V130 V132 -1.8005607967062983e-12
C130_132 V130 V132 -3.181159338478715e-19

R130_133 V130 V133 -310.09717250495345
L130_133 V130 V133 -8.25183215574093e-13
C130_133 V130 V133 -5.864526964219315e-19

R130_134 V130 V134 -318.36794738826455
L130_134 V130 V134 1.170215170351122e-12
C130_134 V130 V134 5.740498798282385e-19

R130_135 V130 V135 -470.12998462898497
L130_135 V130 V135 -3.1935225386705488e-12
C130_135 V130 V135 -7.289753781691263e-20

R130_136 V130 V136 -132.57442766764294
L130_136 V130 V136 -2.271913170752294e-11
C130_136 V130 V136 1.2811972879027084e-19

R130_137 V130 V137 -474.2969202782012
L130_137 V130 V137 -1.377105209459568e-12
C130_137 V130 V137 -3.325706612481139e-19

R130_138 V130 V138 68.06575645182042
L130_138 V130 V138 2.021197993063109e-12
C130_138 V130 V138 -1.2596474891872998e-20

R130_139 V130 V139 79.24194183775482
L130_139 V130 V139 1.126822419483615e-11
C130_139 V130 V139 -1.0892987953803624e-19

R130_140 V130 V140 44.17164257935835
L130_140 V130 V140 3.0619868284967547e-12
C130_140 V130 V140 -1.5052924224385613e-19

R130_141 V130 V141 -226.1526446571738
L130_141 V130 V141 6.326669117427341e-13
C130_141 V130 V141 8.98929231704637e-19

R130_142 V130 V142 126635.66290754384
L130_142 V130 V142 -1.3322151802588858e-12
C130_142 V130 V142 -2.1846695897879147e-19

R130_143 V130 V143 -147.71612651305873
L130_143 V130 V143 2.1199852054508215e-12
C130_143 V130 V143 2.656414188617609e-19

R130_144 V130 V144 -126.91561317941989
L130_144 V130 V144 2.599206370903032e-11
C130_144 V130 V144 1.4099866432742606e-19

R130_145 V130 V145 1426.7922581664357
L130_145 V130 V145 1.4248779789572324e-12
C130_145 V130 V145 2.900075733989401e-19

R130_146 V130 V146 -61.75962388542308
L130_146 V130 V146 3.358096364797517e-12
C130_146 V130 V146 -3.807435474854388e-21

R130_147 V130 V147 -230.3861262343033
L130_147 V130 V147 1.2103374259603418e-11
C130_147 V130 V147 1.0047768934658574e-19

R130_148 V130 V148 -154.5427147544144
L130_148 V130 V148 2.3716698830533824e-12
C130_148 V130 V148 1.4620481681633362e-19

R130_149 V130 V149 111.34000688225885
L130_149 V130 V149 -3.9917711724288185e-13
C130_149 V130 V149 -1.2103149323889505e-18

R130_150 V130 V150 -389.9339410641924
L130_150 V130 V150 -1.2259573514110793e-11
C130_150 V130 V150 6.243618043727096e-19

R130_151 V130 V151 146.39567967026994
L130_151 V130 V151 -9.800366707369933e-12
C130_151 V130 V151 -1.3993375554722945e-19

R130_152 V130 V152 123.68204230918602
L130_152 V130 V152 -1.5667685834332934e-11
C130_152 V130 V152 5.246383278440342e-21

R130_153 V130 V153 -1043.0564577249372
L130_153 V130 V153 -3.0544206100867306e-12
C130_153 V130 V153 -1.3327175708935452e-19

R130_154 V130 V154 78.62734345717902
L130_154 V130 V154 1.9318914376000173e-11
C130_154 V130 V154 -4.599240481273765e-19

R130_155 V130 V155 -227.63894979810993
L130_155 V130 V155 -1.3344586626565887e-12
C130_155 V130 V155 -2.75727061022026e-19

R130_156 V130 V156 -424.75782713107736
L130_156 V130 V156 -4.28842294413437e-12
C130_156 V130 V156 -2.2659023657798025e-19

R130_157 V130 V157 -95.12367710094478
L130_157 V130 V157 4.702444542237546e-13
C130_157 V130 V157 1.0364754386960481e-18

R130_158 V130 V158 -113.00593098187089
L130_158 V130 V158 -6.184727557709598e-12
C130_158 V130 V158 6.669389398336874e-20

R130_159 V130 V159 -171.17540579817057
L130_159 V130 V159 -3.748334086932067e-11
C130_159 V130 V159 -1.778970952028652e-20

R130_160 V130 V160 -131.42352521490253
L130_160 V130 V160 -2.415991331718789e-12
C130_160 V130 V160 -1.261447124138778e-19

R130_161 V130 V161 105.24108333493423
L130_161 V130 V161 3.985044052976731e-12
C130_161 V130 V161 1.1714056786139058e-19

R130_162 V130 V162 713.4390464145623
L130_162 V130 V162 -1.7290744908087768e-12
C130_162 V130 V162 -1.699064204323199e-19

R130_163 V130 V163 80.83691965475207
L130_163 V130 V163 1.2639196807582213e-12
C130_163 V130 V163 2.056621413041728e-19

R130_164 V130 V164 61.22438333101342
L130_164 V130 V164 1.4870346586785559e-12
C130_164 V130 V164 5.788316364543548e-20

R130_165 V130 V165 502.07678305846684
L130_165 V130 V165 -1.0533263355479873e-12
C130_165 V130 V165 -4.467209303148188e-19

R130_166 V130 V166 100.45299530894778
L130_166 V130 V166 3.949879109692934e-12
C130_166 V130 V166 1.208976279913646e-19

R130_167 V130 V167 -476.54822594998194
L130_167 V130 V167 1.2310294602760471e-11
C130_167 V130 V167 7.49034297983607e-20

R130_168 V130 V168 -213.1794181061381
L130_168 V130 V168 6.820459756606873e-12
C130_168 V130 V168 2.2882364155036435e-19

R130_169 V130 V169 -72.49480884739154
L130_169 V130 V169 -5.4344363426415236e-12
C130_169 V130 V169 1.291110778444758e-19

R130_170 V130 V170 -61.68971889179511
L130_170 V130 V170 -3.4752143018947725e-12
C130_170 V130 V170 -2.4346148165365574e-19

R130_171 V130 V171 -87.7308291146652
L130_171 V130 V171 -7.828480217881052e-13
C130_171 V130 V171 -3.9704516703829764e-19

R130_172 V130 V172 -91.6516871156246
L130_172 V130 V172 -1.4168201242050508e-12
C130_172 V130 V172 -2.808720976401575e-19

R130_173 V130 V173 182.7140032333374
L130_173 V130 V173 1.9274700508848984e-12
C130_173 V130 V173 -5.582755582935692e-20

R130_174 V130 V174 -304.45216557298903
L130_174 V130 V174 -1.0360904958402267e-11
C130_174 V130 V174 2.818106186354436e-19

R130_175 V130 V175 227.62258866648546
L130_175 V130 V175 -1.4750017034109782e-11
C130_175 V130 V175 -1.2661381893692849e-19

R130_176 V130 V176 113.60163499982656
L130_176 V130 V176 -8.129642051337894e-12
C130_176 V130 V176 -1.7317194270184698e-19

R130_177 V130 V177 127.96652352408216
L130_177 V130 V177 -2.2054797266104346e-11
C130_177 V130 V177 -1.4138988179493122e-19

R130_178 V130 V178 58.10748521620643
L130_178 V130 V178 2.0275282583914336e-12
C130_178 V130 V178 1.4329239660059307e-19

R130_179 V130 V179 465.0055200839747
L130_179 V130 V179 8.884032466196547e-13
C130_179 V130 V179 4.367591266931701e-19

R130_180 V130 V180 170.79620056218053
L130_180 V130 V180 8.737016571966952e-13
C130_180 V130 V180 3.3926301134864933e-19

R130_181 V130 V181 -119.36786311224981
L130_181 V130 V181 4.3807435438304745e-11
C130_181 V130 V181 4.1826011952721795e-19

R130_182 V130 V182 -70.05708286630417
L130_182 V130 V182 -8.726276737959159e-13
C130_182 V130 V182 -2.9067424371133566e-19

R130_183 V130 V183 5292.9556304993475
L130_183 V130 V183 2.5456066887347983e-12
C130_183 V130 V183 1.3366223470452842e-19

R130_184 V130 V184 -190.02560171449235
L130_184 V130 V184 2.1289112433526182e-11
C130_184 V130 V184 3.369786622996333e-20

R130_185 V130 V185 -293.18845944941364
L130_185 V130 V185 6.453972828214556e-12
C130_185 V130 V185 -1.3592974895821168e-19

R130_186 V130 V186 -124.10297640623791
L130_186 V130 V186 6.1318537742843035e-12
C130_186 V130 V186 8.798715235157584e-20

R130_187 V130 V187 1581.8679392843524
L130_187 V130 V187 -1.21439869805579e-12
C130_187 V130 V187 -3.526161020467549e-19

R130_188 V130 V188 -8172.741545587896
L130_188 V130 V188 -9.448608037514605e-13
C130_188 V130 V188 -2.590731136239651e-19

R130_189 V130 V189 131.9603606242442
L130_189 V130 V189 -1.6611600583051775e-12
C130_189 V130 V189 -4.023068031870588e-19

R130_190 V130 V190 102.60002423040461
L130_190 V130 V190 7.674709276176178e-12
C130_190 V130 V190 2.673637979036597e-19

R130_191 V130 V191 -11063.278667189534
L130_191 V130 V191 -1.1104211504993417e-12
C130_191 V130 V191 -3.362381891321598e-19

R130_192 V130 V192 197.98040569617402
L130_192 V130 V192 -8.542773849773314e-12
C130_192 V130 V192 -2.7452840625953404e-19

R130_193 V130 V193 425.0683558016199
L130_193 V130 V193 3.617143520946779e-12
C130_193 V130 V193 1.8323854708317134e-19

R130_194 V130 V194 -133.1282913563867
L130_194 V130 V194 8.272163611972804e-12
C130_194 V130 V194 1.2048771723447642e-19

R130_195 V130 V195 -1848.172414770605
L130_195 V130 V195 7.369236939774379e-13
C130_195 V130 V195 5.953413612681367e-19

R130_196 V130 V196 -456.3379323030664
L130_196 V130 V196 1.0693518017941696e-12
C130_196 V130 V196 4.823013974070195e-19

R130_197 V130 V197 -224.66908965919072
L130_197 V130 V197 1.5357509895901115e-12
C130_197 V130 V197 2.9987819800932467e-19

R130_198 V130 V198 -172.05671060602984
L130_198 V130 V198 -1.057005983169482e-11
C130_198 V130 V198 -1.150355412522883e-19

R130_199 V130 V199 -2257.8513024471326
L130_199 V130 V199 2.284883429005758e-12
C130_199 V130 V199 2.0671814026937497e-19

R130_200 V130 V200 -1734.7988513156174
L130_200 V130 V200 5.9457803125867985e-12
C130_200 V130 V200 7.86583637630054e-20

R131_131 V131 0 35.28575904558404
L131_131 V131 0 -6.672597377648275e-13
C131_131 V131 0 -1.3670381935912007e-18

R131_132 V131 V132 -46.86866238525558
L131_132 V131 V132 -1.6254400084326263e-12
C131_132 V131 V132 -3.774150954861602e-19

R131_133 V131 V133 -325.3233089381065
L131_133 V131 V133 -2.9944194935616136e-12
C131_133 V131 V133 -2.5564474049381387e-19

R131_134 V131 V134 -82.49545979565634
L131_134 V131 V134 -2.9983638053093875e-12
C131_134 V131 V134 -1.6535574982461503e-19

R131_135 V131 V135 306.8810062763933
L131_135 V131 V135 5.268381183452612e-12
C131_135 V131 V135 1.5800735605900177e-19

R131_136 V131 V136 -59.382629366206906
L131_136 V131 V136 2.020130156658575e-12
C131_136 V131 V136 5.848392068841987e-19

R131_137 V131 V137 -131.46015494023274
L131_137 V131 V137 2.1866083920813484e-09
C131_137 V131 V137 6.143691815597819e-22

R131_138 V131 V138 52.12991773618466
L131_138 V131 V138 1.6297499731286806e-12
C131_138 V131 V138 2.220172170126433e-19

R131_139 V131 V139 53.986762248371015
L131_139 V131 V139 1.3734366232160716e-12
C131_139 V131 V139 1.4022612522685326e-19

R131_140 V131 V140 25.69530046902485
L131_140 V131 V140 -6.461001809526121e-12
C131_140 V131 V140 -6.501665314066218e-19

R131_141 V131 V141 -411.4674687148574
L131_141 V131 V141 3.0674879614165274e-12
C131_141 V131 V141 2.922523953982955e-19

R131_142 V131 V142 60.43613067389167
L131_142 V131 V142 3.310828199802577e-12
C131_142 V131 V142 -1.2600341599272916e-20

R131_143 V131 V143 -82.74837374863478
L131_143 V131 V143 -6.985488072787716e-12
C131_143 V131 V143 -4.390561306409957e-20

R131_144 V131 V144 -219.20063659821298
L131_144 V131 V144 1.5890112140771377e-11
C131_144 V131 V144 1.413875230389267e-19

R131_145 V131 V145 93.42804216330524
L131_145 V131 V145 5.000113832701022e-11
C131_145 V131 V145 1.672050727095301e-20

R131_146 V131 V146 -30.36198322979404
L131_146 V131 V146 -1.2203955608082375e-12
C131_146 V131 V146 -1.0524614007422119e-19

R131_147 V131 V147 113.54831030053244
L131_147 V131 V147 6.504568518680849e-12
C131_147 V131 V147 1.571289569908304e-19

R131_148 V131 V148 -53.083902137729595
L131_148 V131 V148 2.0017323119966783e-12
C131_148 V131 V148 4.1415826424223215e-19

R131_149 V131 V149 -979.1442801459852
L131_149 V131 V149 -2.2090015622143328e-12
C131_149 V131 V149 -3.3389755188644067e-19

R131_150 V131 V150 -55.66945330550671
L131_150 V131 V150 1.5349021868802742e-10
C131_150 V131 V150 1.6927253695487792e-19

R131_151 V131 V151 243.739191742408
L131_151 V131 V151 -8.22806205400918e-12
C131_151 V131 V151 -6.230127050081406e-20

R131_152 V131 V152 92.41797064624734
L131_152 V131 V152 -2.7978658341813406e-12
C131_152 V131 V152 -1.3739124964635215e-19

R131_153 V131 V153 -116.05866284674043
L131_153 V131 V153 -5.150679826837102e-12
C131_153 V131 V153 1.04250684816312e-20

R131_154 V131 V154 43.690653391651466
L131_154 V131 V154 4.632594157048264e-12
C131_154 V131 V154 -1.78650741399199e-20

R131_155 V131 V155 -168.8702796996663
L131_155 V131 V155 -2.160616138224867e-12
C131_155 V131 V155 -1.26843257027785e-19

R131_156 V131 V156 -397.39034520086057
L131_156 V131 V156 -1.361197024941386e-11
C131_156 V131 V156 -3.6240119506190464e-19

R131_157 V131 V157 2094.4111589101835
L131_157 V131 V157 1.3949761585448607e-12
C131_157 V131 V157 3.6034420315994396e-19

R131_158 V131 V158 -2177.1909002149005
L131_158 V131 V158 -4.986868695365883e-11
C131_158 V131 V158 -9.033568489104445e-20

R131_159 V131 V159 -86.57940910568385
L131_159 V131 V159 4.29163615786289e-12
C131_159 V131 V159 7.08785258229873e-20

R131_160 V131 V160 -209.86413853988313
L131_160 V131 V160 7.984315014940739e-12
C131_160 V131 V160 2.2199750718689727e-19

R131_161 V131 V161 72.0496936518526
L131_161 V131 V161 -4.187611262729035e-12
C131_161 V131 V161 -1.5301730727484476e-19

R131_162 V131 V162 -137.69181666374723
L131_162 V131 V162 -2.9742252057500333e-12
C131_162 V131 V162 -9.076179742484801e-20

R131_163 V131 V163 63.277558144099864
L131_163 V131 V163 1.028062110568109e-09
C131_163 V131 V163 -9.802312766457032e-20

R131_164 V131 V164 87.00028682355062
L131_164 V131 V164 4.166414201575635e-12
C131_164 V131 V164 -1.7516785462839768e-19

R131_165 V131 V165 -128.80328892381232
L131_165 V131 V165 -9.649443335942612e-12
C131_165 V131 V165 3.1726979562908545e-20

R131_166 V131 V166 964.8436445321234
L131_166 V131 V166 3.779503652696343e-12
C131_166 V131 V166 1.2813673742011397e-19

R131_167 V131 V167 -77.58165498029173
L131_167 V131 V167 -2.7108246716151485e-12
C131_167 V131 V167 4.437106267008973e-20

R131_168 V131 V168 -1593.8229344498623
L131_168 V131 V168 -2.144469697704896e-12
C131_168 V131 V168 8.142068536983103e-21

R131_169 V131 V169 -57.73690282793563
L131_169 V131 V169 1.494601400798545e-11
C131_169 V131 V169 2.0687744467867225e-19

R131_170 V131 V170 -159.8488643551955
L131_170 V131 V170 -2.492587412212458e-12
C131_170 V131 V170 -6.562212204137669e-20

R131_171 V131 V171 218.52050541878515
L131_171 V131 V171 6.822890891876525e-12
C131_171 V131 V171 -7.940642887585213e-20

R131_172 V131 V172 -118.65717787230194
L131_172 V131 V172 4.0951904244074785e-12
C131_172 V131 V172 8.551068314587669e-20

R131_173 V131 V173 58.49226215584518
L131_173 V131 V173 1.8971554998583104e-11
C131_173 V131 V173 -1.7855772279325726e-19

R131_174 V131 V174 -842.6433340371658
L131_174 V131 V174 7.135376808116419e-12
C131_174 V131 V174 9.498541447914316e-20

R131_175 V131 V175 892.8996559632377
L131_175 V131 V175 -6.611798970796637e-11
C131_175 V131 V175 -8.219649501590672e-20

R131_176 V131 V176 129.42635522532197
L131_176 V131 V176 -9.475468185550313e-12
C131_176 V131 V176 -3.310188603551442e-19

R131_177 V131 V177 455.7899325258878
L131_177 V131 V177 1.3360274845522037e-11
C131_177 V131 V177 2.61137651610772e-20

R131_178 V131 V178 80.87992171566458
L131_178 V131 V178 2.1764698873925407e-12
C131_178 V131 V178 -6.53180508659374e-21

R131_179 V131 V179 -83.07036512594185
L131_179 V131 V179 -3.9791929074042275e-12
C131_179 V131 V179 2.302268967800318e-19

R131_180 V131 V180 172.41476597434277
L131_180 V131 V180 2.355181785274183e-12
C131_180 V131 V180 2.8092168807055505e-19

R131_181 V131 V181 -97.37754595808028
L131_181 V131 V181 -8.045920079435936e-12
C131_181 V131 V181 8.865796746554428e-20

R131_182 V131 V182 -79.20116454718055
L131_182 V131 V182 -2.0755880650710083e-12
C131_182 V131 V182 -4.395750159709266e-20

R131_183 V131 V183 86.49081051990309
L131_183 V131 V183 1.1916473695945168e-12
C131_183 V131 V183 6.216509975423801e-20

R131_184 V131 V184 -161.45571090822466
L131_184 V131 V184 1.2379159882122066e-11
C131_184 V131 V184 1.0400263191821169e-20

R131_185 V131 V185 476.0720679857858
L131_185 V131 V185 -1.5826616105301436e-11
C131_185 V131 V185 -7.386775958605232e-20

R131_186 V131 V186 -109.68370572354318
L131_186 V131 V186 2.52259301589312e-11
C131_186 V131 V186 7.51521541072493e-20

R131_187 V131 V187 204.67052756584482
L131_187 V131 V187 -1.885549581130308e-11
C131_187 V131 V187 -2.2052720590569317e-19

R131_188 V131 V188 344.39687194092335
L131_188 V131 V188 -1.0420935412731794e-12
C131_188 V131 V188 -2.5353788029300817e-19

R131_189 V131 V189 373.9871399056197
L131_189 V131 V189 5.477828651282305e-12
C131_189 V131 V189 1.0606217375447176e-20

R131_190 V131 V190 145.39978249223412
L131_190 V131 V190 4.209124680039896e-12
C131_190 V131 V190 2.1954786569422886e-20

R131_191 V131 V191 -92.91325614148751
L131_191 V131 V191 -9.190168574494527e-13
C131_191 V131 V191 -6.899291873560689e-20

R131_192 V131 V192 221.1683462807539
L131_192 V131 V192 1.3958146636542604e-12
C131_192 V131 V192 2.3332658303159787e-19

R131_193 V131 V193 1417.7530234232447
L131_193 V131 V193 4.295441039574738e-11
C131_193 V131 V193 6.655846924072004e-20

R131_194 V131 V194 -230.13939775453812
L131_194 V131 V194 8.47661587862466e-12
C131_194 V131 V194 2.0849390905290272e-19

R131_195 V131 V195 137.60234200506545
L131_195 V131 V195 7.446656037501358e-13
C131_195 V131 V195 3.1963570683586597e-19

R131_196 V131 V196 -157.6978722847743
L131_196 V131 V196 -1.7219552928028945e-12
C131_196 V131 V196 -3.5977525471829846e-19

R131_197 V131 V197 813.1508305468599
L131_197 V131 V197 -2.278517773821656e-11
C131_197 V131 V197 -3.800330199549593e-20

R131_198 V131 V198 -117.28704524571063
L131_198 V131 V198 -6.004683051134409e-12
C131_198 V131 V198 4.8326303954336855e-20

R131_199 V131 V199 -1250.5875347123676
L131_199 V131 V199 1.565646150596577e-11
C131_199 V131 V199 -1.0400746251324173e-19

R131_200 V131 V200 192.12099416586693
L131_200 V131 V200 1.9109998209532612e-11
C131_200 V131 V200 4.612585192147007e-20

R132_132 V132 0 32.76073492183287
L132_132 V132 0 -4.719108158500524e-13
C132_132 V132 0 -2.665522402245026e-18

R132_133 V132 V133 -159.1047719513219
L132_133 V132 V133 -1.3743627314012254e-12
C132_133 V132 V133 -5.301480868353664e-19

R132_134 V132 V134 -49.992640374734464
L132_134 V132 V134 -2.7758671628583626e-12
C132_134 V132 V134 -2.1857045932304926e-19

R132_135 V132 V135 -132.51738640711645
L132_135 V132 V135 3.915726762178103e-12
C132_135 V132 V135 3.2117796169587356e-19

R132_136 V132 V136 -71.33255362624867
L132_136 V132 V136 1.437767215992992e-12
C132_136 V132 V136 1.005046432978344e-18

R132_137 V132 V137 -88.91241664543598
L132_137 V132 V137 -3.565239993851401e-12
C132_137 V132 V137 -7.542007300687287e-20

R132_138 V132 V138 38.35791641502501
L132_138 V132 V138 1.2376192571380552e-12
C132_138 V132 V138 3.757590425226975e-19

R132_139 V132 V139 36.342382174279976
L132_139 V132 V139 -4.415051559105611e-12
C132_139 V132 V139 -4.497355182742088e-19

R132_140 V132 V140 16.799672153194226
L132_140 V132 V140 1.7368455026122528e-12
C132_140 V132 V140 -7.576627551485133e-19

R132_141 V132 V141 -325.51160730921526
L132_141 V132 V141 1.2533975607209477e-12
C132_141 V132 V141 6.810569828015851e-19

R132_142 V132 V142 36.86988466326877
L132_142 V132 V142 3.053422952807489e-12
C132_142 V132 V142 -2.4251920059153502e-20

R132_143 V132 V143 -94.24484446574165
L132_143 V132 V143 3.742758028210749e-12
C132_143 V132 V143 1.7992772701811013e-19

R132_144 V132 V144 -55.32107328998116
L132_144 V132 V144 -2.361130557601047e-12
C132_144 V132 V144 4.5657994318315954e-20

R132_145 V132 V145 62.98816475868879
L132_145 V132 V145 3.337674052740203e-12
C132_145 V132 V145 8.326867347540063e-20

R132_146 V132 V146 -18.99809070537504
L132_146 V132 V146 -8.966918500733617e-13
C132_146 V132 V146 -2.245865075869814e-19

R132_147 V132 V147 -173.5955415215468
L132_147 V132 V147 3.761788370595079e-12
C132_147 V132 V147 5.372741352174188e-19

R132_148 V132 V148 -1495.3446745419935
L132_148 V132 V148 8.884916560789142e-13
C132_148 V132 V148 7.333988934176692e-19

R132_149 V132 V149 -410.3584524482983
L132_149 V132 V149 -9.254470236667278e-13
C132_149 V132 V149 -7.567473445985842e-19

R132_150 V132 V150 -42.811293040909476
L132_150 V132 V150 9.741121905510378e-12
C132_150 V132 V150 3.8505635416778557e-19

R132_151 V132 V151 135.16757953947388
L132_151 V132 V151 -7.87104568153698e-12
C132_151 V132 V151 -2.2361041387969067e-19

R132_152 V132 V152 64.29510241881547
L132_152 V132 V152 -2.257766057747978e-12
C132_152 V132 V152 -2.2285025107557964e-19

R132_153 V132 V153 -85.01473751291931
L132_153 V132 V153 -2.7294016171534525e-12
C132_153 V132 V153 -6.644144007766296e-21

R132_154 V132 V154 29.80078509469072
L132_154 V132 V154 4.200416735139246e-12
C132_154 V132 V154 -8.559233575128128e-20

R132_155 V132 V155 295.0979121548114
L132_155 V132 V155 -1.1920461731060966e-12
C132_155 V132 V155 -3.8555314115096586e-19

R132_156 V132 V156 -53.383394168291
L132_156 V132 V156 -3.328525581499098e-12
C132_156 V132 V156 -4.886150358520838e-19

R132_157 V132 V157 246.53970982675466
L132_157 V132 V157 7.961724878150651e-13
C132_157 V132 V157 7.607104056339239e-19

R132_158 V132 V158 276.2673520752617
L132_158 V132 V158 4.084705889126905e-11
C132_158 V132 V158 -1.2234423878332633e-19

R132_159 V132 V159 -57.97597166519841
L132_159 V132 V159 3.0852023647622016e-12
C132_159 V132 V159 2.0755502918812177e-19

R132_160 V132 V160 -80.74823221395536
L132_160 V132 V160 1.0029776494430057e-11
C132_160 V132 V160 2.7450765004764636e-19

R132_161 V132 V161 45.671802701997905
L132_161 V132 V161 -5.851650269246919e-12
C132_161 V132 V161 -2.559848493867709e-19

R132_162 V132 V162 -82.60264192581604
L132_162 V132 V162 -1.8147909323872674e-12
C132_162 V132 V162 -2.0489929811121389e-19

R132_163 V132 V163 69.1627177628076
L132_163 V132 V163 4.020145702594342e-12
C132_163 V132 V163 -9.002123167673893e-20

R132_164 V132 V164 34.39202242927321
L132_164 V132 V164 2.289981819777115e-12
C132_164 V132 V164 -3.4749838829389183e-19

R132_165 V132 V165 -85.03527525146762
L132_165 V132 V165 1.0281551077906632e-11
C132_165 V132 V165 9.885449535200918e-20

R132_166 V132 V166 1005.0957095601752
L132_166 V132 V166 2.1777024660095182e-12
C132_166 V132 V166 2.5657588359498876e-19

R132_167 V132 V167 -1109.1209654616866
L132_167 V132 V167 -8.383973362751272e-12
C132_167 V132 V167 -2.88207591539482e-20

R132_168 V132 V168 -50.2979549016113
L132_168 V132 V168 -1.106267806285541e-12
C132_168 V132 V168 1.5116362518319215e-19

R132_169 V132 V169 -39.65360830352126
L132_169 V132 V169 -8.090173315887078e-12
C132_169 V132 V169 3.6493859846821946e-19

R132_170 V132 V170 -134.17781219862422
L132_170 V132 V170 -2.1720162511169638e-12
C132_170 V132 V170 -9.614653243373758e-20

R132_171 V132 V171 -128.3555066242537
L132_171 V132 V171 -3.3088737721541663e-12
C132_171 V132 V171 2.468480557311921e-20

R132_172 V132 V172 128.08931857691132
L132_172 V132 V172 1.1371886580630684e-12
C132_172 V132 V172 4.053381977666203e-20

R132_173 V132 V173 33.58962502097605
L132_173 V132 V173 1.7542602867953348e-11
C132_173 V132 V173 -3.696436954388494e-19

R132_174 V132 V174 -209.003015833582
L132_174 V132 V174 -1.2309324334657541e-11
C132_174 V132 V174 1.619800157537498e-19

R132_175 V132 V175 551.8094976909588
L132_175 V132 V175 -1.0483761187502195e-11
C132_175 V132 V175 -3.0625741839833127e-19

R132_176 V132 V176 86.43964416500718
L132_176 V132 V176 -1.8060883009488081e-12
C132_176 V132 V176 -6.015938526328395e-19

R132_177 V132 V177 235.19085824292483
L132_177 V132 V177 3.99029464026971e-12
C132_177 V132 V177 3.7525499151687175e-20

R132_178 V132 V178 44.79328687255287
L132_178 V132 V178 1.2991002684296355e-12
C132_178 V132 V178 -2.831965928150736e-20

R132_179 V132 V179 152.7199877303871
L132_179 V132 V179 1.7895263256451537e-12
C132_179 V132 V179 3.7141318778380515e-19

R132_180 V132 V180 -31.718232367841143
L132_180 V132 V180 -2.7953372428558556e-12
C132_180 V132 V180 5.890892438142975e-19

R132_181 V132 V181 -58.5876543050195
L132_181 V132 V181 -1.3546440588848387e-11
C132_181 V132 V181 3.076269991475319e-19

R132_182 V132 V182 -59.59839824489549
L132_182 V132 V182 -1.3649680761942572e-12
C132_182 V132 V182 -1.0003986315871991e-19

R132_183 V132 V183 -202.97075778793854
L132_183 V132 V183 2.9056836908159553e-12
C132_183 V132 V183 1.5847977201736385e-19

R132_184 V132 V184 51.9414682312293
L132_184 V132 V184 8.831873264716144e-13
C132_184 V132 V184 -5.873039204566042e-20

R132_185 V132 V185 145.8366170876936
L132_185 V132 V185 -3.3222600999060134e-11
C132_185 V132 V185 -2.0843927757078834e-19

R132_186 V132 V186 -63.2300461982257
L132_186 V132 V186 5.607399061675291e-12
C132_186 V132 V186 1.770758936448344e-19

R132_187 V132 V187 -646.9533757364105
L132_187 V132 V187 -1.6364637495491371e-12
C132_187 V132 V187 -4.794566403804947e-19

R132_188 V132 V188 59.39713367765917
L132_188 V132 V188 -9.852951706596104e-13
C132_188 V132 V188 -3.5519816493796096e-19

R132_189 V132 V189 304.5867592316803
L132_189 V132 V189 -1.1790740056138402e-11
C132_189 V132 V189 -8.80093809911804e-20

R132_190 V132 V190 78.37644987610267
L132_190 V132 V190 2.7359493730558193e-12
C132_190 V132 V190 7.823714198290945e-20

R132_191 V132 V191 189.9876763951103
L132_191 V132 V191 -2.5534926461186046e-12
C132_191 V132 V191 -6.2555672691376576e-21

R132_192 V132 V192 -66.1049395847597
L132_192 V132 V192 -5.194234661210606e-12
C132_192 V132 V192 2.313392610671915e-19

R132_193 V132 V193 -204.80065027597678
L132_193 V132 V193 3.689708534422673e-11
C132_193 V132 V193 1.3756471804742584e-19

R132_194 V132 V194 -182.07155801510842
L132_194 V132 V194 -1.8123718767980603e-11
C132_194 V132 V194 3.6517403886414497e-19

R132_195 V132 V195 -458.2744059405611
L132_195 V132 V195 1.3729133656407042e-12
C132_195 V132 V195 3.2814344481371115e-19

R132_196 V132 V196 136.2588348563818
L132_196 V132 V196 1.6048759195258998e-12
C132_196 V132 V196 -3.3668108373810397e-19

R132_197 V132 V197 250.08867063778322
L132_197 V132 V197 9.196731969583592e-12
C132_197 V132 V197 -9.352859156929478e-21

R132_198 V132 V198 -84.35462449334035
L132_198 V132 V198 -3.881100900342393e-12
C132_198 V132 V198 4.293164109146914e-20

R132_199 V132 V199 -220.76649621860628
L132_199 V132 V199 -3.107860821290821e-11
C132_199 V132 V199 -4.996272651196665e-20

R132_200 V132 V200 88.25425721891138
L132_200 V132 V200 5.683061946144973e-12
C132_200 V132 V200 1.723616266288045e-20

R133_133 V133 0 403.68190577981306
L133_133 V133 0 -2.0905452924479055e-13
C133_133 V133 0 -3.269482824923427e-18

R133_134 V133 V134 1272.196249576481
L133_134 V133 V134 1.1694208318278662e-12
C133_134 V133 V134 4.606854362007905e-19

R133_135 V133 V135 270.7553402024991
L133_135 V133 V135 -2.5296592965112857e-12
C133_135 V133 V135 -2.778402523666457e-19

R133_136 V133 V136 291.20093088525294
L133_136 V133 V136 1.732775216914988e-11
C133_136 V133 V136 2.5284236582150296e-19

R133_137 V133 V137 114.83087949553274
L133_137 V133 V137 -2.2213645562935806e-12
C133_137 V133 V137 -1.944585814851441e-19

R133_138 V133 V138 547.4246894988052
L133_138 V133 V138 -1.4641448895348977e-11
C133_138 V133 V138 -1.4676642269535928e-19

R133_139 V133 V139 -511.2584246171133
L133_139 V133 V139 3.844436345366724e-12
C133_139 V133 V139 1.889965338534969e-19

R133_140 V133 V140 1873.1550962098265
L133_140 V133 V140 4.438898678910064e-12
C133_140 V133 V140 -2.0875368063813172e-19

R133_141 V133 V141 531.0777859630927
L133_141 V133 V141 4.58004858491668e-13
C133_141 V133 V141 1.3617335292992703e-18

R133_142 V133 V142 -215.78234421724716
L133_142 V133 V142 -1.1095935484606237e-12
C133_142 V133 V142 -1.3634248435703229e-19

R133_143 V133 V143 -228.5379231586966
L133_143 V133 V143 4.842385657557464e-12
C133_143 V133 V143 2.1415059880657667e-19

R133_144 V133 V144 -160.05038095406778
L133_144 V133 V144 -9.336789214557828e-12
C133_144 V133 V144 1.4955987320040636e-19

R133_145 V133 V145 -117.3108784633823
L133_145 V133 V145 2.271146326359436e-12
C133_145 V133 V145 2.6392044220252245e-20

R133_146 V133 V146 -541.8913317111563
L133_146 V133 V146 1.0839422997165445e-12
C133_146 V133 V146 2.911991992492832e-20

R133_147 V133 V147 355.25803458371877
L133_147 V133 V147 6.994589339073143e-12
C133_147 V133 V147 -5.206886795175854e-21

R133_148 V133 V148 201.3405949988091
L133_148 V133 V148 1.786922308305181e-12
C133_148 V133 V148 2.686215110724893e-19

R133_149 V133 V149 450.4394472439681
L133_149 V133 V149 -4.183130520542839e-13
C133_149 V133 V149 -1.2027883764778182e-18

R133_150 V133 V150 104.38659757367584
L133_150 V133 V150 1.782722455411696e-11
C133_150 V133 V150 7.319490950041724e-19

R133_151 V133 V151 130.16800496295662
L133_151 V133 V151 2.4902543250832844e-11
C133_151 V133 V151 -1.176011177112945e-19

R133_152 V133 V152 214.35818254217713
L133_152 V133 V152 -1.1775796062681569e-11
C133_152 V133 V152 -7.166011389965014e-20

R133_153 V133 V153 133.90506749073054
L133_153 V133 V153 -3.435354620424243e-12
C133_153 V133 V153 -5.880909007655202e-20

R133_154 V133 V154 -625.6506303498178
L133_154 V133 V154 -2.732209679047239e-12
C133_154 V133 V154 -5.913628439166277e-19

R133_155 V133 V155 -93.46317587123632
L133_155 V133 V155 -1.7234864991997282e-12
C133_155 V133 V155 -2.0476502887662555e-19

R133_156 V133 V156 -225.62196324246065
L133_156 V133 V156 -3.928659760700099e-12
C133_156 V133 V156 -3.099532191023499e-19

R133_157 V133 V157 -397.9205765368993
L133_157 V133 V157 5.178338390971147e-13
C133_157 V133 V157 9.44434632382649e-19

R133_158 V133 V158 -261.2680582495368
L133_158 V133 V158 -4.0650601164486554e-12
C133_158 V133 V158 1.0703709660913403e-19

R133_159 V133 V159 -707.4949609118532
L133_159 V133 V159 -4.861842399254473e-12
C133_159 V133 V159 -6.690769724559754e-20

R133_160 V133 V160 -156.9624990389876
L133_160 V133 V160 -2.5884801895936054e-12
C133_160 V133 V160 -2.892411793207396e-20

R133_161 V133 V161 387.13242492299634
L133_161 V133 V161 1.0396471020507542e-11
C133_161 V133 V161 1.3998244133675856e-19

R133_162 V133 V162 220.97994330244111
L133_162 V133 V162 -4.421477343804638e-12
C133_162 V133 V162 -1.785263563632672e-19

R133_163 V133 V163 173.3066998443563
L133_163 V133 V163 1.764159827956922e-12
C133_163 V133 V163 2.2572942575724446e-19

R133_164 V133 V164 111.44941936427847
L133_164 V133 V164 2.013614271107894e-12
C133_164 V133 V164 -1.9456010010478057e-20

R133_165 V133 V165 1074.507865444276
L133_165 V133 V165 -1.975378171364141e-12
C133_165 V133 V165 -3.766807541633161e-19

R133_166 V133 V166 203.79798764962592
L133_166 V133 V166 4.868316766731887e-12
C133_166 V133 V166 1.1689485742952253e-19

R133_167 V133 V167 687.0313026630193
L133_167 V133 V167 4.125318176981727e-12
C133_167 V133 V167 9.759765199845792e-20

R133_168 V133 V168 -345.33219673578753
L133_168 V133 V168 3.85135556427939e-12
C133_168 V133 V168 2.977825607327448e-19

R133_169 V133 V169 -3334.016777922733
L133_169 V133 V169 6.031312396591462e-12
C133_169 V133 V169 1.8585353438693511e-19

R133_170 V133 V170 -101.54596626534477
L133_170 V133 V170 -4.133069284124684e-12
C133_170 V133 V170 -2.13116255313888e-19

R133_171 V133 V171 -174.35201517366667
L133_171 V133 V171 -1.0087055520808943e-12
C133_171 V133 V171 -4.2742915019104924e-19

R133_172 V133 V172 -186.43766472830433
L133_172 V133 V172 -1.82087868343914e-12
C133_172 V133 V172 -2.932308476709794e-19

R133_173 V133 V173 444.32553912808834
L133_173 V133 V173 -1.0950010154121375e-11
C133_173 V133 V173 -1.9224482111542175e-19

R133_174 V133 V174 -686.1877889713508
L133_174 V133 V174 -4.889061053098565e-12
C133_174 V133 V174 3.1606398719259143e-19

R133_175 V133 V175 554.6215162380684
L133_175 V133 V175 -4.176577520748039e-12
C133_175 V133 V175 -1.6914423180066848e-19

R133_176 V133 V176 278.9093865711667
L133_176 V133 V176 -2.450826673091206e-12
C133_176 V133 V176 -3.9411401824877872e-19

R133_177 V133 V177 -347.8931144116959
L133_177 V133 V177 1.2919032924136657e-11
C133_177 V133 V177 3.385175026513782e-20

R133_178 V133 V178 83.0425767318914
L133_178 V133 V178 1.789893396001981e-12
C133_178 V133 V178 8.701234127618992e-20

R133_179 V133 V179 7890.169682327164
L133_179 V133 V179 1.0014429012599918e-12
C133_179 V133 V179 5.046766757316385e-19

R133_180 V133 V180 669.9912698320636
L133_180 V133 V180 1.0004318224125637e-12
C133_180 V133 V180 5.331585574752035e-19

R133_181 V133 V181 1642.0749135139035
L133_181 V133 V181 7.265907982501415e-12
C133_181 V133 V181 3.247589111286094e-19

R133_182 V133 V182 -154.24291461772404
L133_182 V133 V182 -7.9212278911526e-13
C133_182 V133 V182 -3.3078345175728955e-19

R133_183 V133 V183 -742.083352332935
L133_183 V133 V183 2.320172199471661e-12
C133_183 V133 V183 2.130932453921174e-19

R133_184 V133 V184 -290.4536112878945
L133_184 V133 V184 2.6011523461465454e-12
C133_184 V133 V184 4.476836547409758e-20

R133_185 V133 V185 233.43590396445765
L133_185 V133 V185 1.1256343460064981e-11
C133_185 V133 V185 -2.116300616683224e-19

R133_186 V133 V186 -111.4126933805587
L133_186 V133 V186 3.8481788961808276e-12
C133_186 V133 V186 2.5934115637736716e-19

R133_187 V133 V187 18279.31681514441
L133_187 V133 V187 -1.8060573945815865e-12
C133_187 V133 V187 -4.1018563549961426e-19

R133_188 V133 V188 389.5981314261475
L133_188 V133 V188 -1.124440241291394e-12
C133_188 V133 V188 -3.457428017359975e-19

R133_189 V133 V189 -437.9111859093255
L133_189 V133 V189 -1.5650014220406159e-12
C133_189 V133 V189 -3.8970359443763813e-19

R133_190 V133 V190 105.30920011025572
L133_190 V133 V190 2.6043922553393443e-12
C133_190 V133 V190 2.7217671643172532e-19

R133_191 V133 V191 158.68109243833078
L133_191 V133 V191 -1.074994274238381e-12
C133_191 V133 V191 -4.877659026530241e-19

R133_192 V133 V192 272.3856256403018
L133_192 V133 V192 -2.0401773039975316e-12
C133_192 V133 V192 -3.1165600518297157e-19

R133_193 V133 V193 -711.560946837196
L133_193 V133 V193 6.634268483252417e-12
C133_193 V133 V193 1.2150092216395718e-19

R133_194 V133 V194 4022.832827408039
L133_194 V133 V194 -2.138568933083207e-12
C133_194 V133 V194 1.2685379448254716e-19

R133_195 V133 V195 -290.64805689062
L133_195 V133 V195 7.417229016489269e-13
C133_195 V133 V195 9.006337145364746e-19

R133_196 V133 V196 -1280.8447213420304
L133_196 V133 V196 9.356849508846494e-13
C133_196 V133 V196 4.660771591711594e-19

R133_197 V133 V197 -844.5632289885325
L133_197 V133 V197 1.4038148410556137e-12
C133_197 V133 V197 5.23276081259159e-19

R133_198 V133 V198 -172.19441735898667
L133_198 V133 V198 -7.877042107371316e-12
C133_198 V133 V198 -3.176357178817822e-20

R133_199 V133 V199 -211.03025509007213
L133_199 V133 V199 1.8784791568901562e-12
C133_199 V133 V199 2.634836736490748e-19

R133_200 V133 V200 -157.15647005104083
L133_200 V133 V200 2.4690821556571963e-12
C133_200 V133 V200 1.8285607948461183e-19

R134_134 V134 0 80.96130318620176
L134_134 V134 0 -1.0929022753068211e-11
C134_134 V134 0 1.1936397263461548e-18

R134_135 V134 V135 -165.3364964779304
L134_135 V134 V135 1.9435127578448275e-12
C134_135 V134 V135 3.215743820334654e-19

R134_136 V134 V136 -95.53144414935505
L134_136 V134 V136 1.730388208486415e-12
C134_136 V134 V136 6.706376290191688e-19

R134_137 V134 V137 -63.44947556883073
L134_137 V134 V137 1.9690004735744197e-12
C134_137 V134 V137 5.310444717019484e-19

R134_138 V134 V138 53.10832697262533
L134_138 V134 V138 1.0315562589762152e-12
C134_138 V134 V138 7.680358561871805e-19

R134_139 V134 V139 81.59327132928777
L134_139 V134 V139 -7.841000387510545e-12
C134_139 V134 V139 -1.4348714911864583e-19

R134_140 V134 V140 46.29139855385528
L134_140 V134 V140 -2.194415376953323e-12
C134_140 V134 V140 -7.116492736398161e-19

R134_141 V134 V141 -414.4693397806428
L134_141 V134 V141 -8.729234196329474e-13
C134_141 V134 V141 -8.773118477075554e-19

R134_142 V134 V142 37.6722160617051
L134_142 V134 V142 7.664831541668199e-13
C134_142 V134 V142 3.222074755291362e-19

R134_143 V134 V143 -432.2466935060159
L134_143 V134 V143 -2.609697670834769e-12
C134_143 V134 V143 -3.293020461190151e-19

R134_144 V134 V144 -719.1983174408991
L134_144 V134 V144 1.74293234952856e-11
C134_144 V134 V144 -6.216318422649753e-20

R134_145 V134 V145 39.18853166277636
L134_145 V134 V145 -8.155577499211831e-12
C134_145 V134 V145 -4.2336256152512192e-19

R134_146 V134 V146 -56.55880753091011
L134_146 V134 V146 -6.195787672381765e-13
C134_146 V134 V146 -3.1656273996410896e-19

R134_147 V134 V147 269.65795323375625
L134_147 V134 V147 3.754002135153725e-12
C134_147 V134 V147 3.484960292172541e-19

R134_148 V134 V148 -630.3516632523714
L134_148 V134 V148 4.329820415775876e-12
C134_148 V134 V148 4.85480050790081e-19

R134_149 V134 V149 -73.70499618359725
L134_149 V134 V149 5.328484380128952e-13
C134_149 V134 V149 1.4645970045397077e-18

R134_150 V134 V150 -18.303630483652565
L134_150 V134 V150 -1.8275613427801658e-11
C134_150 V134 V150 -8.040381116243909e-19

R134_151 V134 V151 197.5612849253115
L134_151 V134 V151 7.878476514710752e-12
C134_151 V134 V151 1.0286458999398499e-19

R134_152 V134 V152 80.54929544661269
L134_152 V134 V152 -2.7329184569587586e-12
C134_152 V134 V152 -2.1553147483966301e-19

R134_153 V134 V153 -57.80152097831002
L134_153 V134 V153 -5.576030406266993e-12
C134_153 V134 V153 1.6757900314986504e-19

R134_154 V134 V154 43.533343157303825
L134_154 V134 V154 3.0672467505824244e-12
C134_154 V134 V154 8.263790781751961e-19

R134_155 V134 V155 1003.7236370406446
L134_155 V134 V155 3.624510586270707e-11
C134_155 V134 V155 1.2605358420833564e-19

R134_156 V134 V156 -64.38418784644486
L134_156 V134 V156 7.99680299187434e-12
C134_156 V134 V156 -1.6685773323412234e-19

R134_157 V134 V157 156.4655694882666
L134_157 V134 V157 -6.472439022141969e-13
C134_157 V134 V157 -1.240973744272326e-18

R134_158 V134 V158 28.891257465745962
L134_158 V134 V158 2.498679677446855e-12
C134_158 V134 V158 -1.954159382701237e-19

R134_159 V134 V159 -59.88752886669652
L134_159 V134 V159 1.2806301104927784e-11
C134_159 V134 V159 1.643899486334969e-19

R134_160 V134 V160 -81.36449139254033
L134_160 V134 V160 2.1953125262772195e-12
C134_160 V134 V160 4.475052304471141e-19

R134_161 V134 V161 52.38498127882482
L134_161 V134 V161 -3.552781476620904e-12
C134_161 V134 V161 -3.3676747920040995e-19

R134_162 V134 V162 -177.55368517913962
L134_162 V134 V162 -6.977468885954474e-12
C134_162 V134 V162 4.2334842367860125e-20

R134_163 V134 V163 78.10479416244289
L134_163 V134 V163 -1.7155526650512114e-12
C134_163 V134 V163 -4.2217846198851696e-19

R134_164 V134 V164 52.183108122089926
L134_164 V134 V164 -3.043980964714897e-12
C134_164 V134 V164 -3.1274294187287114e-19

R134_165 V134 V165 -108.30274316520656
L134_165 V134 V165 6.588585125301264e-13
C134_165 V134 V165 1.0210438563574869e-18

R134_166 V134 V166 -18.48610283965906
L134_166 V134 V166 -4.945032252249862e-11
C134_166 V134 V166 5.2890544315993595e-20

R134_167 V134 V167 103.23964337356858
L134_167 V134 V167 -4.654821189132873e-12
C134_167 V134 V167 -1.645428580557553e-19

R134_168 V134 V168 87.49679938269921
L134_168 V134 V168 -1.6334328921673156e-12
C134_168 V134 V168 -3.343351311723405e-19

R134_169 V134 V169 -50.6301328427845
L134_169 V134 V169 6.18734693170563e-12
C134_169 V134 V169 1.9637211937054604e-19

R134_170 V134 V170 29.181352196998795
L134_170 V134 V170 2.2537465947089467e-12
C134_170 V134 V170 3.9995075884486217e-19

R134_171 V134 V171 -98.62872479218258
L134_171 V134 V171 7.87121322262359e-13
C134_171 V134 V171 8.190509991682185e-19

R134_172 V134 V172 -81.51072237766857
L134_172 V134 V172 8.376508102126041e-13
C134_172 V134 V172 6.042119577997686e-19

R134_173 V134 V173 40.647930421368656
L134_173 V134 V173 -9.691901492928172e-13
C134_173 V134 V173 -5.571590515472157e-19

R134_174 V134 V174 34.735214792829304
L134_174 V134 V174 -6.476016239200584e-11
C134_174 V134 V174 -3.901901570003648e-19

R134_175 V134 V175 -149.09753976766783
L134_175 V134 V175 -8.270349024899e-12
C134_175 V134 V175 -7.315318900080818e-20

R134_176 V134 V176 -170.75404491248878
L134_176 V134 V176 -2.4168356572382075e-12
C134_176 V134 V176 -2.93231285291922e-19

R134_177 V134 V177 379.35627837507667
L134_177 V134 V177 3.4592972723569116e-12
C134_177 V134 V177 2.9932082703286097e-19

R134_178 V134 V178 -35.466694529502945
L134_178 V134 V178 -2.041166711493762e-12
C134_178 V134 V178 -2.7361835075829617e-19

R134_179 V134 V179 116.36617682952168
L134_179 V134 V179 -1.0783895092779333e-12
C134_179 V134 V179 -5.506139690950962e-19

R134_180 V134 V180 124.51529454613295
L134_180 V134 V180 -1.0755583551086264e-12
C134_180 V134 V180 -2.083178869296413e-19

R134_181 V134 V181 -70.23697617657277
L134_181 V134 V181 1.2956736914190172e-11
C134_181 V134 V181 -2.141512998963133e-19

R134_182 V134 V182 -60.69387081071394
L134_182 V134 V182 8.851862988608613e-13
C134_182 V134 V182 4.672180111457621e-19

R134_183 V134 V183 7142.374004033114
L134_183 V134 V183 -1.2124555609653444e-11
C134_183 V134 V183 -3.5856019346483326e-20

R134_184 V134 V184 450.774504547531
L134_184 V134 V184 2.3142158772950016e-12
C134_184 V134 V184 3.342628394128312e-21

R134_185 V134 V185 148.26481608977588
L134_185 V134 V185 -5.65325951514625e-12
C134_185 V134 V185 -6.49623618328944e-20

R134_186 V134 V186 200.54654447395905
L134_186 V134 V186 2.2811448415404183e-12
C134_186 V134 V186 4.114600418200883e-21

R134_187 V134 V187 -537.5085135404431
L134_187 V134 V187 1.4511729079312299e-12
C134_187 V134 V187 2.75915664336815e-19

R134_188 V134 V188 587.9483928281988
L134_188 V134 V188 4.801185195500765e-12
C134_188 V134 V188 1.688382808169865e-19

R134_189 V134 V189 -2673.9682216478227
L134_189 V134 V189 2.0533616097327644e-12
C134_189 V134 V189 5.97551843728997e-19

R134_190 V134 V190 501.024099238178
L134_190 V134 V190 -2.0942487676373635e-12
C134_190 V134 V190 -4.5943100855027e-19

R134_191 V134 V191 -10139.993075310711
L134_191 V134 V191 1.9499241000803752e-12
C134_191 V134 V191 5.053393571403154e-19

R134_192 V134 V192 -497.55323436393724
L134_192 V134 V192 1.9362784932519363e-12
C134_192 V134 V192 6.644820359851354e-19

R134_193 V134 V193 -402.0561370497311
L134_193 V134 V193 -3.430829849538143e-12
C134_193 V134 V193 -2.391531505771861e-19

R134_194 V134 V194 387.73125721785993
L134_194 V134 V194 5.755490911917141e-12
C134_194 V134 V194 2.6097240790672624e-19

R134_195 V134 V195 -3322.888421037616
L134_195 V134 V195 -1.0067744835703461e-12
C134_195 V134 V195 -6.931600892582322e-19

R134_196 V134 V196 7142.1795135028815
L134_196 V134 V196 -6.468289928890204e-13
C134_196 V134 V196 -1.2933879075435339e-18

R134_197 V134 V197 170.03534180933542
L134_197 V134 V197 -1.6078996818226255e-12
C134_197 V134 V197 -4.668601932754835e-19

R134_198 V134 V198 -77.44502487142168
L134_198 V134 V198 3.240878538610063e-12
C134_198 V134 V198 2.1288303215469899e-19

R134_199 V134 V199 -293.41389592448706
L134_199 V134 V199 -1.6853762109448333e-12
C134_199 V134 V199 -4.042889932764309e-19

R134_200 V134 V200 135.04510752792174
L134_200 V134 V200 -1.099112471014683e-11
C134_200 V134 V200 -1.045130684838503e-19

R135_135 V135 0 70.1534454300592
L135_135 V135 0 -5.178279449503793e-13
C135_135 V135 0 -9.131450856413285e-19

R135_136 V135 V136 -160.24435644989407
L135_136 V135 V136 1.922895508714212e-12
C135_136 V135 V136 6.020930841874105e-19

R135_137 V135 V137 -67.31797291765926
L135_137 V135 V137 -2.4151343278161583e-12
C135_137 V135 V137 9.638841959259108e-21

R135_138 V135 V138 188.6578236361557
L135_138 V135 V138 -1.8110901107990194e-12
C135_138 V135 V138 -4.3147628138712395e-19

R135_139 V135 V139 42.3449579571041
L135_139 V135 V139 2.760055079060048e-13
C135_139 V135 V139 2.6020111874473704e-18

R135_140 V135 V140 69.90242744740168
L135_140 V135 V140 -1.5785258030486922e-12
C135_140 V135 V140 -8.529279414616092e-19

R135_141 V135 V141 -253.324648520719
L135_141 V135 V141 2.7157401739078736e-12
C135_141 V135 V141 1.6714945849864972e-19

R135_142 V135 V142 109.44741771611746
L135_142 V135 V142 -5.677301209241079e-12
C135_142 V135 V142 -3.1947243564723505e-20

R135_143 V135 V143 79.7963080296909
L135_143 V135 V143 -3.488420672312626e-12
C135_143 V135 V143 -2.713603203916082e-19

R135_144 V135 V144 -279.711518667318
L135_144 V135 V144 8.93492148466778e-12
C135_144 V135 V144 2.5782918303986257e-19

R135_145 V135 V145 49.511898390042774
L135_145 V135 V145 2.269751679735633e-12
C135_145 V135 V145 -6.753339457360822e-20

R135_146 V135 V146 -136.57795533220943
L135_146 V135 V146 1.7728776434957733e-12
C135_146 V135 V146 2.445055320403509e-19

R135_147 V135 V147 -44.50719131364823
L135_147 V135 V147 -5.624389518177487e-13
C135_147 V135 V147 -1.4660827982585002e-18

R135_148 V135 V148 163.3874500859931
L135_148 V135 V148 9.987470452568804e-13
C135_148 V135 V148 4.1138792424629444e-19

R135_149 V135 V149 -120.94092979135219
L135_149 V135 V149 -2.1989518304381684e-12
C135_149 V135 V149 7.740725667722068e-20

R135_150 V135 V150 -60.215515327789056
L135_150 V135 V150 -1.1985734681080796e-11
C135_150 V135 V150 3.1311691719161783e-19

R135_151 V135 V151 -38.14235476473911
L135_151 V135 V151 5.097334468782464e-12
C135_151 V135 V151 6.114967774983932e-19

R135_152 V135 V152 396.8569871685894
L135_152 V135 V152 -1.3182714749939178e-12
C135_152 V135 V152 -2.499842592851312e-19

R135_153 V135 V153 -100.57963837577685
L135_153 V135 V153 -1.7826075824296703e-12
C135_153 V135 V153 -3.056964634871786e-19

R135_154 V135 V154 155.78527076324886
L135_154 V135 V154 -2.738164453373983e-12
C135_154 V135 V154 -4.343425131672761e-19

R135_155 V135 V155 26.484733708012204
L135_155 V135 V155 5.237228488120805e-13
C135_155 V135 V155 8.570700788370138e-19

R135_156 V135 V156 -189.2768626608715
L135_156 V135 V156 -3.4993424661395206e-11
C135_156 V135 V156 -4.1517996154405903e-19

R135_157 V135 V157 474.155343253754
L135_157 V135 V157 1.3935373380768418e-12
C135_157 V135 V157 2.9318747766076046e-19

R135_158 V135 V158 328.03271710595396
L135_158 V135 V158 8.792666515859205e-12
C135_158 V135 V158 2.106663641656512e-19

R135_159 V135 V159 66.10856778582261
L135_159 V135 V159 -6.470609554083831e-13
C135_159 V135 V159 -1.1479419194621235e-18

R135_160 V135 V160 -93.52259782523979
L135_160 V135 V160 9.433033094160919e-12
C135_160 V135 V160 2.97389825256419e-19

R135_161 V135 V161 167.56242684421144
L135_161 V135 V161 2.002693169506191e-12
C135_161 V135 V161 3.213154776084752e-19

R135_162 V135 V162 -178.32712483310078
L135_162 V135 V162 3.726589313786783e-12
C135_162 V135 V162 1.9851453931080007e-19

R135_163 V135 V163 -69.3483978549927
L135_163 V135 V163 3.654396969698334e-12
C135_163 V135 V163 7.707041784737732e-19

R135_164 V135 V164 139.4611620777559
L135_164 V135 V164 6.4558597998486686e-12
C135_164 V135 V164 1.7504862066963105e-20

R135_165 V135 V165 -293.7680712535449
L135_165 V135 V165 -1.4434234514601528e-12
C135_165 V135 V165 -4.121147005485481e-19

R135_166 V135 V166 -262.2790168016956
L135_166 V135 V166 -4.573596714510956e-11
C135_166 V135 V166 -2.5694350191825228e-20

R135_167 V135 V167 -66.80361276344824
L135_167 V135 V167 1.8416773494577334e-12
C135_167 V135 V167 5.42597146439752e-20

R135_168 V135 V168 160.4047744212881
L135_168 V135 V168 6.161571111542482e-12
C135_168 V135 V168 2.1860907011666047e-19

R135_169 V135 V169 -178.3833061485173
L135_169 V135 V169 -1.7221146915586884e-12
C135_169 V135 V169 -3.1685827621491026e-19

R135_170 V135 V170 128.6659292858382
L135_170 V135 V170 -4.725106604027202e-12
C135_170 V135 V170 -9.718603400915566e-20

R135_171 V135 V171 62.296013998921424
L135_171 V135 V171 -9.08786903171861e-13
C135_171 V135 V171 -5.283499509962074e-19

R135_172 V135 V172 -1463.47565351557
L135_172 V135 V172 -1.1604432405157683e-11
C135_172 V135 V172 -2.7722762956014326e-19

R135_173 V135 V173 157.74059322981114
L135_173 V135 V173 1.2423917985531605e-12
C135_173 V135 V173 3.792909222385997e-19

R135_174 V135 V174 -237.60298167780502
L135_174 V135 V174 -1.322814331130322e-11
C135_174 V135 V174 -2.8839992413392654e-20

R135_175 V135 V175 1571.3310904290454
L135_175 V135 V175 8.036379891661034e-13
C135_175 V135 V175 8.356549218562348e-19

R135_176 V135 V176 -520.5900823788638
L135_176 V135 V176 -1.7057338691334399e-12
C135_176 V135 V176 -4.117446679471159e-19

R135_177 V135 V177 -1697.613187987167
L135_177 V135 V177 -1.106795265008099e-11
C135_177 V135 V177 -5.205147342669096e-20

R135_178 V135 V178 -306.46862772154356
L135_178 V135 V178 2.0691187691352566e-11
C135_178 V135 V178 1.0204979719947976e-19

R135_179 V135 V179 986.0740151329978
L135_179 V135 V179 4.130941089490758e-12
C135_179 V135 V179 -4.309217009416609e-19

R135_180 V135 V180 -262.0264058355004
L135_180 V135 V180 2.0780842048303147e-12
C135_180 V135 V180 4.010061053192413e-19

R135_181 V135 V181 -222.79702855376232
L135_181 V135 V181 7.918915932813337e-12
C135_181 V135 V181 4.21772878969175e-20

R135_182 V135 V182 585.2443657822738
L135_182 V135 V182 -1.8337655824157786e-11
C135_182 V135 V182 1.1172660544282516e-20

R135_183 V135 V183 -223.38815532272073
L135_183 V135 V183 -1.3762310476920204e-12
C135_183 V135 V183 1.3011411997521175e-19

R135_184 V135 V184 175.53129333049344
L135_184 V135 V184 1.2240768612680141e-11
C135_184 V135 V184 -1.9838592906855353e-19

R135_185 V135 V185 234.320745416433
L135_185 V135 V185 6.956754963849886e-12
C135_185 V135 V185 1.918082487551703e-20

R135_186 V135 V186 -3253.482486966195
L135_186 V135 V186 -7.473437753575535e-12
C135_186 V135 V186 -2.1601609899071698e-19

R135_187 V135 V187 -309.8700895250535
L135_187 V135 V187 8.049883379290813e-13
C135_187 V135 V187 5.5062245276589825e-19

R135_188 V135 V188 541.1295821377445
L135_188 V135 V188 -1.937159038291825e-12
C135_188 V135 V188 1.0968540511463045e-20

R135_189 V135 V189 -2718.046871965443
L135_189 V135 V189 -1.7101591188852547e-12
C135_189 V135 V189 -3.056236055368109e-19

R135_190 V135 V190 -206.65277717920796
L135_190 V135 V190 -1.4910983717933502e-09
C135_190 V135 V190 1.8705104176889383e-19

R135_191 V135 V191 484.90584088010513
L135_191 V135 V191 -1.6152378594607557e-12
C135_191 V135 V191 -9.438468254140499e-19

R135_192 V135 V192 -171.46719700277905
L135_192 V135 V192 2.2209832511817208e-12
C135_192 V135 V192 3.3232341806115764e-20

R135_193 V135 V193 -222.81905547823837
L135_193 V135 V193 4.249066426477023e-12
C135_193 V135 V193 1.173209585778547e-19

R135_194 V135 V194 442.9339666868319
L135_194 V135 V194 -7.260256916363274e-12
C135_194 V135 V194 -1.8539614664656933e-19

R135_195 V135 V195 233.48444643062194
L135_195 V135 V195 1.066019903386107e-12
C135_195 V135 V195 1.523134767589872e-18

R135_196 V135 V196 692.1579680810574
L135_196 V135 V196 -1.272350589279175e-12
C135_196 V135 V196 -6.811545444624872e-19

R135_197 V135 V197 413.5983896710894
L135_197 V135 V197 1.855243279348906e-12
C135_197 V135 V197 2.3086507614633173e-19

R135_198 V135 V198 -890.9558397235859
L135_198 V135 V198 9.11367278700721e-12
C135_198 V135 V198 7.864643691526532e-20

R135_199 V135 V199 -231.20142127494725
L135_199 V135 V199 3.740868445074772e-12
C135_199 V135 V199 2.092451201181681e-19

R135_200 V135 V200 360.0204035976871
L135_200 V135 V200 1.4275442770152903e-12
C135_200 V135 V200 5.067246917718255e-19

R136_136 V136 0 28.397609224046377
L136_136 V136 0 3.4562840698733393e-13
C136_136 V136 0 2.871889158876912e-18

R136_137 V136 V137 -56.20707318372565
L136_137 V136 V137 -1.4849828850689193e-12
C136_137 V136 V137 -1.961902737597911e-19

R136_138 V136 V138 78.6704766575883
L136_138 V136 V138 -1.419828277192524e-12
C136_138 V136 V138 -6.386650595734053e-19

R136_139 V136 V139 57.50015334520301
L136_139 V136 V139 -9.844897191128423e-13
C136_139 V136 V139 -9.007871558746575e-19

R136_140 V136 V140 24.92455019889659
L136_140 V136 V140 3.9676342526600766e-13
C136_140 V136 V140 1.990044789954788e-18

R136_141 V136 V141 -263.34387980891614
L136_141 V136 V141 -1.2573976224897162e-11
C136_141 V136 V141 -1.6625409559815368e-19

R136_142 V136 V142 56.38622106678791
L136_142 V136 V142 -6.6309226607803744e-12
C136_142 V136 V142 -1.0265816317357999e-19

R136_143 V136 V143 -252.05147942954486
L136_143 V136 V143 -1.280094540560635e-10
C136_143 V136 V143 1.0984441872490316e-19

R136_144 V136 V144 114.89050937111048
L136_144 V136 V144 -1.3271671118155041e-11
C136_144 V136 V144 -1.7944581151720516e-19

R136_145 V136 V145 41.478358145017104
L136_145 V136 V145 1.6215056844314788e-12
C136_145 V136 V145 1.0196488839889902e-19

R136_146 V136 V146 -48.36622641350057
L136_146 V136 V146 1.4355288259278052e-12
C136_146 V136 V146 3.3085110399694855e-19

R136_147 V136 V147 -858.3163620692579
L136_147 V136 V147 1.650250357709362e-11
C136_147 V136 V147 8.205876048787621e-20

R136_148 V136 V148 -34.05394430574891
L136_148 V136 V148 -3.9341652047763236e-13
C136_148 V136 V148 -1.316600099512668e-18

R136_149 V136 V149 -101.19433814901086
L136_149 V136 V149 -8.421309544332751e-12
C136_149 V136 V149 1.170558591232534e-19

R136_150 V136 V150 -37.41235606225797
L136_150 V136 V150 -2.17529012139889e-12
C136_150 V136 V150 -1.3560882028580687e-19

R136_151 V136 V151 -1099.158379570706
L136_151 V136 V151 3.245642169854881e-12
C136_151 V136 V151 -9.563563909968223e-20

R136_152 V136 V152 -132.54916246203464
L136_152 V136 V152 7.216819487002133e-13
C136_152 V136 V152 4.879297333235841e-19

R136_153 V136 V153 -69.53246728967777
L136_153 V136 V153 7.326612933830652e-12
C136_153 V136 V153 1.6030284399743278e-21

R136_154 V136 V154 58.42230002600309
L136_154 V136 V154 2.23701159361612e-12
C136_154 V136 V154 -1.9145426710336314e-19

R136_155 V136 V155 154.3222772251591
L136_155 V136 V155 -1.0109116516691914e-11
C136_155 V136 V155 -9.326562009437924e-20

R136_156 V136 V156 76.72090529764188
L136_156 V136 V156 2.0989581294202968e-12
C136_156 V136 V156 9.068506437634468e-19

R136_157 V136 V157 245.7597159875859
L136_157 V136 V157 -2.2127783836315575e-12
C136_157 V136 V157 -5.109390379215068e-19

R136_158 V136 V158 302.2772091195204
L136_158 V136 V158 -4.430199684423762e-12
C136_158 V136 V158 1.3396836347264474e-19

R136_159 V136 V159 -68.75951297421551
L136_159 V136 V159 4.5481479914523794e-12
C136_159 V136 V159 2.1621581825873753e-19

R136_160 V136 V160 53.814035640061064
L136_160 V136 V160 -1.4321690371269512e-12
C136_160 V136 V160 -7.9995398353905895e-19

R136_161 V136 V161 105.63409548303378
L136_161 V136 V161 1.0212156998067064e-12
C136_161 V136 V161 3.8284365904544034e-19

R136_162 V136 V162 -108.94906106128339
L136_162 V136 V162 2.6923305899863026e-12
C136_162 V136 V162 8.659491561002641e-20

R136_163 V136 V163 144.53249282000036
L136_163 V136 V163 1.8455161377278094e-11
C136_163 V136 V163 -1.5245744121276401e-19

R136_164 V136 V164 -87.66061265454381
L136_164 V136 V164 -7.587345524250384e-12
C136_164 V136 V164 5.446634817193672e-19

R136_165 V136 V165 -107.91890863704636
L136_165 V136 V165 -1.5615954266331531e-12
C136_165 V136 V165 -2.2289436172947075e-19

R136_166 V136 V166 -168.64215158828114
L136_166 V136 V166 -4.5753669391412014e-12
C136_166 V136 V166 -2.968141614988498e-19

R136_167 V136 V167 -607.328256290418
L136_167 V136 V167 6.3794786140944534e-12
C136_167 V136 V167 1.6791762437158972e-19

R136_168 V136 V168 -130.36568295683776
L136_168 V136 V168 8.926916533802797e-13
C136_168 V136 V168 8.530295911235245e-20

R136_169 V136 V169 -85.98036431322552
L136_169 V136 V169 -2.079528266657374e-12
C136_169 V136 V169 -4.94188152862934e-19

R136_170 V136 V170 194.8240795120937
L136_170 V136 V170 4.8556596568294044e-12
C136_170 V136 V170 7.587068067001135e-20

R136_171 V136 V171 -620.4156478660317
L136_171 V136 V171 2.7673828657599147e-12
C136_171 V136 V171 -2.6886687527765435e-20

R136_172 V136 V172 81.40838605116684
L136_172 V136 V172 -7.56924766395612e-13
C136_172 V136 V172 -2.758969457967964e-19

R136_173 V136 V173 72.96653209889458
L136_173 V136 V173 1.4689358007596551e-12
C136_173 V136 V173 3.310305981414886e-19

R136_174 V136 V174 -820.499965811322
L136_174 V136 V174 -3.857495804242037e-12
C136_174 V136 V174 -1.097619528111286e-19

R136_175 V136 V175 -5707.324601731803
L136_175 V136 V175 -1.3073161427945912e-12
C136_175 V136 V175 -2.403269107090403e-19

R136_176 V136 V176 610.3524028240888
L136_176 V136 V176 9.940504619893465e-13
C136_176 V136 V176 9.06212162954527e-19

R136_177 V136 V177 -1010.0149827667841
L136_177 V136 V177 -5.2235586193945946e-11
C136_177 V136 V177 -3.3800796661817676e-20

R136_178 V136 V178 1313.2711715444157
L136_178 V136 V178 -6.674843069035603e-12
C136_178 V136 V178 3.4374931966858975e-20

R136_179 V136 V179 424.9487044117827
L136_179 V136 V179 -1.2318377180814854e-11
C136_179 V136 V179 4.232044566273281e-20

R136_180 V136 V180 -191.7857119866851
L136_180 V136 V180 -5.817080760386977e-12
C136_180 V136 V180 -7.572160294073651e-19

R136_181 V136 V181 -130.9054698292812
L136_181 V136 V181 -1.3152957636665917e-11
C136_181 V136 V181 -1.688054281597549e-21

R136_182 V136 V182 -244.71243031859277
L136_182 V136 V182 -1.4677940594091664e-11
C136_182 V136 V182 -7.477618365408652e-20

R136_183 V136 V183 388.3967830991708
L136_183 V136 V183 -4.483561375162903e-10
C136_183 V136 V183 -1.9884525562561644e-19

R136_184 V136 V184 164.5836514249342
L136_184 V136 V184 -1.294617781566002e-12
C136_184 V136 V184 2.1679417491118528e-19

R136_185 V136 V185 169.2332474544387
L136_185 V136 V185 7.670605585272881e-12
C136_185 V136 V185 1.4853251418086053e-20

R136_186 V136 V186 -4393.955382934523
L136_186 V136 V186 -2.252226537506245e-12
C136_186 V136 V186 9.296494395538655e-20

R136_187 V136 V187 546.1219162545934
L136_187 V136 V187 -2.4881010952042747e-12
C136_187 V136 V187 1.246876879433362e-19

R136_188 V136 V188 -159.6332593858381
L136_188 V136 V188 4.57337313738317e-13
C136_188 V136 V188 4.476323746941681e-19

R136_189 V136 V189 1302.7199195752128
L136_189 V136 V189 -1.939692457140187e-12
C136_189 V136 V189 -1.8753124670470037e-19

R136_190 V136 V190 -268.02924213818716
L136_190 V136 V190 1.0375735813673432e-11
C136_190 V136 V190 -1.064582859351174e-20

R136_191 V136 V191 -124.62231847324445
L136_191 V136 V191 1.174106163213806e-12
C136_191 V136 V191 2.628078689539818e-19

R136_192 V136 V192 318.7090653145206
L136_192 V136 V192 -7.267931570465447e-13
C136_192 V136 V192 -8.632804192618266e-19

R136_193 V136 V193 -241.81427604293958
L136_193 V136 V193 5.1139431771181963e-11
C136_193 V136 V193 -1.0158291365706748e-19

R136_194 V136 V194 1153.5429296194295
L136_194 V136 V194 -1.4887064850991376e-12
C136_194 V136 V194 -6.187092080809078e-19

R136_195 V136 V195 193.62762096861908
L136_195 V136 V195 -9.362566677562023e-13
C136_195 V136 V195 -8.93044425309651e-19

R136_196 V136 V196 670.1318202593467
L136_196 V136 V196 6.400897342267152e-13
C136_196 V136 V196 1.5662727138865784e-18

R136_197 V136 V197 184.24272556851264
L136_197 V136 V197 1.963550381022109e-12
C136_197 V136 V197 3.4112651891649646e-19

R136_198 V136 V198 -163.28222952165694
L136_198 V136 V198 1.530142903243034e-11
C136_198 V136 V198 -1.6191700522494294e-19

R136_199 V136 V199 -199.85414770267394
L136_199 V136 V199 2.532508468746488e-12
C136_199 V136 V199 1.4206328574301214e-19

R136_200 V136 V200 297.0805654233002
L136_200 V136 V200 -6.566655797209372e-12
C136_200 V136 V200 -1.7006113680866398e-19

R137_137 V137 0 27.852229534173883
L137_137 V137 0 -3.639735931073345e-13
C137_137 V137 0 -1.1895368990365517e-18

R137_138 V137 V138 118.57488443875
L137_138 V137 V138 -4.126405828450086e-12
C137_138 V137 V138 -2.76057412245618e-19

R137_139 V137 V139 62.12192542828601
L137_139 V137 V139 9.215060198433635e-12
C137_139 V137 V139 -1.276128373688927e-19

R137_140 V137 V140 51.31887196770677
L137_140 V137 V140 1.5799659461151582e-12
C137_140 V137 V140 2.1539311710638556e-19

R137_141 V137 V141 -382.6241670409312
L137_141 V137 V141 7.713043711967682e-13
C137_141 V137 V141 6.4257786443696005e-19

R137_142 V137 V142 35.459129744162745
L137_142 V137 V142 -2.571593220577721e-11
C137_142 V137 V142 -1.4225632103018574e-19

R137_143 V137 V143 64.71928497643331
L137_143 V137 V143 1.58297778877955e-12
C137_143 V137 V143 1.9393158409802737e-19

R137_144 V137 V144 47.67649762290068
L137_144 V137 V144 2.38799277709129e-12
C137_144 V137 V144 1.0249083399657837e-19

R137_145 V137 V145 17.881256653744554
L137_145 V137 V145 6.230996950034506e-13
C137_145 V137 V145 4.003163165406592e-19

R137_146 V137 V146 228.45359708553383
L137_146 V137 V146 1.4911082268662888e-12
C137_146 V137 V146 9.231093315693573e-20

R137_147 V137 V147 -361.494213113346
L137_147 V137 V147 -4.537154504463697e-12
C137_147 V137 V147 6.674178439403561e-20

R137_148 V137 V148 -63.400667958476994
L137_148 V137 V148 -4.287810194169659e-12
C137_148 V137 V148 -1.0989957531886502e-19

R137_149 V137 V149 -88.4193426452001
L137_149 V137 V149 -4.955764646761812e-13
C137_149 V137 V149 -9.052458691622351e-19

R137_150 V137 V150 -16.218958646670764
L137_150 V137 V150 -1.9771420858912438e-12
C137_150 V137 V150 5.245408222702273e-19

R137_151 V137 V151 -32.8538098322684
L137_151 V137 V151 -3.9876273999217185e-12
C137_151 V137 V151 -1.3791602312779146e-19

R137_152 V137 V152 -105.536537589527
L137_152 V137 V152 -6.93148261364616e-12
C137_152 V137 V152 4.9778142401419e-20

R137_153 V137 V153 -21.569817857906664
L137_153 V137 V153 -1.2249882092502984e-12
C137_153 V137 V153 -1.9468842191974884e-19

R137_154 V137 V154 -190.29067187108376
L137_154 V137 V154 -2.7816109364500267e-12
C137_154 V137 V154 -4.622370901363121e-19

R137_155 V137 V155 40.02716097877918
L137_155 V137 V155 -3.1190536942974417e-12
C137_155 V137 V155 -1.2752342609990082e-19

R137_156 V137 V156 -88.37394348444133
L137_156 V137 V156 -5.273705458450158e-12
C137_156 V137 V156 -3.6144619151639215e-20

R137_157 V137 V157 -79.9790338515868
L137_157 V137 V157 8.909779068201377e-13
C137_157 V137 V157 7.42911299442839e-19

R137_158 V137 V158 27.164319600009026
L137_158 V137 V158 9.346826379924794e-12
C137_158 V137 V158 -1.554126739831079e-20

R137_159 V137 V159 275.8629969003835
L137_159 V137 V159 3.757939098639345e-12
C137_159 V137 V159 -1.0278154784237368e-19

R137_160 V137 V160 43.67064441528503
L137_160 V137 V160 1.339121535972978e-11
C137_160 V137 V160 -2.196759088893145e-19

R137_161 V137 V161 39.42319234307231
L137_161 V137 V161 1.7156629669989179e-12
C137_161 V137 V161 1.9610019075059033e-19

R137_162 V137 V162 89.82403001084609
L137_162 V137 V162 1.792633968645687e-11
C137_162 V137 V162 -4.1309713134790134e-20

R137_163 V137 V163 189.6332051137725
L137_163 V137 V163 3.6210613338345986e-12
C137_163 V137 V163 1.9001521742009868e-19

R137_164 V137 V164 275.0580142348538
L137_164 V137 V164 2.7021782544176117e-12
C137_164 V137 V164 1.6019794046753597e-19

R137_165 V137 V165 149.60327877161419
L137_165 V137 V165 -2.4103058279162237e-12
C137_165 V137 V165 -5.326458310109939e-19

R137_166 V137 V166 -19.361410841437362
L137_166 V137 V166 3.2472808433905395e-11
C137_166 V137 V166 1.2506084620188445e-19

R137_167 V137 V167 -79.14286057138744
L137_167 V137 V167 9.313585408085387e-12
C137_167 V137 V167 1.0699839727399657e-19

R137_168 V137 V168 482.9542412190964
L137_168 V137 V168 7.73868399123889e-12
C137_168 V137 V168 2.6406890600709937e-19

R137_169 V137 V169 -39.17997529944938
L137_169 V137 V169 -1.8073427457195132e-12
C137_169 V137 V169 -1.7112917082327514e-19

R137_170 V137 V170 47.86522650169508
L137_170 V137 V170 -5.684306539210013e-12
C137_170 V137 V170 -2.450687236856826e-19

R137_171 V137 V171 191.70703294110308
L137_171 V137 V171 -1.9233489818514398e-12
C137_171 V137 V171 -3.4605131702372153e-19

R137_172 V137 V172 1845.3027976459073
L137_172 V137 V172 -1.8274468113359606e-12
C137_172 V137 V172 -3.2821058236020703e-19

R137_173 V137 V173 147.72055925806458
L137_173 V137 V173 2.285291555623492e-12
C137_173 V137 V173 3.233029845664431e-19

R137_174 V137 V174 32.483555048283634
L137_174 V137 V174 -4.1363833494064875e-12
C137_174 V137 V174 6.23522507699179e-20

R137_175 V137 V175 2156.0042955041913
L137_175 V137 V175 -4.493736447903297e-12
C137_175 V137 V175 -1.5170860871758373e-19

R137_176 V137 V176 -630.6926748501088
L137_176 V137 V176 -9.069864238904359e-12
C137_176 V137 V176 -3.4214647917235944e-20

R137_177 V137 V177 101.66687655182174
L137_177 V137 V177 2.6905860679035132e-12
C137_177 V137 V177 -2.2581507170743927e-20

R137_178 V137 V178 -44.32578754949
L137_178 V137 V178 4.130304904371341e-12
C137_178 V137 V178 2.007528036950007e-19

R137_179 V137 V179 200.40686478256228
L137_179 V137 V179 1.9707499261623517e-12
C137_179 V137 V179 3.951859766982003e-19

R137_180 V137 V180 1287.8459763012113
L137_180 V137 V180 1.7381808419974493e-12
C137_180 V137 V180 2.2953122525522237e-19

R137_181 V137 V181 -106.6227777071816
L137_181 V137 V181 -4.2442502290873296e-12
C137_181 V137 V181 1.8113715134247494e-19

R137_182 V137 V182 -72.79272411543683
L137_182 V137 V182 -1.6361838259671504e-12
C137_182 V137 V182 -2.6240401566410363e-19

R137_183 V137 V183 -265.5190574464053
L137_183 V137 V183 7.039778569296513e-12
C137_183 V137 V183 7.257554784189286e-21

R137_184 V137 V184 283.37175136881854
L137_184 V137 V184 5.140250332253859e-11
C137_184 V137 V184 1.5968879306636918e-20

R137_185 V137 V185 -138.66295636124167
L137_185 V137 V185 1.1099063050690976e-11
C137_185 V137 V185 -1.6908052783923053e-19

R137_186 V137 V186 83.10484394384235
L137_186 V137 V186 4.099422764405541e-12
C137_186 V137 V186 6.326719119241749e-20

R137_187 V137 V187 333.844554540286
L137_187 V137 V187 -3.710749009141838e-12
C137_187 V137 V187 -2.3867289792842044e-19

R137_188 V137 V188 -2761.350950561324
L137_188 V137 V188 -5.318987880688947e-11
C137_188 V137 V188 -1.1445434401027604e-19

R137_189 V137 V189 135.06314860249793
L137_189 V137 V189 -2.755246932584361e-12
C137_189 V137 V189 -2.7745990380061794e-19

R137_190 V137 V190 -968.1524877080916
L137_190 V137 V190 -1.3125881859323204e-09
C137_190 V137 V190 2.6192769172358583e-19

R137_191 V137 V191 -182.37032584220117
L137_191 V137 V191 -3.082998413356315e-12
C137_191 V137 V191 -1.3386433882218015e-19

R137_192 V137 V192 -530.8293392252411
L137_192 V137 V192 -1.8090301022101166e-12
C137_192 V137 V192 -2.8084114963435665e-19

R137_193 V137 V193 234.89397225681256
L137_193 V137 V193 -2.9856918020274643e-12
C137_193 V137 V193 1.555654446782375e-19

R137_194 V137 V194 -155.73554864194594
L137_194 V137 V194 -2.238433859070663e-12
C137_194 V137 V194 -1.9603144617793268e-19

R137_195 V137 V195 812.493576571594
L137_195 V137 V195 1.84030333019616e-12
C137_195 V137 V195 2.6120553262996593e-19

R137_196 V137 V196 -282.5258572910465
L137_196 V137 V196 1.1293756952583791e-12
C137_196 V137 V196 5.252570063276665e-19

R137_197 V137 V197 -322.06678394835825
L137_197 V137 V197 1.1208979690790354e-12
C137_197 V137 V197 3.216408022711934e-19

R137_198 V137 V198 -101.94037827014179
L137_198 V137 V198 9.009123438490878e-12
C137_198 V137 V198 -6.178343152079324e-20

R137_199 V137 V199 -295.80143173451626
L137_199 V137 V199 2.833098484592587e-12
C137_199 V137 V199 1.3367488820825438e-19

R137_200 V137 V200 93.27848461394488
L137_200 V137 V200 3.3963276332032432e-12
C137_200 V137 V200 8.061257885719213e-20

R138_138 V138 0 -53.885029328745226
L138_138 V138 0 3.8260548050841424e-13
C138_138 V138 0 -1.3978272972257268e-19

R138_139 V138 V139 -54.11226767466952
L138_139 V138 V139 2.563708753235516e-12
C138_139 V138 V139 3.914056496367578e-19

R138_140 V138 V140 -29.946878397702935
L138_140 V138 V140 2.4963091871754663e-12
C138_140 V138 V140 6.747784034294849e-19

R138_141 V138 V141 189.82780595274554
L138_141 V138 V141 7.156453722466577e-12
C138_141 V138 V141 3.070272694670188e-19

R138_142 V138 V142 -56.58607538403886
L138_142 V138 V142 -1.7428732051057748e-12
C138_142 V138 V142 -6.975446568505353e-20

R138_143 V138 V143 120.04071862828629
L138_143 V138 V143 3.9109166404713344e-11
C138_143 V138 V143 1.304773158313715e-19

R138_144 V138 V144 127.20889313641798
L138_144 V138 V144 -3.7192146219091556e-11
C138_144 V138 V144 -2.051836833599004e-20

R138_145 V138 V145 -65.06753476962406
L138_145 V138 V145 -8.47996956539998e-12
C138_145 V138 V145 1.82591377073989e-19

R138_146 V138 V146 33.79268277481013
L138_146 V138 V146 6.485818581219326e-13
C138_146 V138 V146 3.4820098339421813e-19

R138_147 V138 V147 -2412.5260743178187
L138_147 V138 V147 -2.0141817562976665e-12
C138_147 V138 V147 -5.306911453622211e-19

R138_148 V138 V148 180.08777068798773
L138_148 V138 V148 -1.5104072542104455e-12
C138_148 V138 V148 -4.908282640552724e-19

R138_149 V138 V149 183.56204055287992
L138_149 V138 V149 -5.49714925522838e-12
C138_149 V138 V149 -5.823231955075735e-19

R138_150 V138 V150 28.532136854595894
L138_150 V138 V150 -2.069345356994101e-11
C138_150 V138 V150 4.108116998527407e-19

R138_151 V138 V151 -118.68394471108543
L138_151 V138 V151 4.044462911675816e-11
C138_151 V138 V151 9.147688353398606e-20

R138_152 V138 V152 -76.79703732956638
L138_152 V138 V152 2.932848161046748e-12
C138_152 V138 V152 1.823436293764265e-19

R138_153 V138 V153 124.56867490073334
L138_153 V138 V153 3.5325218727542437e-12
C138_153 V138 V153 -8.646653758116305e-20

R138_154 V138 V154 -31.460426133635153
L138_154 V138 V154 -2.2991958983960776e-12
C138_154 V138 V154 -5.664063718563183e-19

R138_155 V138 V155 1178.2165594941
L138_155 V138 V155 1.500465202710875e-12
C138_155 V138 V155 4.835481441401145e-20

R138_156 V138 V156 94.31274411260165
L138_156 V138 V156 7.339618514853763e-12
C138_156 V138 V156 2.7544782750674358e-19

R138_157 V138 V157 -375.68168836173726
L138_157 V138 V157 -1.472770075429234e-10
C138_157 V138 V157 5.696075343454454e-19

R138_158 V138 V158 -103.38805682069501
L138_158 V138 V158 -6.226816931308884e-12
C138_158 V138 V158 1.4691761237257227e-19

R138_159 V138 V159 62.13417711605569
L138_159 V138 V159 -4.617049621618539e-12
C138_159 V138 V159 -1.8407839149119766e-19

R138_160 V138 V160 82.82022007250592
L138_160 V138 V160 -1.2974930794936021e-11
C138_160 V138 V160 -3.5722489523859563e-19

R138_161 V138 V161 -58.61577193400131
L138_161 V138 V161 5.0077943921382466e-12
C138_161 V138 V161 2.4002576477731285e-19

R138_162 V138 V162 91.35957715880475
L138_162 V138 V162 2.1182068094758514e-12
C138_162 V138 V162 1.1376889956312473e-19

R138_163 V138 V163 -65.88358839414771
L138_163 V138 V163 1.357791827251359e-11
C138_163 V138 V163 3.258019235353302e-19

R138_164 V138 V164 -47.8124163180322
L138_164 V138 V164 -4.88061452943552e-12
C138_164 V138 V164 2.843468781171652e-19

R138_165 V138 V165 107.92587782632613
L138_165 V138 V165 -1.4129160384668485e-12
C138_165 V138 V165 -7.026810679332764e-19

R138_166 V138 V166 54.84833730169045
L138_166 V138 V166 -4.425251616414455e-12
C138_166 V138 V166 -8.174927790198465e-20

R138_167 V138 V167 -583.0112131352898
L138_167 V138 V167 4.860831009957974e-12
C138_167 V138 V167 1.2630918652166196e-19

R138_168 V138 V168 1259.8862611297375
L138_168 V138 V168 1.7703719650945301e-12
C138_168 V138 V168 1.7045830993477975e-19

R138_169 V138 V169 51.67667946634407
L138_169 V138 V169 -5.2097094992597785e-12
C138_169 V138 V169 -2.6987072808373863e-19

R138_170 V138 V170 -70.73966679245018
L138_170 V138 V170 -7.107802848073636e-12
C138_170 V138 V170 -2.290055278656554e-19

R138_171 V138 V171 101.2842439655542
L138_171 V138 V171 -2.374367573330924e-12
C138_171 V138 V171 -5.598357049986121e-19

R138_172 V138 V172 104.42814885855037
L138_172 V138 V172 -1.3057521943053175e-12
C138_172 V138 V172 -4.530928356377184e-19

R138_173 V138 V173 -42.64222154927076
L138_173 V138 V173 1.551827571469766e-12
C138_173 V138 V173 5.854100880177719e-19

R138_174 V138 V174 -234.17711489898232
L138_174 V138 V174 4.277247494834124e-12
C138_174 V138 V174 2.161927381400396e-19

R138_175 V138 V175 941.5617422009043
L138_175 V138 V175 4.9782556167560415e-12
C138_175 V138 V175 2.0345811077119042e-19

R138_176 V138 V176 -230.22438845562505
L138_176 V138 V176 3.226194594066174e-12
C138_176 V138 V176 3.5775750558857615e-19

R138_177 V138 V177 -258.82546209906593
L138_177 V138 V177 -7.889520217570945e-12
C138_177 V138 V177 -1.7843247485086284e-19

R138_178 V138 V178 193.2329650619569
L138_178 V138 V178 1.4855198428061852e-11
C138_178 V138 V178 1.3712409446145512e-19

R138_179 V138 V179 -182.1112353969015
L138_179 V138 V179 1.2005595866573841e-11
C138_179 V138 V179 1.847741705807347e-19

R138_180 V138 V180 -332.5729268890617
L138_180 V138 V180 4.744916977883021e-12
C138_180 V138 V180 1.1086910881838136e-20

R138_181 V138 V181 71.30056508098049
L138_181 V138 V181 -5.7387764276597135e-12
C138_181 V138 V181 -4.03128557532592e-20

R138_182 V138 V182 75.33108956650227
L138_182 V138 V182 -3.746967810146762e-12
C138_182 V138 V182 -2.4606164580743747e-19

R138_183 V138 V183 -2661.365759720047
L138_183 V138 V183 -3.931012406928189e-12
C138_183 V138 V183 -2.924264584553867e-20

R138_184 V138 V184 -5484.711648625292
L138_184 V138 V184 -2.127183181188756e-12
C138_184 V138 V184 -5.538198723331634e-20

R138_185 V138 V185 -196.94605670189853
L138_185 V138 V185 1.8908488852709744e-11
C138_185 V138 V185 1.1133415266994626e-19

R138_186 V138 V186 233.40227096818052
L138_186 V138 V186 -1.5026091370427938e-12
C138_186 V138 V186 -9.422375739191151e-20

R138_187 V138 V187 663.874690508548
L138_187 V138 V187 3.138217980126605e-11
C138_187 V138 V187 -2.523718629419993e-20

R138_188 V138 V188 -293.50465346358334
L138_188 V138 V188 1.6251237468429262e-12
C138_188 V138 V188 2.2186905176965318e-20

R138_189 V138 V189 -924.9072217512091
L138_189 V138 V189 -2.0223358127571425e-11
C138_189 V138 V189 -3.4150833288950115e-19

R138_190 V138 V190 -459.8487195766846
L138_190 V138 V190 2.186922397019116e-12
C138_190 V138 V190 2.96730064394231e-19

R138_191 V138 V191 3289.977257929564
L138_191 V138 V191 6.956505955299671e-12
C138_191 V138 V191 -2.968817319504082e-19

R138_192 V138 V192 -14124.955227532799
L138_192 V138 V192 -2.013372008647086e-12
C138_192 V138 V192 -4.502923959173211e-19

R138_193 V138 V193 1319.2130458469444
L138_193 V138 V193 5.641492083119966e-11
C138_193 V138 V193 1.3588981411519323e-19

R138_194 V138 V194 3190.5927906029715
L138_194 V138 V194 -2.162187525395785e-12
C138_194 V138 V194 -3.2335612362783996e-19

R138_195 V138 V195 -4233.287870478716
L138_195 V138 V195 -4.762577899246125e-11
C138_195 V138 V195 3.9687314041917464e-19

R138_196 V138 V196 1095.286508522456
L138_196 V138 V196 1.2031414654324874e-12
C138_196 V138 V196 8.889830292108247e-19

R138_197 V138 V197 -216.25869154823977
L138_197 V138 V197 4.149740147626819e-12
C138_197 V138 V197 2.8524101916159567e-19

R138_198 V138 V198 116.05057141902704
L138_198 V138 V198 -9.165425130523875e-12
C138_198 V138 V198 -4.3772479490130665e-20

R138_199 V138 V199 386.2461628250616
L138_199 V138 V199 3.7016310661630006e-12
C138_199 V138 V199 3.0488278115450126e-19

R138_200 V138 V200 -166.02047262448167
L138_200 V138 V200 2.6829476894970543e-11
C138_200 V138 V200 2.8304747610793535e-20

R139_139 V139 0 -25.776713676383455
L139_139 V139 0 4.579405468926503e-13
C139_139 V139 0 4.660635578260954e-19

R139_140 V139 V140 -22.209074587693163
L139_140 V139 V140 1.1068188563418662e-12
C139_140 V139 V140 1.2314183992988119e-18

R139_141 V139 V141 110.41416744579175
L139_141 V139 V141 1.626336927776478e-11
C139_141 V139 V141 1.787616487402088e-20

R139_142 V139 V142 -62.276352872486285
L139_142 V139 V142 -6.29908168774186e-12
C139_142 V139 V142 -2.2669745613596708e-21

R139_143 V139 V143 203.2373986657312
L139_143 V139 V143 8.107382249451879e-13
C139_143 V139 V143 6.345931042090903e-19

R139_144 V139 V144 108.68377226121872
L139_144 V139 V144 -4.450917510904489e-11
C139_144 V139 V144 -3.4272372509460482e-19

R139_145 V139 V145 -48.17008974428139
L139_145 V139 V145 -4.8579450023286954e-12
C139_145 V139 V145 1.40427574458214e-19

R139_146 V139 V146 30.99327935190922
L139_146 V139 V146 7.323741153533027e-12
C139_146 V139 V146 -2.5536914299681486e-19

R139_147 V139 V147 40.07914984548369
L139_147 V139 V147 3.9009731463261645e-13
C139_147 V139 V147 1.9084798705308467e-18

R139_148 V139 V148 103.54012940491297
L139_148 V139 V148 -6.955389538348843e-13
C139_148 V139 V148 -5.980497026132883e-19

R139_149 V139 V149 1047.8843099188248
L139_149 V139 V149 -1.7578681732599804e-12
C139_149 V139 V149 -4.513089333623713e-19

R139_150 V139 V150 42.583297066949086
L139_150 V139 V150 4.030710252519111e-11
C139_150 V139 V150 -1.4071228761259449e-19

R139_151 V139 V151 130.35984293665067
L139_151 V139 V151 -1.6622664165835923e-12
C139_151 V139 V151 -8.676744945876031e-19

R139_152 V139 V152 -91.15544374103655
L139_152 V139 V152 9.921479071249462e-13
C139_152 V139 V152 3.650747725087019e-19

R139_153 V139 V153 99.60780264986194
L139_153 V139 V153 1.396866130837744e-12
C139_153 V139 V153 4.0885409063660007e-19

R139_154 V139 V154 -36.65373785192841
L139_154 V139 V154 4.750889292080323e-12
C139_154 V139 V154 3.278864201818901e-19

R139_155 V139 V155 -29.600409437874475
L139_155 V139 V155 -3.6069461573067564e-13
C139_155 V139 V155 -1.1934750464307462e-18

R139_156 V139 V156 140.22906133886548
L139_156 V139 V156 6.6038428927367325e-12
C139_156 V139 V156 5.978676504835518e-19

R139_157 V139 V157 676.6394305767185
L139_157 V139 V157 -3.050592420047262e-11
C139_157 V139 V157 2.132278141959615e-20

R139_158 V139 V158 353.41397228229425
L139_158 V139 V158 -9.010265944947437e-12
C139_158 V139 V158 -2.135515198746819e-19

R139_159 V139 V159 96.84082580649395
L139_159 V139 V159 4.236886010568323e-13
C139_159 V139 V159 1.412626946216311e-18

R139_160 V139 V160 93.72488070416661
L139_160 V139 V160 -5.043854599106653e-12
C139_160 V139 V160 -5.342464183100539e-19

R139_161 V139 V161 -69.44058571028762
L139_161 V139 V161 -1.797030057620221e-12
C139_161 V139 V161 -3.9689001639643323e-19

R139_162 V139 V162 88.58928951983205
L139_162 V139 V162 -2.7781556832101645e-12
C139_162 V139 V162 -2.4904399868407045e-19

R139_163 V139 V163 -1267.7924847363106
L139_163 V139 V163 -7.083026681821523e-11
C139_163 V139 V163 -7.605876970843018e-19

R139_164 V139 V164 -67.12206046585587
L139_164 V139 V164 -4.113720156009098e-12
C139_164 V139 V164 8.00281690941962e-20

R139_165 V139 V165 115.94292921968103
L139_165 V139 V165 3.780464131105318e-12
C139_165 V139 V165 2.335274900690169e-19

R139_166 V139 V166 -649.2390214227187
L139_166 V139 V166 -6.769647845639199e-12
C139_166 V139 V166 5.141443954759872e-20

R139_167 V139 V167 161.7129488417364
L139_167 V139 V167 -1.019656946419778e-12
C139_167 V139 V167 -9.470884699771121e-20

R139_168 V139 V168 2589.219549439879
L139_168 V139 V168 6.026688544885857e-12
C139_168 V139 V168 -2.2725652965571825e-19

R139_169 V139 V169 53.107130150622275
L139_169 V139 V169 1.219804994790262e-12
C139_169 V139 V169 4.1448096080636875e-19

R139_170 V139 V170 989.1452331348643
L139_170 V139 V170 1.9301158687773657e-12
C139_170 V139 V170 4.555961825855304e-21

R139_171 V139 V171 -954.2872103883277
L139_171 V139 V171 8.521308988329478e-13
C139_171 V139 V171 5.53164066073504e-19

R139_172 V139 V172 257.1046542082997
L139_172 V139 V172 -6.427421380746407e-12
C139_172 V139 V172 1.7397615762179316e-19

R139_173 V139 V173 -57.36811301981732
L139_173 V139 V173 -1.2701590831376205e-12
C139_173 V139 V173 -3.016358297976832e-19

R139_174 V139 V174 186.4599470844122
L139_174 V139 V174 -2.356974075981082e-09
C139_174 V139 V174 1.5630119367723949e-19

R139_175 V139 V175 -13155.730866174315
L139_175 V139 V175 -7.497456308654541e-13
C139_175 V139 V175 -1.0714375695077112e-18

R139_176 V139 V176 -178.07169018404795
L139_176 V139 V176 1.4059420018726316e-12
C139_176 V139 V176 6.231631810565657e-19

R139_177 V139 V177 -239.8591604746998
L139_177 V139 V177 3.666182881597853e-12
C139_177 V139 V177 2.4329826658336046e-20

R139_178 V139 V178 -138.60134897368587
L139_178 V139 V178 -7.446473384380157e-12
C139_178 V139 V178 -3.9528023836869474e-20

R139_179 V139 V179 -137.36380728387854
L139_179 V139 V179 9.700206481562738e-12
C139_179 V139 V179 6.4364435970805335e-19

R139_180 V139 V180 204.63234412147972
L139_180 V139 V180 -3.433935515217718e-12
C139_180 V139 V180 -4.418017105422706e-19

R139_181 V139 V181 79.11516213293623
L139_181 V139 V181 -4.418116810440316e-12
C139_181 V139 V181 -1.086927152411375e-19

R139_182 V139 V182 131.29300543468773
L139_182 V139 V182 -4.188671281038425e-12
C139_182 V139 V182 -1.5985266961910838e-19

R139_183 V139 V183 226.64245194083813
L139_183 V139 V183 1.1979513880862099e-12
C139_183 V139 V183 -1.520243272907015e-19

R139_184 V139 V184 -222.052921972896
L139_184 V139 V184 3.4844859771000707e-10
C139_184 V139 V184 2.0237978898998754e-19

R139_185 V139 V185 -317.7153924611311
L139_185 V139 V185 -3.1224367210734386e-12
C139_185 V139 V185 6.647294548086385e-21

R139_186 V139 V186 158.37289554037395
L139_186 V139 V186 8.194786335787197e-12
C139_186 V139 V186 2.470583737620232e-19

R139_187 V139 V187 362.8763894139554
L139_187 V139 V187 -4.973331429569824e-13
C139_187 V139 V187 -7.967557343621458e-19

R139_188 V139 V188 -180.20413115017794
L139_188 V139 V188 2.19039528040106e-12
C139_188 V139 V188 -3.7647111648389284e-20

R139_189 V139 V189 -241.9998458506908
L139_189 V139 V189 1.842656433823875e-12
C139_189 V139 V189 2.739943276314597e-19

R139_190 V139 V190 -5188.8188366494205
L139_190 V139 V190 -5.387923408268619e-10
C139_190 V139 V190 -6.674490941974032e-20

R139_191 V139 V191 -5852.708890952645
L139_191 V139 V191 8.692014947368901e-13
C139_191 V139 V191 1.1589385234897004e-18

R139_192 V139 V192 217.32050067303257
L139_192 V139 V192 -1.045648536810195e-12
C139_192 V139 V192 -1.6794085285152033e-19

R139_193 V139 V193 483.67441414858297
L139_193 V139 V193 -1.9177632554949794e-11
C139_193 V139 V193 -7.853948732766896e-20

R139_194 V139 V194 445.59690084545196
L139_194 V139 V194 3.4701611541071356e-12
C139_194 V139 V194 2.365689245309764e-19

R139_195 V139 V195 -333.79607162741763
L139_195 V139 V195 -6.64257080097964e-13
C139_195 V139 V195 -1.8892136570971756e-18

R139_196 V139 V196 1287.2007373557785
L139_196 V139 V196 4.800418829294137e-13
C139_196 V139 V196 1.1871937369266667e-18

R139_197 V139 V197 -731.9828781491782
L139_197 V139 V197 -2.80950724709319e-12
C139_197 V139 V197 -1.8617512636033117e-19

R139_198 V139 V198 159.4362904515992
L139_198 V139 V198 -4.495974348106784e-12
C139_198 V139 V198 -1.5607020815880299e-19

R139_199 V139 V199 233.2040685722119
L139_199 V139 V199 -3.988449885480992e-12
C139_199 V139 V199 -2.830740243811809e-20

R139_200 V139 V200 -127.21961230603857
L139_200 V139 V200 -1.0974682210984735e-12
C139_200 V139 V200 -6.947860355697729e-19

R140_140 V140 0 -19.795791395016323
L140_140 V140 0 -4.037116536825477e-13
C140_140 V140 0 -2.953887538659882e-18

R140_141 V140 V141 101.33913070502686
L140_141 V140 V141 -1.0980937425078874e-11
C140_141 V140 V141 1.0271327118767943e-19

R140_142 V140 V142 -31.60883445016001
L140_142 V140 V142 3.229771805455747e-11
C140_142 V140 V142 1.8035588076364512e-19

R140_143 V140 V143 65.65811751371999
L140_143 V140 V143 3.6891154408596464e-11
C140_143 V140 V143 -1.6090925068751292e-19

R140_144 V140 V144 47.36203052432629
L140_144 V140 V144 1.146275016631256e-12
C140_144 V140 V144 4.461231613578376e-19

R140_145 V140 V145 -38.68043950309357
L140_145 V140 V145 -1.7136230956599813e-12
C140_145 V140 V145 -1.329159197050223e-19

R140_146 V140 V146 15.623042002113493
L140_146 V140 V146 2.4818342588080742e-11
C140_146 V140 V146 -3.742630419657193e-19

R140_147 V140 V147 83.37934138939384
L140_147 V140 V147 1.6013231608976654e-11
C140_147 V140 V147 -2.286943264176715e-19

R140_148 V140 V148 35.57401528162986
L140_148 V140 V148 3.9161936427854084e-13
C140_148 V140 V148 1.4396283281366348e-18

R140_149 V140 V149 241.78851664375674
L140_149 V140 V149 2.635617543724366e-12
C140_149 V140 V149 9.609364958386523e-20

R140_150 V140 V150 25.420943905601376
L140_150 V140 V150 2.4613444023104098e-12
C140_150 V140 V150 1.2775313078566902e-19

R140_151 V140 V151 -203.06014598691743
L140_151 V140 V151 -3.2954478324127132e-12
C140_151 V140 V151 2.1542623536338515e-19

R140_152 V140 V152 -59.40720235353734
L140_152 V140 V152 -6.225284089968428e-13
C140_152 V140 V152 -5.6355145740677865e-19

R140_153 V140 V153 69.57914209138846
L140_153 V140 V153 -5.2603221870746446e-12
C140_153 V140 V153 -1.010985167283325e-19

R140_154 V140 V154 -19.85742348828738
L140_154 V140 V154 -1.2058437515283361e-12
C140_154 V140 V154 2.1732475303564923e-19

R140_155 V140 V155 -67.6672597135354
L140_155 V140 V155 3.663754808644974e-12
C140_155 V140 V155 1.6579061373016143e-19

R140_156 V140 V156 -131.64545674958197
L140_156 V140 V156 -1.827414008348706e-12
C140_156 V140 V156 -1.0548589031114342e-18

R140_157 V140 V157 -185.46560919204416
L140_157 V140 V157 6.406904351679393e-12
C140_157 V140 V157 4.459346331655517e-19

R140_158 V140 V158 -4406.283299308453
L140_158 V140 V158 2.1819403438954944e-12
C140_158 V140 V158 -1.3103549195999722e-19

R140_159 V140 V159 42.578055079008244
L140_159 V140 V159 -2.5578876070072606e-12
C140_159 V140 V159 -3.7156169889556834e-19

R140_160 V140 V160 51.509124163423955
L140_160 V140 V160 9.182309251652584e-13
C140_160 V140 V160 8.007218059280418e-19

R140_161 V140 V161 -42.7773993859704
L140_161 V140 V161 -9.347935979927919e-13
C140_161 V140 V161 -3.526478763324734e-19

R140_162 V140 V162 49.37429913981529
L140_162 V140 V162 -7.876141305204013e-12
C140_162 V140 V162 -8.39950244973445e-20

R140_163 V140 V163 -50.433950647872315
L140_163 V140 V163 -3.65914484155517e-12
C140_163 V140 V163 2.0296202754562898e-19

R140_164 V140 V164 -44.36612842425002
L140_164 V140 V164 -9.586473878140325e-12
C140_164 V140 V164 -4.805070205714996e-19

R140_165 V140 V165 57.32712632664379
L140_165 V140 V165 1.0122152304643636e-12
C140_165 V140 V165 2.326557568783926e-19

R140_166 V140 V166 -1309.9360635940795
L140_166 V140 V166 -2.7773531646720442e-11
C140_166 V140 V166 3.734781692813548e-19

R140_167 V140 V167 123.4025383249619
L140_167 V140 V167 1.1107674499506759e-11
C140_167 V140 V167 -1.392490492149096e-19

R140_168 V140 V168 193.37887827999847
L140_168 V140 V168 -9.873490565798668e-13
C140_168 V140 V168 -5.2412288143205864e-20

R140_169 V140 V169 30.420054842599917
L140_169 V140 V169 2.301660816520531e-12
C140_169 V140 V169 3.6479339865114457e-19

R140_170 V140 V170 195.72773829055672
L140_170 V140 V170 8.374530863595362e-12
C140_170 V140 V170 -1.1234290636874889e-19

R140_171 V140 V171 110.14641815123412
L140_171 V140 V171 -9.991548371298114e-12
C140_171 V140 V171 3.1325841737968013e-20

R140_172 V140 V172 1018.2492290872652
L140_172 V140 V172 8.199031044140462e-13
C140_172 V140 V172 2.717678406446876e-19

R140_173 V140 V173 -28.200807748852636
L140_173 V140 V173 -9.737389038434445e-13
C140_173 V140 V173 -2.560441105295797e-19

R140_174 V140 V174 199.52658311847352
L140_174 V140 V174 3.98633134731249e-10
C140_174 V140 V174 4.91534681437073e-21

R140_175 V140 V175 -207.79081005397657
L140_175 V140 V175 1.596608894731104e-12
C140_175 V140 V175 3.241922004717871e-19

R140_176 V140 V176 -119.35478579902288
L140_176 V140 V176 -1.1583057460004209e-12
C140_176 V140 V176 -9.821748214525048e-19

R140_177 V140 V177 -146.41669795118364
L140_177 V140 V177 2.842615086286286e-12
C140_177 V140 V177 1.426164923813495e-19

R140_178 V140 V178 -55.05954238149907
L140_178 V140 V178 -4.052194567423461e-12
C140_178 V140 V178 1.633377370386607e-20

R140_179 V140 V179 -197.66706301678718
L140_179 V140 V179 -1.3345662491626542e-11
C140_179 V140 V179 -1.6338436781139966e-19

R140_180 V140 V180 97.79515730542366
L140_180 V140 V180 4.311292477405913e-12
C140_180 V140 V180 7.144226544608989e-19

R140_181 V140 V181 42.572783794505774
L140_181 V140 V181 6.6805003176265284e-12
C140_181 V140 V181 -8.015779881151301e-20

R140_182 V140 V182 47.33895026992435
L140_182 V140 V182 1.570000878246002e-12
C140_182 V140 V182 1.452873317237645e-19

R140_183 V140 V183 -2122.9611635942047
L140_183 V140 V183 -1.8366258405331065e-11
C140_183 V140 V183 1.7681792682955188e-19

R140_184 V140 V184 -85.70846494020938
L140_184 V140 V184 2.4218890333795655e-12
C140_184 V140 V184 -2.1223136757691218e-19

R140_185 V140 V185 -137.68652847920086
L140_185 V140 V185 -2.9329499853829067e-12
C140_185 V140 V185 -6.171558180879649e-20

R140_186 V140 V186 87.43957080056619
L140_186 V140 V186 1.8727807735090733e-12
C140_186 V140 V186 -1.3604451599392663e-19

R140_187 V140 V187 -569.9790105158581
L140_187 V140 V187 1.585351244057309e-12
C140_187 V140 V187 -8.740239354218392e-21

R140_188 V140 V188 -10919.903028781353
L140_188 V140 V188 -5.834350843494525e-13
C140_188 V140 V188 -3.7612905359717595e-19

R140_189 V140 V189 -133.10647015776195
L140_189 V140 V189 2.663481966134664e-12
C140_189 V140 V189 2.427182541136761e-19

R140_190 V140 V190 -133.45069760149468
L140_190 V140 V190 -1.9966295425096302e-12
C140_190 V140 V190 1.2620056481821213e-20

R140_191 V140 V191 147.72432776995763
L140_191 V140 V191 -1.2709904408789386e-12
C140_191 V140 V191 -2.71197879837719e-19

R140_192 V140 V192 338.45463174132925
L140_192 V140 V192 5.374413182055055e-13
C140_192 V140 V192 9.742332129911233e-19

R140_193 V140 V193 184.62570599864742
L140_193 V140 V193 1.0571158891847286e-11
C140_193 V140 V193 8.704877387562813e-20

R140_194 V140 V194 190.71408618182303
L140_194 V140 V194 1.4194427031874963e-12
C140_194 V140 V194 5.773535883433409e-19

R140_195 V140 V195 -173.6177386685796
L140_195 V140 V195 1.0320392497303426e-12
C140_195 V140 V195 9.694955897923706e-19

R140_196 V140 V196 -288.51312082595166
L140_196 V140 V196 -4.5367068892894347e-13
C140_196 V140 V196 -1.874855507402474e-18

R140_197 V140 V197 -224.108025097237
L140_197 V140 V197 -2.402469285363422e-12
C140_197 V140 V197 -3.1556993143558954e-19

R140_198 V140 V198 70.91159420752777
L140_198 V140 V198 4.3937780142234065e-12
C140_198 V140 V198 1.8271768097508894e-19

R140_199 V140 V199 267.6671950909767
L140_199 V140 V199 -3.1933085057977644e-12
C140_199 V140 V199 -1.801339939542612e-19

R140_200 V140 V200 -92.82799238042163
L140_200 V140 V200 -1.4348247773516998e-11
C140_200 V140 V200 2.1584436191510638e-19

R141_141 V141 0 654.0314409930634
L141_141 V141 0 1.2857496215484305e-13
C141_141 V141 0 4.518997879039322e-18

R141_142 V141 V142 3414.4107838662344
L141_142 V141 V142 1.08057069941741e-12
C141_142 V141 V142 2.4120455063294277e-19

R141_143 V141 V143 -331.9628093881958
L141_143 V141 V143 -1.4447698534036913e-12
C141_143 V141 V143 -3.9080331531878495e-19

R141_144 V141 V144 -354.5435510882885
L141_144 V141 V144 -7.2353526764148745e-12
C141_144 V141 V144 -2.747546539349134e-19

R141_145 V141 V145 171.5218018991375
L141_145 V141 V145 -9.74737377182023e-13
C141_145 V141 V145 -3.924693469614618e-19

R141_146 V141 V146 -233.11284982630153
L141_146 V141 V146 -8.560239797033026e-13
C141_146 V141 V146 -4.189774867160572e-20

R141_147 V141 V147 -331.54997689033087
L141_147 V141 V147 -3.0492617858363573e-12
C141_147 V141 V147 -1.469577031079015e-19

R141_148 V141 V148 -304.4768569059076
L141_148 V141 V148 -1.0343695701626216e-12
C141_148 V141 V148 -2.1683069699701954e-19

R141_149 V141 V149 296.53906468488503
L141_149 V141 V149 2.2550804952066678e-13
C141_149 V141 V149 2.2523389823851884e-18

R141_150 V141 V150 -149.5178653828865
L141_150 V141 V150 2.0957919117805538e-10
C141_150 V141 V150 -1.2412709836827954e-18

R141_151 V141 V151 -572.4590216221585
L141_151 V141 V151 1.9426220930719046e-11
C141_151 V141 V151 2.3053715482557534e-19

R141_152 V141 V152 447.95465035191546
L141_152 V141 V152 3.654308583820421e-12
C141_152 V141 V152 4.3229716035299535e-20

R141_153 V141 V153 -1068.8616446387712
L141_153 V141 V153 1.4685787966938434e-12
C141_153 V141 V153 4.332759252625453e-19

R141_154 V141 V154 154.9442372404814
L141_154 V141 V154 1.7463390844891564e-12
C141_154 V141 V154 1.0057259470207445e-18

R141_155 V141 V155 123.93424777030593
L141_155 V141 V155 8.645738345647895e-13
C141_155 V141 V155 4.220445193746162e-19

R141_156 V141 V156 7047.776340074476
L141_156 V141 V156 2.094278258343303e-12
C141_156 V141 V156 3.90438212677905e-19

R141_157 V141 V157 -172.87304035548243
L141_157 V141 V157 -3.002831833462768e-13
C141_157 V141 V157 -1.769733670275597e-18

R141_158 V141 V158 -892.5238897108235
L141_158 V141 V158 3.2043999814567525e-12
C141_158 V141 V158 -5.2928172326634127e-20

R141_159 V141 V159 -244.68911184885013
L141_159 V141 V159 2.8356304226369218e-11
C141_159 V141 V159 1.2876903068364663e-19

R141_160 V141 V160 -397.7074611046777
L141_160 V141 V160 2.1333191516285045e-12
C141_160 V141 V160 1.8494629878978377e-19

R141_161 V141 V161 180.1836047387117
L141_161 V141 V161 -3.369968627330277e-12
C141_161 V141 V161 -5.175538582795007e-19

R141_162 V141 V162 -3469.820380152341
L141_162 V141 V162 1.6963846370010889e-12
C141_162 V141 V162 2.572116049409197e-19

R141_163 V141 V163 367.63837031804184
L141_163 V141 V163 -1.7470329370172296e-12
C141_163 V141 V163 -3.005787421601492e-19

R141_164 V141 V164 348.5379591554364
L141_164 V141 V164 -1.5549914858267038e-12
C141_164 V141 V164 -7.181637863033788e-20

R141_165 V141 V165 663.140607282309
L141_165 V141 V165 1.6032856612232712e-12
C141_165 V141 V165 6.63765600255922e-19

R141_166 V141 V166 -433.56497480156185
L141_166 V141 V166 -1.6816023997841145e-12
C141_166 V141 V166 -3.4217852399816163e-19

R141_167 V141 V167 -636.2851106313536
L141_167 V141 V167 -2.044119348587432e-12
C141_167 V141 V167 -2.513523941161077e-19

R141_168 V141 V168 365.5696534483755
L141_168 V141 V168 -2.88068490626862e-12
C141_168 V141 V168 -5.862944172685584e-19

R141_169 V141 V169 -134.67694333663871
L141_169 V141 V169 3.849512051441989e-12
C141_169 V141 V169 2.812954121305802e-19

R141_170 V141 V170 1253.8996309647823
L141_170 V141 V170 2.2758816348767303e-12
C141_170 V141 V170 4.6488347590969335e-19

R141_171 V141 V171 -501.16494483599496
L141_171 V141 V171 7.200298690064649e-13
C141_171 V141 V171 7.140762603076623e-19

R141_172 V141 V172 -352.26184284230055
L141_172 V141 V172 1.3012662723821333e-12
C141_172 V141 V172 5.946887336692672e-19

R141_173 V141 V173 229.8377910182078
L141_173 V141 V173 4.798646957856563e-12
C141_173 V141 V173 -7.454543623242367e-20

R141_174 V141 V174 672.8006776376297
L141_174 V141 V174 1.749977462949068e-12
C141_174 V141 V174 -2.2639913149838735e-19

R141_175 V141 V175 -16821.139404261303
L141_175 V141 V175 1.5483643902430157e-12
C141_175 V141 V175 4.2193750633610193e-19

R141_176 V141 V176 -2409.2170906317797
L141_176 V141 V176 1.1226450200856526e-12
C141_176 V141 V176 5.443706709674417e-19

R141_177 V141 V177 285.49507665269454
L141_177 V141 V177 -1.9043155086265106e-12
C141_177 V141 V177 -2.2997701758766773e-20

R141_178 V141 V178 -598.476412929707
L141_178 V141 V178 -1.226065939945857e-12
C141_178 V141 V178 -3.169275680084806e-19

R141_179 V141 V179 224.6017372700052
L141_179 V141 V179 -7.172481813113284e-13
C141_179 V141 V179 -9.040056210754067e-19

R141_180 V141 V180 390.8400878557616
L141_180 V141 V180 -6.153376724557672e-13
C141_180 V141 V180 -8.4720970683260765e-19

R141_181 V141 V181 -295.76960512187225
L141_181 V141 V181 3.321459883402641e-12
C141_181 V141 V181 -6.679235029721094e-19

R141_182 V141 V182 -430.73797530800204
L141_182 V141 V182 6.67493075422181e-13
C141_182 V141 V182 5.257344925075552e-19

R141_183 V141 V183 -402.68655994123446
L141_183 V141 V183 -1.3003781272121214e-12
C141_183 V141 V183 -2.089311905223041e-19

R141_184 V141 V184 -3171.9068521668537
L141_184 V141 V184 -1.769682147672725e-12
C141_184 V141 V184 -5.568137181757587e-20

R141_185 V141 V185 -560.5760540534774
L141_185 V141 V185 -2.615179172896927e-12
C141_185 V141 V185 3.696553818374374e-19

R141_186 V141 V186 1549.0432348818665
L141_186 V141 V186 -1.6303236471570145e-12
C141_186 V141 V186 -3.6444981513202715e-19

R141_187 V141 V187 -1783.0248177470203
L141_187 V141 V187 1.2168703134247338e-12
C141_187 V141 V187 6.04495543689036e-19

R141_188 V141 V188 2908.7338547241193
L141_188 V141 V188 7.858636570666068e-13
C141_188 V141 V188 4.2072351216966646e-19

R141_189 V141 V189 -3465.9645818590857
L141_189 V141 V189 1.7504381064967647e-12
C141_189 V141 V189 6.436078301351959e-19

R141_190 V141 V190 -2404.7718415207323
L141_190 V141 V190 -4.736639682784073e-12
C141_190 V141 V190 -4.871787779665989e-19

R141_191 V141 V191 1502.7490973904667
L141_191 V141 V191 7.021008290031769e-13
C141_191 V141 V191 5.477024631664781e-19

R141_192 V141 V192 7372.525474306288
L141_192 V141 V192 1.2530532218452501e-12
C141_192 V141 V192 5.961116856314992e-19

R141_193 V141 V193 259.86552319982076
L141_193 V141 V193 3.3796392676979193e-12
C141_193 V141 V193 -1.7317467923425516e-19

R141_194 V141 V194 -445.12628156707837
L141_194 V141 V194 1.5279771008019836e-12
C141_194 V141 V194 1.8066621726445737e-19

R141_195 V141 V195 -594.8355096489809
L141_195 V141 V195 -5.119117759141302e-13
C141_195 V141 V195 -1.0238442718950937e-18

R141_196 V141 V196 -437.2533111998385
L141_196 V141 V196 -6.71489889619309e-13
C141_196 V141 V196 -8.275059457452305e-19

R141_197 V141 V197 1705.510697791164
L141_197 V141 V197 -9.474169430916818e-13
C141_197 V141 V197 -7.372284685143768e-19

R141_198 V141 V198 -885.8818654464122
L141_198 V141 V198 3.118943574509489e-11
C141_198 V141 V198 8.326863566794528e-20

R141_199 V141 V199 3655.8544420335675
L141_199 V141 V199 -1.522730692606006e-12
C141_199 V141 V199 -2.770355345682049e-19

R141_200 V141 V200 276.894766450029
L141_200 V141 V200 -1.5674021973500845e-12
C141_200 V141 V200 -3.103326387786734e-19

R142_142 V142 0 -38.705155088732134
L142_142 V142 0 -1.5984719514719861e-12
C142_142 V142 0 -3.3512773903983735e-19

R142_143 V142 V143 -425.70764459322186
L142_143 V142 V143 3.580836724526838e-12
C142_143 V142 V143 8.531947768181447e-20

R142_144 V142 V144 -228.40082764288496
L142_144 V142 V144 -8.898728226325707e-12
C142_144 V142 V144 -2.1385656399238876e-20

R142_145 V142 V145 -26.594002727848398
L142_145 V142 V145 -4.416840759127958e-12
C142_145 V142 V145 1.3190624374482568e-19

R142_146 V142 V146 35.62875632639872
L142_146 V142 V146 5.950063428748414e-13
C142_146 V142 V146 1.1440570836852108e-19

R142_147 V142 V147 -1149.3899713700837
L142_147 V142 V147 -1.793389482175932e-11
C142_147 V142 V147 -4.681843440700786e-21

R142_148 V142 V148 104.96123819672002
L142_148 V142 V148 -1.1068667632222952e-11
C142_148 V142 V148 -9.116110094350038e-20

R142_149 V142 V149 56.85627431557922
L142_149 V142 V149 -6.795098816677606e-13
C142_149 V142 V149 -5.092869391554061e-19

R142_150 V142 V150 15.740565350664289
L142_150 V142 V150 1.6871192259141454e-12
C142_150 V142 V150 2.3086990498557414e-19

R142_151 V142 V151 -98302.00528867802
L142_151 V142 V151 -6.67120836128788e-12
C142_151 V142 V151 -1.1521418210175215e-19

R142_152 V142 V152 -86.87189672888188
L142_152 V142 V152 4.371669429581458e-12
C142_152 V142 V152 6.51955144055214e-20

R142_153 V142 V153 32.51899699698688
L142_153 V142 V153 3.161174952160335e-12
C142_153 V142 V153 -5.933412870938488e-21

R142_154 V142 V154 -47.27706439243897
L142_154 V142 V154 -2.0025848567408173e-12
C142_154 V142 V154 -2.053839124649277e-19

R142_155 V142 V155 -278.1975880218026
L142_155 V142 V155 -6.5792637992185774e-12
C142_155 V142 V155 1.4326132566020143e-20

R142_156 V142 V156 59.233765184892114
L142_156 V142 V156 3.650141078109678e-11
C142_156 V142 V156 -1.1175666151095864e-20

R142_157 V142 V157 -109.48508318858973
L142_157 V142 V157 7.617148659226233e-13
C142_157 V142 V157 4.290097815817013e-19

R142_158 V142 V158 -21.776682168706667
L142_158 V142 V158 -1.065015869847672e-12
C142_158 V142 V158 2.2748761059512575e-20

R142_159 V142 V159 60.75360273554329
L142_159 V142 V159 2.834253803937583e-11
C142_159 V142 V159 -4.024061462859229e-20

R142_160 V142 V160 143.0304900873701
L142_160 V142 V160 -2.8718633961549085e-12
C142_160 V142 V160 -7.624942867639627e-20

R142_161 V142 V161 -45.71962700639966
L142_161 V142 V161 5.78830513378517e-12
C142_161 V142 V161 4.9758982203683443e-20

R142_162 V142 V162 112.21572004071119
L142_162 V142 V162 2.6655265526382246e-12
C142_162 V142 V162 -4.124689114236195e-21

R142_163 V142 V163 -73.47116908223752
L142_163 V142 V163 2.2321497455139473e-12
C142_163 V142 V163 1.3168313043427097e-19

R142_164 V142 V164 -54.02281379093928
L142_164 V142 V164 4.860242434457821e-12
C142_164 V142 V164 5.294666821239027e-20

R142_165 V142 V165 85.27424521082789
L142_165 V142 V165 -8.198568749140534e-13
C142_165 V142 V165 -3.0271095139655015e-19

R142_166 V142 V166 15.690045130970368
L142_166 V142 V166 3.1631216909472737e-12
C142_166 V142 V166 -5.687643672717519e-20

R142_167 V142 V167 -146.46069897496554
L142_167 V142 V167 7.690935637434797e-12
C142_167 V142 V167 -5.958856909465119e-21

R142_168 V142 V168 -108.956633773024
L142_168 V142 V168 2.1844340972791798e-12
C142_168 V142 V168 6.983357387781207e-20

R142_169 V142 V169 43.140477518535235
L142_169 V142 V169 1.0364843367905907e-11
C142_169 V142 V169 6.372189989668145e-20

R142_170 V142 V170 -24.101580735095443
L142_170 V142 V170 -1.34721068623281e-12
C142_170 V142 V170 -9.144191338290327e-20

R142_171 V142 V171 125.37390828378307
L142_171 V142 V171 -9.532915785232011e-13
C142_171 V142 V171 -2.013411132573257e-19

R142_172 V142 V172 128.92861546522604
L142_172 V142 V172 -1.0709046485052374e-12
C142_172 V142 V172 -1.300681081325844e-19

R142_173 V142 V173 -39.3444478931768
L142_173 V142 V173 1.964534999438459e-12
C142_173 V142 V173 7.546542286893568e-20

R142_174 V142 V174 -28.915511209528105
L142_174 V142 V174 6.217168935881821e-12
C142_174 V142 V174 1.4290329463913776e-19

R142_175 V142 V175 181.95062833382062
L142_175 V142 V175 -1.1222645622047785e-11
C142_175 V142 V175 -1.1833142511739535e-20

R142_176 V142 V176 170.39942004051642
L142_176 V142 V176 5.1481800354280915e-12
C142_176 V142 V176 5.630809414593356e-20

R142_177 V142 V177 -335.57971329711125
L142_177 V142 V177 -2.5644506464159795e-12
C142_177 V142 V177 -1.175841186945282e-19

R142_178 V142 V178 28.761944345676
L142_178 V142 V178 1.6328900689816941e-12
C142_178 V142 V178 6.43520992867132e-20

R142_179 V142 V179 -146.81366616525565
L142_179 V142 V179 1.1571223136028484e-12
C142_179 V142 V179 2.260373937781646e-19

R142_180 V142 V180 -460.0083292070078
L142_180 V142 V180 1.3038299366304707e-12
C142_180 V142 V180 9.809895845956803e-20

R142_181 V142 V181 63.29195782214504
L142_181 V142 V181 2.8725590182640844e-12
C142_181 V142 V181 8.046448467902678e-20

R142_182 V142 V182 67.28720958579625
L142_182 V142 V182 -8.474854307874149e-13
C142_182 V142 V182 -1.6856911859510464e-19

R142_183 V142 V183 -1938.8083906201894
L142_183 V142 V183 6.820000801989731e-12
C142_183 V142 V183 2.4008871699016477e-20

R142_184 V142 V184 -155.3029120314623
L142_184 V142 V184 -5.942199973736587e-12
C142_184 V142 V184 1.8012601134336355e-20

R142_185 V142 V185 -164.46496115958522
L142_185 V142 V185 2.7370624701391746e-10
C142_185 V142 V185 3.9241633777351145e-20

R142_186 V142 V186 -101.11230956877937
L142_186 V142 V186 -7.637894964377398e-12
C142_186 V142 V186 3.575207473555024e-20

R142_187 V142 V187 -123388.59815057197
L142_187 V142 V187 -1.4091355705344974e-12
C142_187 V142 V187 -1.3327054911739618e-19

R142_188 V142 V188 -890.0609685776591
L142_188 V142 V188 -2.0843182218441286e-12
C142_188 V142 V188 -1.1249489930131716e-19

R142_189 V142 V189 -484.96611861928363
L142_189 V142 V189 -1.4684323002382098e-12
C142_189 V142 V189 -1.7187824771064814e-19

R142_190 V142 V190 -14554.766647707473
L142_190 V142 V190 2.3085652294243562e-12
C142_190 V142 V190 1.1244287818592928e-19

R142_191 V142 V191 253.45686546568544
L142_191 V142 V191 -1.7937556030676131e-12
C142_191 V142 V191 -1.721814793237607e-19

R142_192 V142 V192 195.49075262905097
L142_192 V142 V192 -2.2210075738111446e-12
C142_192 V142 V192 -1.5717110324867972e-19

R142_193 V142 V193 233.18340560613044
L142_193 V142 V193 1.7446448425588548e-12
C142_193 V142 V193 8.278413759896773e-20

R142_194 V142 V194 -472.96458299749554
L142_194 V142 V194 -4.751927175793968e-12
C142_194 V142 V194 8.592548095153807e-21

R142_195 V142 V195 -555.5540050512744
L142_195 V142 V195 1.1628932941656241e-12
C142_195 V142 V195 2.282580035708908e-19

R142_196 V142 V196 -518.6987094237583
L142_196 V142 V196 7.613331640271154e-13
C142_196 V142 V196 3.254867015783465e-19

R142_197 V142 V197 -156.73054518346552
L142_197 V142 V197 2.435070463124932e-12
C142_197 V142 V197 9.274828829288142e-20

R142_198 V142 V198 78.67695921348043
L142_198 V142 V198 -6.2816024776799e-12
C142_198 V142 V198 -1.0042167842583683e-19

R142_199 V142 V199 408.44720758632883
L142_199 V142 V199 1.9829433991821154e-12
C142_199 V142 V199 1.2157679318841112e-19

R142_200 V142 V200 -96.98317761383196
L142_200 V142 V200 3.447391612664224e-09
C142_200 V142 V200 3.2542042134947543e-20

R143_143 V143 0 156.6754747252363
L143_143 V143 0 2.2554153960572625e-12
C143_143 V143 0 9.728187283463552e-19

R143_144 V143 V144 -149.56569885957478
L143_144 V143 V144 -4.912469598896656e-12
C143_144 V143 V144 -1.3499536020376604e-20

R143_145 V143 V145 -50.8845144731864
L143_145 V143 V145 -1.7492130121151828e-12
C143_145 V143 V145 -1.3562711915188127e-19

R143_146 V143 V146 -59.94245958441021
L143_146 V143 V146 -1.811326625271354e-12
C143_146 V143 V146 -3.4670240289170156e-20

R143_147 V143 V147 66.33666302933685
L143_147 V143 V147 4.487139420489451e-12
C143_147 V143 V147 -1.9231991628346575e-19

R143_148 V143 V148 -70.40484920528058
L143_148 V143 V148 -3.6126704983583753e-12
C143_148 V143 V148 1.0166620089404603e-19

R143_149 V143 V149 89.35411903780248
L143_149 V143 V149 5.559362753773283e-13
C143_149 V143 V149 7.290528589269441e-19

R143_150 V143 V150 294.08525595042045
L143_150 V143 V150 5.0078880784261745e-12
C143_150 V143 V150 -3.695479862006251e-19

R143_151 V143 V151 23.34291780410628
L143_151 V143 V151 9.297819809589005e-13
C143_151 V143 V151 1.7906438337812532e-19

R143_152 V143 V152 136.1286768059586
L143_152 V143 V152 1.7849621900388875e-11
C143_152 V143 V152 -8.826370792688847e-20

R143_153 V143 V153 67.79558096812755
L143_153 V143 V153 1.1351569403264954e-11
C143_153 V143 V153 -8.047900137075329e-20

R143_154 V143 V154 50.924872486271475
L143_154 V143 V154 3.6347410514903057e-12
C143_154 V143 V154 2.7348743785992717e-19

R143_155 V143 V155 -42.05864985633799
L143_155 V143 V155 2.1080709410696786e-12
C143_155 V143 V155 4.1674898116539514e-19

R143_156 V143 V156 307.8384443373959
L143_156 V143 V156 4.159971685462895e-12
C143_156 V143 V156 -2.69685179004033e-20

R143_157 V143 V157 8109.183693967708
L143_157 V143 V157 -7.258331944033717e-13
C143_157 V143 V157 -6.943356651174203e-19

R143_158 V143 V158 -198.19056250388627
L143_158 V143 V158 1.2153581651960408e-11
C143_158 V143 V158 9.490939311165184e-21

R143_159 V143 V159 -20.590430050387596
L143_159 V143 V159 -6.396491328230548e-13
C143_159 V143 V159 -2.3280456257530556e-19

R143_160 V143 V160 391.50716194632906
L143_160 V143 V160 1.0646015899835891e-11
C143_160 V143 V160 1.6154431486150354e-19

R143_161 V143 V161 3880.0241594869703
L143_161 V143 V161 4.759278993262066e-12
C143_161 V143 V161 9.723848803735409e-20

R143_162 V143 V162 -259.40390013139154
L143_162 V143 V162 3.4156055145053133e-12
C143_162 V143 V162 3.6891600837555707e-20

R143_163 V143 V163 42.39266016277532
L143_163 V143 V163 7.657742250819902e-12
C143_163 V143 V163 -8.954916491511222e-20

R143_164 V143 V164 1151.8742984970354
L143_164 V143 V164 -4.0531865046955546e-12
C143_164 V143 V164 -7.494666394227414e-20

R143_165 V143 V165 -160.73592206476576
L143_165 V143 V165 1.088378096966913e-12
C143_165 V143 V165 4.109214718173245e-19

R143_166 V143 V166 3183.6842948792555
L143_166 V143 V166 9.603658640094136e-12
C143_166 V143 V166 -3.4359178352067344e-20

R143_167 V143 V167 29.9081962785049
L143_167 V143 V167 1.2868312766756381e-12
C143_167 V143 V167 7.127019254031656e-21

R143_168 V143 V168 -155.17098273263701
L143_168 V143 V168 8.352602652988182e-12
C143_168 V143 V168 -1.967699799876865e-20

R143_169 V143 V169 -171.0203914269586
L143_169 V143 V169 -3.017843107366387e-12
C143_169 V143 V169 -1.531079962905742e-19

R143_170 V143 V170 -142.9983224324076
L143_170 V143 V170 -8.757519679660232e-12
C143_170 V143 V170 2.0999955881017224e-19

R143_171 V143 V171 -30.385843002396083
L143_171 V143 V171 1.8619440840626827e-11
C143_171 V143 V171 2.4280313157174303e-19

R143_172 V143 V172 -329.57081432429356
L143_172 V143 V172 5.01000215873121e-12
C143_172 V143 V172 1.6100254060853509e-19

R143_173 V143 V173 109.52872486397877
L143_173 V143 V173 -3.7444074326604756e-12
C143_173 V143 V173 -1.7751392131860143e-19

R143_174 V143 V174 135.35958188824324
L143_174 V143 V174 -1.2340844342583299e-11
C143_174 V143 V174 -2.662065153783577e-19

R143_175 V143 V175 -145.3192649997645
L143_175 V143 V175 2.1295665681429836e-11
C143_175 V143 V175 1.2969751955345295e-19

R143_176 V143 V176 228.96386083713233
L143_176 V143 V176 -8.242982131343282e-12
C143_176 V143 V176 -1.2474369546842363e-19

R143_177 V143 V177 375.91397310184175
L143_177 V143 V177 -5.715243675368418e-11
C143_177 V143 V177 1.1420088574522701e-19

R143_178 V143 V178 234.19923209785043
L143_178 V143 V178 -4.577348838104107e-12
C143_178 V143 V178 -1.1682759480252285e-19

R143_179 V143 V179 60.95695371712392
L143_179 V143 V179 -2.9635285349419023e-12
C143_179 V143 V179 -3.497656221646655e-19

R143_180 V143 V180 409.61619347434754
L143_180 V143 V180 -2.2625707313676963e-12
C143_180 V143 V180 -1.4165865192326467e-19

R143_181 V143 V181 -197.10165085029945
L143_181 V143 V181 4.682410780156567e-12
C143_181 V143 V181 3.569074327168421e-20

R143_182 V143 V182 -101.50999351699002
L143_182 V143 V182 1.428169402682978e-12
C143_182 V143 V182 2.5196182671415344e-19

R143_183 V143 V183 -477.1799652430226
L143_183 V143 V183 -1.9679568019729782e-12
C143_183 V143 V183 -2.2201956234656996e-20

R143_184 V143 V184 -363.95298106599876
L143_184 V143 V184 -8.714426669511158e-12
C143_184 V143 V184 1.552637138308876e-20

R143_185 V143 V185 11240.697429021642
L143_185 V143 V185 5.9503232287601065e-12
C143_185 V143 V185 -6.248817204077489e-20

R143_186 V143 V186 -280.8547247889853
L143_186 V143 V186 1.3566116372246354e-11
C143_186 V143 V186 -1.038481397189857e-20

R143_187 V143 V187 9726.364569627456
L143_187 V143 V187 8.506623254229907e-13
C143_187 V143 V187 3.3695270415522506e-19

R143_188 V143 V188 612.1433231378409
L143_188 V143 V188 1.0992398969667933e-12
C143_188 V143 V188 1.9977189117334508e-19

R143_189 V143 V189 446.47931092522305
L143_189 V143 V189 -5.147764545877229e-12
C143_189 V143 V189 1.2410768554906913e-19

R143_190 V143 V190 144.7312718279426
L143_190 V143 V190 -4.373806252996429e-12
C143_190 V143 V190 -2.144628474606608e-19

R143_191 V143 V191 603.676506800277
L143_191 V143 V191 4.027819366888386e-12
C143_191 V143 V191 -3.0304349731558414e-20

R143_192 V143 V192 223.3823325716117
L143_192 V143 V192 9.371488735467053e-12
C143_192 V143 V192 9.063411864714592e-20

R143_193 V143 V193 342.50547661504106
L143_193 V143 V193 -7.56324285042936e-12
C143_193 V143 V193 -1.3141887902371162e-19

R143_194 V143 V194 -537.8581139485622
L143_194 V143 V194 -2.4368920545978932e-12
C143_194 V143 V194 -9.518823146418419e-20

R143_195 V143 V195 -128.0054875961557
L143_195 V143 V195 -1.819185321635668e-12
C143_195 V143 V195 7.006659366135407e-21

R143_196 V143 V196 -618.8373984301963
L143_196 V143 V196 -8.950503773304256e-13
C143_196 V143 V196 -5.095269151363993e-19

R143_197 V143 V197 -1159.55997726049
L143_197 V143 V197 -5.3834487752345e-12
C143_197 V143 V197 -8.235601125667733e-20

R143_198 V143 V198 -182.55576991017128
L143_198 V143 V198 4.463616461395471e-12
C143_198 V143 V198 9.053513261081223e-20

R143_199 V143 V199 346.3409862416207
L143_199 V143 V199 -4.729100795423436e-11
C143_199 V143 V199 -1.898732301854992e-19

R143_200 V143 V200 602.205288038843
L143_200 V143 V200 4.767710948770334e-12
C143_200 V143 V200 9.858224021387317e-20

R144_144 V144 0 -30.519896770007932
L144_144 V144 0 9.4345627502675e-13
C144_144 V144 0 8.225733383597845e-19

R144_145 V144 V145 -37.40066550730252
L144_145 V144 V145 -1.92230509930238e-12
C144_145 V144 V145 -7.301511663997046e-20

R144_146 V144 V146 -44.8242443396911
L144_146 V144 V146 -2.966763540801473e-12
C144_146 V144 V146 4.146326175025779e-20

R144_147 V144 V147 -105.41475174992841
L144_147 V144 V147 -6.679227578021268e-12
C144_147 V144 V147 1.119521900871185e-19

R144_148 V144 V148 26.162924957524318
L144_148 V144 V148 5.066757431838458e-12
C144_148 V144 V148 -1.7119931379636564e-19

R144_149 V144 V149 89.31464154015164
L144_149 V144 V149 2.5174248670104006e-12
C144_149 V144 V149 2.210801446010474e-19

R144_150 V144 V150 117.59441191732974
L144_150 V144 V150 4.7207490129924785e-12
C144_150 V144 V150 -1.842087006354977e-19

R144_151 V144 V151 292.94481971232204
L144_151 V144 V151 8.945817407581335e-12
C144_151 V144 V151 -6.887364993931766e-20

R144_152 V144 V152 26.307392324781503
L144_152 V144 V152 1.2466469035008242e-12
C144_152 V144 V152 9.547279846277941e-20

R144_153 V144 V153 48.283158141835486
L144_153 V144 V153 2.6357917821049494e-12
C144_153 V144 V153 1.4946586694368584e-19

R144_154 V144 V154 45.65636610732239
L144_154 V144 V154 2.459960196508634e-12
C144_154 V144 V154 1.3134915907737603e-19

R144_155 V144 V155 91.85297235090194
L144_155 V144 V155 6.142810766486797e-12
C144_155 V144 V155 2.1818260428748533e-20

R144_156 V144 V156 -90.49414907413467
L144_156 V144 V156 -8.971485119024527e-12
C144_156 V144 V156 2.5082046856404575e-19

R144_157 V144 V157 178.15167925058913
L144_157 V144 V157 -5.207835072138593e-12
C144_157 V144 V157 -2.5796004999220787e-19

R144_158 V144 V158 -1034.6307273160935
L144_158 V144 V158 -5.654051034554348e-12
C144_158 V144 V158 1.8187830407454522e-20

R144_159 V144 V159 135.4893959638526
L144_159 V144 V159 9.760702787909901e-12
C144_159 V144 V159 1.8454298279605832e-19

R144_160 V144 V160 -12.680817536305609
L144_160 V144 V160 -1.0590296259302334e-12
C144_160 V144 V160 -6.44175512568799e-20

R144_161 V144 V161 4735.2738044204725
L144_161 V144 V161 1.0628761966339498e-11
C144_161 V144 V161 -6.077533461255081e-20

R144_162 V144 V162 -167.78746053706027
L144_162 V144 V162 -5.100131722299721e-11
C144_162 V144 V162 5.338627264488612e-20

R144_163 V144 V163 463.40839421347175
L144_163 V144 V163 5.272487914016728e-11
C144_163 V144 V163 -8.327997500821363e-20

R144_164 V144 V164 19.761136542032286
L144_164 V144 V164 2.7811901995647777e-12
C144_164 V144 V164 4.4947853880826544e-21

R144_165 V144 V165 -336.17494945518007
L144_165 V144 V165 -7.24639115349306e-12
C144_165 V144 V165 9.652211720228057e-20

R144_166 V144 V166 306.8020831045607
L144_166 V144 V166 1.1216219689733627e-11
C144_166 V144 V166 -1.2395255126304012e-19

R144_167 V144 V167 -248.3318716776941
L144_167 V144 V167 -7.0059654239745e-12
C144_167 V144 V167 -5.277205996845624e-20

R144_168 V144 V168 37.952661581603834
L144_168 V144 V168 1.940943617297779e-12
C144_168 V144 V168 -1.3758347250587823e-19

R144_169 V144 V169 -132.9868467654237
L144_169 V144 V169 2.0200949700283236e-11
C144_169 V144 V169 1.2491083090446237e-19

R144_170 V144 V170 -167.52575543668326
L144_170 V144 V170 -5.111527071260285e-12
C144_170 V144 V170 1.0235630655194884e-19

R144_171 V144 V171 -342.52040443895066
L144_171 V144 V171 3.8867389203341935e-11
C144_171 V144 V171 1.1954523525023965e-19

R144_172 V144 V172 -28.074326826528498
L144_172 V144 V172 -3.202903885579973e-12
C144_172 V144 V172 4.388910417048909e-20

R144_173 V144 V173 84.39010882750449
L144_173 V144 V173 4.8968443168823795e-12
C144_173 V144 V173 -5.222982303712165e-20

R144_174 V144 V174 288.09373091163735
L144_174 V144 V174 4.579610148504106e-12
C144_174 V144 V174 4.7860142998202536e-20

R144_175 V144 V175 374.24805173096763
L144_175 V144 V175 6.6174669665023755e-12
C144_175 V144 V175 -3.056359477021601e-20

R144_176 V144 V176 -429.73828438912324
L144_176 V144 V176 -3.721515079087304e-12
C144_176 V144 V176 2.3440667535665453e-19

R144_177 V144 V177 140.11262714571046
L144_177 V144 V177 -4.595688426804123e-12
C144_177 V144 V177 -7.856469053378551e-20

R144_178 V144 V178 158.76880558039866
L144_178 V144 V178 4.13483523891925e-11
C144_178 V144 V178 -9.432515907726829e-20

R144_179 V144 V179 1298.350137646905
L144_179 V144 V179 -9.891087457052332e-12
C144_179 V144 V179 -3.6757085684497263e-20

R144_180 V144 V180 83.48436786274922
L144_180 V144 V180 1.228994473220909e-11
C144_180 V144 V180 -1.7207332634063889e-19

R144_181 V144 V181 -94.87935678776746
L144_181 V144 V181 -1.9914916588689083e-10
C144_181 V144 V181 -7.598279424193776e-20

R144_182 V144 V182 -67.72509801278981
L144_182 V144 V182 -5.708763064751532e-12
C144_182 V144 V182 2.5751227153076138e-20

R144_183 V144 V183 -256.7711732710434
L144_183 V144 V183 -7.639136215944605e-12
C144_183 V144 V183 -3.5859043738820054e-20

R144_184 V144 V184 -513.9875079600521
L144_184 V144 V184 1.1554880955657387e-11
C144_184 V144 V184 -1.6724757944363554e-20

R144_185 V144 V185 -11959.520320200312
L144_185 V144 V185 6.184516968710483e-12
C144_185 V144 V185 1.1985409821010372e-19

R144_186 V144 V186 -135.00327599204587
L144_186 V144 V186 -8.53579168799986e-12
C144_186 V144 V186 -3.3427833586750633e-20

R144_187 V144 V187 -462.2981865363409
L144_187 V144 V187 1.6946099385763864e-11
C144_187 V144 V187 -1.514762726139899e-20

R144_188 V144 V188 171.35406362278576
L144_188 V144 V188 2.8889931393258416e-12
C144_188 V144 V188 1.0974273112277863e-19

R144_189 V144 V189 212.81735714891212
L144_189 V144 V189 -2.7931915097829738e-11
C144_189 V144 V189 5.588371153948914e-20

R144_190 V144 V190 74.81193662569089
L144_190 V144 V190 5.058519032008743e-12
C144_190 V144 V190 -5.630840306293013e-20

R144_191 V144 V191 118.4891037845108
L144_191 V144 V191 3.7791435037774305e-12
C144_191 V144 V191 1.416326717864157e-19

R144_192 V144 V192 -137.26892327728115
L144_192 V144 V192 -2.326202167872582e-12
C144_192 V144 V192 -9.509057591024061e-20

R144_193 V144 V193 -1085.0852054468896
L144_193 V144 V193 3.209028699066202e-11
C144_193 V144 V193 -4.963966554705974e-20

R144_194 V144 V194 -351.722442684486
L144_194 V144 V194 -8.409072566654564e-12
C144_194 V144 V194 3.145929382209109e-20

R144_195 V144 V195 -461.02997420207146
L144_195 V144 V195 -3.7558550100848124e-12
C144_195 V144 V195 -2.9457418674690606e-19

R144_196 V144 V196 752.5696692695382
L144_196 V144 V196 3.4446569489649707e-12
C144_196 V144 V196 2.478111769281412e-19

R144_197 V144 V197 -202.42384409283645
L144_197 V144 V197 -7.259211789263279e-12
C144_197 V144 V197 -1.225496268329386e-19

R144_198 V144 V198 -331.72204375167064
L144_198 V144 V198 -5.125185554338955e-12
C144_198 V144 V198 -2.500531533895409e-21

R144_199 V144 V199 122.77056479598419
L144_199 V144 V199 -8.910458229964102e-12
C144_199 V144 V199 5.3978363970865544e-20

R144_200 V144 V200 746.024172711006
L144_200 V144 V200 3.8997624580762936e-12
C144_200 V144 V200 -1.3958291562122346e-19

R145_145 V145 0 -29.95389648521652
L145_145 V145 0 2.1198013102837466e-13
C145_145 V145 0 1.1680685123989946e-18

R145_146 V145 V146 -187.6918469740648
L145_146 V145 V146 -3.549055370644224e-12
C145_146 V145 V146 -4.385167353489466e-20

R145_147 V145 V147 790.0770308170173
L145_147 V145 V147 8.002003231528951e-12
C145_147 V145 V147 -1.344537673616624e-19

R145_148 V145 V148 54.478126369716875
L145_148 V145 V148 5.571467421033567e-12
C145_148 V145 V148 4.830391775142199e-20

R145_149 V145 V149 34.41989209161124
L145_149 V145 V149 4.867267299486783e-13
C145_149 V145 V149 8.568044043072038e-19

R145_150 V145 V150 11.343313440250812
L145_150 V145 V150 2.243316369359656e-12
C145_150 V145 V150 -4.3329726928340282e-19

R145_151 V145 V151 26.30645225382627
L145_151 V145 V151 5.1797706976520586e-12
C145_151 V145 V151 1.1590464761762423e-19

R145_152 V145 V152 71.01203022746891
L145_152 V145 V152 3.446407734457498e-12
C145_152 V145 V152 -3.453431303651833e-20

R145_153 V145 V153 18.886990292000355
L145_153 V145 V153 6.297736048680517e-13
C145_153 V145 V153 3.1050670845297332e-19

R145_154 V145 V154 340.32146790200244
L145_154 V145 V154 1.9846054638753822e-12
C145_154 V145 V154 3.8098759375754967e-19

R145_155 V145 V155 -32.22422659881744
L145_155 V145 V155 2.2527933148338756e-12
C145_155 V145 V155 1.2856751399580227e-19

R145_156 V145 V156 78.76991968972216
L145_156 V145 V156 5.203103604017703e-12
C145_156 V145 V156 6.852404013375523e-20

R145_157 V145 V157 118.74233872447245
L145_157 V145 V157 -1.0536998553292304e-12
C145_157 V145 V157 -6.302537800219107e-19

R145_158 V145 V158 -18.88481331520806
L145_158 V145 V158 -3.450139997055387e-12
C145_158 V145 V158 2.1116114226975022e-20

R145_159 V145 V159 -269.4724738909967
L145_159 V145 V159 -4.03321642865366e-12
C145_159 V145 V159 1.0288686777699314e-19

R145_160 V145 V160 -35.65360830502918
L145_160 V145 V160 -2.5306532674663554e-11
C145_160 V145 V160 1.5747068172600795e-19

R145_161 V145 V161 -27.904324638490095
L145_161 V145 V161 -1.0331469660609162e-12
C145_161 V145 V161 -3.1145093323076366e-19

R145_162 V145 V162 -89.11438212622669
L145_162 V145 V162 -1.4259877168793065e-10
C145_162 V145 V162 8.062211571718735e-20

R145_163 V145 V163 -248.3856039887407
L145_163 V145 V163 -1.2897620214779834e-11
C145_163 V145 V163 -1.109436534613664e-19

R145_164 V145 V164 -930.6835456139903
L145_164 V145 V164 -3.1672046817620972e-12
C145_164 V145 V164 -1.0717438935526418e-19

R145_165 V145 V165 -165.65073406871514
L145_165 V145 V165 -5.273039196630553e-12
C145_165 V145 V165 4.844480401797989e-19

R145_166 V145 V166 12.599613160078928
L145_166 V145 V166 -1.9215854190076974e-11
C145_166 V145 V166 -1.7190432290370847e-19

R145_167 V145 V167 70.40308685739963
L145_167 V145 V167 -5.098842455164643e-12
C145_167 V145 V167 -1.3182573710134953e-19

R145_168 V145 V168 -170.34819330791882
L145_168 V145 V168 -3.984906356359378e-12
C145_168 V145 V168 -2.587719571577595e-19

R145_169 V145 V169 30.91772888070639
L145_169 V145 V169 9.103887407947935e-13
C145_169 V145 V169 1.5300859830493007e-19

R145_170 V145 V170 -25.191708908820207
L145_170 V145 V170 -4.462567821563423e-12
C145_170 V145 V170 2.099769947820617e-19

R145_171 V145 V171 -101.19955792381735
L145_171 V145 V171 6.191852648316758e-12
C145_171 V145 V171 2.5268540093870435e-19

R145_172 V145 V172 -329.7493467294225
L145_172 V145 V172 2.7010260157298693e-12
C145_172 V145 V172 2.6503676403712803e-19

R145_173 V145 V173 -54.16362770905244
L145_173 V145 V173 -2.2298685135793596e-12
C145_173 V145 V173 -2.246804741152319e-19

R145_174 V145 V174 -23.847599745785534
L145_174 V145 V174 1.3538593870523615e-12
C145_174 V145 V174 5.020327368385096e-20

R145_175 V145 V175 261.25097006871465
L145_175 V145 V175 1.5486917145366882e-12
C145_175 V145 V175 1.7546697792991022e-19

R145_176 V145 V176 121.0315191806695
L145_176 V145 V176 1.8527334875554335e-12
C145_176 V145 V176 8.832495584492632e-20

R145_177 V145 V177 -141.149446725841
L145_177 V145 V177 -3.1785310271179866e-12
C145_177 V145 V177 -2.2138607357086235e-21

R145_178 V145 V178 28.30538686724783
L145_178 V145 V178 -1.0061509939055161e-11
C145_178 V145 V178 -2.0867756545502786e-19

R145_179 V145 V179 -135.16411396844046
L145_179 V145 V179 -1.982728773788044e-12
C145_179 V145 V179 -3.34482468332324e-19

R145_180 V145 V180 -232.2736930694168
L145_180 V145 V180 -1.6334076384434634e-12
C145_180 V145 V180 -2.308058401761562e-19

R145_181 V145 V181 63.12033722485886
L145_181 V145 V181 1.6519459638745485e-11
C145_181 V145 V181 -1.7924243704410632e-19

R145_182 V145 V182 54.38426022951734
L145_182 V145 V182 6.084789003207263e-12
C145_182 V145 V182 2.005378724688801e-19

R145_183 V145 V183 295.3872765083063
L145_183 V145 V183 -4.158380560797981e-12
C145_183 V145 V183 1.4556088610577094e-20

R145_184 V145 V184 -158.1219764911
L145_184 V145 V184 -3.39231708947016e-12
C145_184 V145 V184 -1.056431540531055e-20

R145_185 V145 V185 -269.61702310167436
L145_185 V145 V185 -2.8758718015082994e-12
C145_185 V145 V185 1.9575296999379199e-19

R145_186 V145 V186 -82.28538094814449
L145_186 V145 V186 -2.8317629039921e-12
C145_186 V145 V186 -5.0870620050198743e-20

R145_187 V145 V187 -499.84472776171566
L145_187 V145 V187 4.675459524607658e-12
C145_187 V145 V187 1.646911242036423e-19

R145_188 V145 V188 315.1574057451551
L145_188 V145 V188 4.2551425232649613e-11
C145_188 V145 V188 7.337106273774357e-20

R145_189 V145 V189 -21478.967224740874
L145_189 V145 V189 9.781311749187314e-13
C145_189 V145 V189 1.8194349393551693e-19

R145_190 V145 V190 1124.2178630723668
L145_190 V145 V190 7.868540047491544e-12
C145_190 V145 V190 -2.1201968172343867e-19

R145_191 V145 V191 275.9689576435123
L145_191 V145 V191 3.7103701947742935e-12
C145_191 V145 V191 6.697824163214605e-20

R145_192 V145 V192 -1392.5040414140335
L145_192 V145 V192 1.4062446361884152e-12
C145_192 V145 V192 2.195916354566995e-19

R145_193 V145 V193 1320.2640240651253
L145_193 V145 V193 -2.4720170761394038e-11
C145_193 V145 V193 -1.1637814669194536e-19

R145_194 V145 V194 1324.153730372756
L145_194 V145 V194 1.3602963809627647e-12
C145_194 V145 V194 2.230101959343521e-19

R145_195 V145 V195 -437.8023720102463
L145_195 V145 V195 -3.2517514917235283e-12
C145_195 V145 V195 -1.3569544480615482e-19

R145_196 V145 V196 322.9401660014935
L145_196 V145 V196 -2.2809337560178696e-12
C145_196 V145 V196 -3.416230362857764e-19

R145_197 V145 V197 -177.54402641707597
L145_197 V145 V197 -1.3551978197306774e-12
C145_197 V145 V197 -2.773955293979308e-19

R145_198 V145 V198 50.25546240698652
L145_198 V145 V198 -3.99841887842473e-12
C145_198 V145 V198 4.9215759053684133e-20

R145_199 V145 V199 78.15906257146922
L145_199 V145 V199 -3.642709176416444e-12
C145_199 V145 V199 -5.419574408504751e-20

R145_200 V145 V200 -111.99005847981951
L145_200 V145 V200 -1.9723272059569068e-12
C145_200 V145 V200 -1.0113899198600365e-19

R146_146 V146 0 29.127555611950047
L146_146 V146 0 -2.101888087576254e-12
C146_146 V146 0 -3.472159288954284e-19

R146_147 V146 V147 -83.83405248338158
L146_147 V146 V147 3.3897795731224073e-12
C146_147 V146 V147 2.7133292815178946e-19

R146_148 V146 V148 -68.99761534622168
L146_148 V146 V148 1.6172813468353981e-12
C146_148 V146 V148 2.77380647972586e-19

R146_149 V146 V149 -894.2452552493759
L146_149 V146 V149 5.636332166487331e-13
C146_149 V146 V149 2.464882451580212e-19

R146_150 V146 V150 81.60095699367078
L146_150 V146 V150 3.0644669080522954e-11
C146_150 V146 V150 -8.32907156698228e-20

R146_151 V146 V151 59.138929141549106
L146_151 V146 V151 3.0923562456713443e-12
C146_151 V146 V151 -5.5312859691093745e-21

R146_152 V146 V152 39.88391486347338
L146_152 V146 V152 -5.22434484062299e-12
C146_152 V146 V152 -1.167085364089737e-19

R146_153 V146 V153 136.62250980256786
L146_153 V146 V153 -2.014446654204795e-11
C146_153 V146 V153 -5.907459909865917e-20

R146_154 V146 V154 18.158729801421035
L146_154 V146 V154 8.266466773009558e-13
C146_154 V146 V154 2.403527622051175e-19

R146_155 V146 V155 -996.8967289579637
L146_155 V146 V155 -4.515172400857605e-12
C146_155 V146 V155 -1.3953068833833448e-19

R146_156 V146 V156 -131.4059994212268
L146_156 V146 V156 -7.317773774273538e-11
C146_156 V146 V156 -1.2231009068888715e-19

R146_157 V146 V157 49.34671976406695
L146_157 V146 V157 -9.15136532286106e-13
C146_157 V146 V157 -2.5059591870293414e-19

R146_158 V146 V158 -37.17874910455895
L146_158 V146 V158 2.8905001726062192e-12
C146_158 V146 V158 -4.2739557916598435e-20

R146_159 V146 V159 -50.429255253302195
L146_159 V146 V159 -1.3996502309948117e-11
C146_159 V146 V159 1.219914931769857e-19

R146_160 V146 V160 -43.00417228085512
L146_160 V146 V160 -2.2189148710924894e-09
C146_160 V146 V160 1.4130818814924145e-19

R146_161 V146 V161 256.7458932933293
L146_161 V146 V161 -2.027717048172726e-12
C146_161 V146 V161 -4.8117986802392934e-20

R146_162 V146 V162 -21.78160085041183
L146_162 V146 V162 -1.0910250264920793e-12
C146_162 V146 V162 -1.1771943051296922e-19

R146_163 V146 V163 69.36270278534292
L146_163 V146 V163 -2.092890223670912e-12
C146_163 V146 V163 -2.121157650779828e-19

R146_164 V146 V164 42.15009331170222
L146_164 V146 V164 -4.0479789097288046e-11
C146_164 V146 V164 -1.5424505739167976e-19

R146_165 V146 V165 -38.11220965977107
L146_165 V146 V165 7.270574986137959e-13
C146_165 V146 V165 3.853273707647904e-19

R146_166 V146 V166 20.909948324002897
L146_166 V146 V166 1.8030891764076244e-12
C146_166 V146 V166 1.0321511477657184e-19

R146_167 V146 V167 -71.8308603927003
L146_167 V146 V167 -2.946343827020485e-12
C146_167 V146 V167 2.1767421590945578e-20

R146_168 V146 V168 -41.37212957506098
L146_168 V146 V168 -1.1027536790089151e-12
C146_168 V146 V168 -1.8507770805879123e-20

R146_169 V146 V169 -132.08497236322597
L146_169 V146 V169 1.5702361907214557e-11
C146_169 V146 V169 4.2320197660898453e-20

R146_170 V146 V170 528.8371080765531
L146_170 V146 V170 1.9867385332855164e-12
C146_170 V146 V170 9.130100011185295e-20

R146_171 V146 V171 -768.2618077822273
L146_171 V146 V171 8.807610548862516e-13
C146_171 V146 V171 2.470966773799358e-19

R146_172 V146 V172 174.54121400940036
L146_172 V146 V172 7.253944399423593e-13
C146_172 V146 V172 1.889536458715863e-19

R146_173 V146 V173 39.40131869434116
L146_173 V146 V173 -1.3813969920189344e-12
C146_173 V146 V173 -3.0844360420046155e-19

R146_174 V146 V174 -20.88541384459205
L146_174 V146 V174 -1.2083572785396035e-12
C146_174 V146 V174 -1.495666144110759e-19

R146_175 V146 V175 97.436388339075
L146_175 V146 V175 -3.5249289807154305e-10
C146_175 V146 V175 -1.5384945264734285e-19

R146_176 V146 V176 49.52509897160574
L146_176 V146 V176 -2.395658336017121e-12
C146_176 V146 V176 -2.450542398058025e-19

R146_177 V146 V177 -175.6677213981961
L146_177 V146 V177 3.0996017500974773e-12
C146_177 V146 V177 1.4155167147672706e-19

R146_178 V146 V178 52.10195905802815
L146_178 V146 V178 -4.8248468244967646e-12
C146_178 V146 V178 -3.234236972232484e-20

R146_179 V146 V179 -222.5672800666996
L146_179 V146 V179 -1.176647766560057e-12
C146_179 V146 V179 -7.823106428398378e-20

R146_180 V146 V180 -39.48870733000089
L146_180 V146 V180 -1.0472426921925528e-12
C146_180 V146 V180 3.4858895908273586e-20

R146_181 V146 V181 -94.44845627120554
L146_181 V146 V181 -4.075702539843941e-12
C146_181 V146 V181 8.187887137579547e-20

R146_182 V146 V182 64.41939523898054
L146_182 V146 V182 6.950555858996543e-13
C146_182 V146 V182 1.391665708613682e-19

R146_183 V146 V183 -409.5010806828184
L146_183 V146 V183 -1.9111875168292257e-11
C146_183 V146 V183 8.593824434141635e-21

R146_184 V146 V184 131.33335617926414
L146_184 V146 V184 2.0718456021501617e-12
C146_184 V146 V184 6.786317759259898e-21

R146_185 V146 V185 81.4129877769135
L146_185 V146 V185 2.1390269019876927e-11
C146_185 V146 V185 -1.119766141264689e-19

R146_186 V146 V186 -72.77689259692477
L146_186 V146 V186 3.0414066950940873e-12
C146_186 V146 V186 6.036336383300235e-20

R146_187 V146 V187 2369.91383927661
L146_187 V146 V187 1.842721809529315e-12
C146_187 V146 V187 9.148812564191382e-21

R146_188 V146 V188 83.46958053635711
L146_188 V146 V188 -1.7639249175307227e-11
C146_188 V146 V188 2.973303705902724e-20

R146_189 V146 V189 -301.02018532327577
L146_189 V146 V189 1.7461378427388154e-12
C146_189 V146 V189 1.3511817054839181e-19

R146_190 V146 V190 -85.9239669581497
L146_190 V146 V190 -1.5925472713269984e-12
C146_190 V146 V190 -1.0198386917705247e-19

R146_191 V146 V191 12228.93731179016
L146_191 V146 V191 2.9567095694310574e-12
C146_191 V146 V191 1.8370836027827936e-19

R146_192 V146 V192 -129.61488429835842
L146_192 V146 V192 1.5199046441194307e-12
C146_192 V146 V192 1.7679310179321647e-19

R146_193 V146 V193 -157.28713080844054
L146_193 V146 V193 -2.0572276073650024e-12
C146_193 V146 V193 -8.552195775687688e-20

R146_194 V146 V194 184.78815873121772
L146_194 V146 V194 2.07503915038299e-12
C146_194 V146 V194 1.0050657413029256e-19

R146_195 V146 V195 589.7795810744531
L146_195 V146 V195 -1.383788849262679e-12
C146_195 V146 V195 -2.1547547498193364e-19

R146_196 V146 V196 379.11030548177564
L146_196 V146 V196 -5.676102241064124e-13
C146_196 V146 V196 -4.1481136655657496e-19

R146_197 V146 V197 88.63664610898861
L146_197 V146 V197 -1.6784788349054546e-12
C146_197 V146 V197 -8.161131828752311e-20

R146_198 V146 V198 94.88829713519809
L146_198 V146 V198 3.253298636556204e-12
C146_198 V146 V198 4.5658628440345006e-20

R146_199 V146 V199 831.1834741938679
L146_199 V146 V199 -1.568561875776085e-12
C146_199 V146 V199 -1.6525474146554362e-19

R146_200 V146 V200 169.7094981994147
L146_200 V146 V200 -2.985628622218551e-11
C146_200 V146 V200 -3.4173069752228484e-22

R147_147 V147 0 133.59626504619365
L147_147 V147 0 9.537207483830385e-13
C147_147 V147 0 4.226348775968419e-19

R147_148 V147 V148 137.1896025162813
L147_148 V147 V148 2.713449470140752e-12
C147_148 V147 V148 -5.690903298743288e-20

R147_149 V147 V149 522.1456491849887
L147_149 V147 V149 4.275537274962644e-12
C147_149 V147 V149 3.1764925211051433e-19

R147_150 V147 V150 64.93631160487192
L147_150 V147 V150 -1.0248331298853657e-11
C147_150 V147 V150 1.2933614991547671e-19

R147_151 V147 V151 -79.41035907470602
L147_151 V147 V151 -5.5751613212947085e-12
C147_151 V147 V151 7.310557278558944e-19

R147_152 V147 V152 133.40629179458222
L147_152 V147 V152 -1.6914850113051053e-11
C147_152 V147 V152 -2.552633256358161e-20

R147_153 V147 V153 751.1848902650187
L147_153 V147 V153 2.951845256304262e-11
C147_153 V147 V153 -1.2116568602272884e-19

R147_154 V147 V154 194.55908895089715
L147_154 V147 V154 3.80912148777917e-11
C147_154 V147 V154 -2.729112314389565e-19

R147_155 V147 V155 52.21654962046041
L147_155 V147 V155 4.70452039931624e-13
C147_155 V147 V155 3.900216029853923e-19

R147_156 V147 V156 -427.17382078017226
L147_156 V147 V156 -7.415106721929209e-12
C147_156 V147 V156 -4.2824705392992185e-20

R147_157 V147 V157 471.7392302230364
L147_157 V147 V157 4.947578365698375e-11
C147_157 V147 V157 1.1752637117123324e-20

R147_158 V147 V158 -57.34782286945678
L147_158 V147 V158 -7.237940215488109e-12
C147_158 V147 V158 1.9956223314343492e-19

R147_159 V147 V159 33.151490979042755
L147_159 V147 V159 -2.5228805259234984e-12
C147_159 V147 V159 -6.3476790859035685e-19

R147_160 V147 V160 -57.12012371870631
L147_160 V147 V160 -6.904685571585691e-12
C147_160 V147 V160 7.267381775207202e-20

R147_161 V147 V161 -260.8053072447237
L147_161 V147 V161 9.581369628765286e-12
C147_161 V147 V161 1.8360888680039669e-19

R147_162 V147 V162 -105.80749176137016
L147_162 V147 V162 5.858316891334766e-12
C147_162 V147 V162 2.5902341491579903e-19

R147_163 V147 V163 -48.9387022564137
L147_163 V147 V163 -1.6799589030365932e-12
C147_163 V147 V163 4.921976470495983e-19

R147_164 V147 V164 101.65911958405691
L147_164 V147 V164 1.2045241186627174e-11
C147_164 V147 V164 1.2136143028712165e-19

R147_165 V147 V165 -544.6379696575912
L147_165 V147 V165 -1.6928494517288435e-12
C147_165 V147 V165 -3.222732535002515e-19

R147_166 V147 V166 35.08607203627504
L147_166 V147 V166 -3.100036629284388e-11
C147_166 V147 V166 -1.7633005771117684e-19

R147_167 V147 V167 -67.18808898479136
L147_167 V147 V167 2.8992171541181245e-12
C147_167 V147 V167 9.874417897934588e-20

R147_168 V147 V168 -356.51672644271883
L147_168 V147 V168 4.5494406090706177e-11
C147_168 V147 V168 1.7050747373782315e-20

R147_169 V147 V169 307.63647943869285
L147_169 V147 V169 -7.176789736230189e-12
C147_169 V147 V169 -2.2382648377367553e-19

R147_170 V147 V170 -122.2224332157031
L147_170 V147 V170 -5.6792810770919545e-12
C147_170 V147 V170 -5.073298087084847e-20

R147_171 V147 V171 78.33678391797703
L147_171 V147 V171 -5.771198327435704e-12
C147_171 V147 V171 -4.994070825086288e-19

R147_172 V147 V172 2143.1855322671195
L147_172 V147 V172 -1.4043758738611367e-11
C147_172 V147 V172 -2.0020577737517404e-19

R147_173 V147 V173 -305.00367822935937
L147_173 V147 V173 1.5934681682897968e-12
C147_173 V147 V173 3.9261900617258256e-19

R147_174 V147 V174 -40.865294063850165
L147_174 V147 V174 5.881752645236364e-12
C147_174 V147 V174 9.095064868390944e-20

R147_175 V147 V175 155.82306372538653
L147_175 V147 V175 2.111237435827164e-12
C147_175 V147 V175 7.233873299853289e-19

R147_176 V147 V176 260.1711734484906
L147_176 V147 V176 2.524124630858849e-10
C147_176 V147 V176 3.4792504795081216e-21

R147_177 V147 V177 561.2220782003469
L147_177 V147 V177 -3.3752029911594613e-12
C147_177 V147 V177 -1.6219965675304967e-19

R147_178 V147 V178 73.67197905387278
L147_178 V147 V178 3.911043490694048e-11
C147_178 V147 V178 8.682831876361592e-21

R147_179 V147 V179 -116.59132274139318
L147_179 V147 V179 -6.176754058279935e-12
C147_179 V147 V179 -4.457163205602571e-19

R147_180 V147 V180 -127.10325856679651
L147_180 V147 V180 -6.84578013274889e-10
C147_180 V147 V180 6.996350442576147e-20

R147_181 V147 V181 -775.725237794735
L147_181 V147 V181 -5.4188705323701214e-11
C147_181 V147 V181 -4.746163511000273e-20

R147_182 V147 V182 122.15128279168898
L147_182 V147 V182 -2.4328860941523278e-11
C147_182 V147 V182 3.053492137118958e-20

R147_183 V147 V183 449.64950070360794
L147_183 V147 V183 -1.1502588443120813e-11
C147_183 V147 V183 5.945719108251116e-20

R147_184 V147 V184 208.52412191933826
L147_184 V147 V184 -1.1311861198587797e-11
C147_184 V147 V184 -1.5874073629785895e-19

R147_185 V147 V185 -1883.826018015716
L147_185 V147 V185 5.856901641364322e-12
C147_185 V147 V185 1.7233095114546292e-19

R147_186 V147 V186 -243.5971490821497
L147_186 V147 V186 -4.134440218623067e-12
C147_186 V147 V186 -2.0718621157827617e-19

R147_187 V147 V187 -186.67019475504415
L147_187 V147 V187 5.483328688779065e-12
C147_187 V147 V187 4.494418890778154e-19

R147_188 V147 V188 850.9516877728593
L147_188 V147 V188 2.1769224186949223e-11
C147_188 V147 V188 6.55559778843291e-20

R147_189 V147 V189 438.1299850477294
L147_189 V147 V189 -1.5657852976513663e-11
C147_189 V147 V189 -2.2965318411371326e-19

R147_190 V147 V190 -196.57926693928297
L147_190 V147 V190 1.5019911307451363e-11
C147_190 V147 V190 1.0472366541228957e-19

R147_191 V147 V191 -847.2083622512222
L147_191 V147 V191 -5.929208319254444e-12
C147_191 V147 V191 -5.836073574389659e-19

R147_192 V147 V192 -131.25132392646944
L147_192 V147 V192 5.7351031100854584e-12
C147_192 V147 V192 -3.1211059120044706e-20

R147_193 V147 V193 -372.2724812398992
L147_193 V147 V193 7.132600815212872e-11
C147_193 V147 V193 8.375252367051134e-20

R147_194 V147 V194 -975.0052836094925
L147_194 V147 V194 1.1600935050202652e-11
C147_194 V147 V194 -1.625332624394271e-19

R147_195 V147 V195 115.12057366668047
L147_195 V147 V195 1.9865052949029663e-12
C147_195 V147 V195 8.797258112667947e-19

R147_196 V147 V196 173.46770146685213
L147_196 V147 V196 -2.7359783687415003e-12
C147_196 V147 V196 -1.7821250621331424e-19

R147_197 V147 V197 2541.101091955641
L147_197 V147 V197 7.481570401369174e-12
C147_197 V147 V197 1.1707422289953432e-19

R147_198 V147 V198 119.88862662857534
L147_198 V147 V198 -2.8537218545167877e-11
C147_198 V147 V198 2.676935203410294e-20

R147_199 V147 V199 -1934.3977097759246
L147_199 V147 V199 1.4849581354780107e-11
C147_199 V147 V199 1.9673944722555332e-19

R147_200 V147 V200 1281.511249963291
L147_200 V147 V200 2.8943156007817584e-12
C147_200 V147 V200 2.710516025084517e-19

R148_148 V148 0 15.824297127045114
L148_148 V148 0 2.1373850531132565e-13
C148_148 V148 0 2.0411885053315066e-18

R148_149 V148 V149 -449.2563566301461
L148_149 V148 V149 9.40582789652589e-13
C148_149 V148 V149 8.498817377017638e-20

R148_150 V148 V150 -468.7532845313059
L148_150 V148 V150 -2.391589879819632e-12
C148_150 V148 V150 -1.2790938236931043e-19

R148_151 V148 V151 47.91567321839352
L148_151 V148 V151 3.0187391321875715e-12
C148_151 V148 V151 -4.643029180193797e-20

R148_152 V148 V152 -44.15992399694666
L148_152 V148 V152 8.485396686364473e-13
C148_152 V148 V152 4.4305964628622125e-19

R148_153 V148 V153 -93.16360264899946
L148_153 V148 V153 1.914697527538509e-12
C148_153 V148 V153 8.559633681414433e-20

R148_154 V148 V154 128.58112434353072
L148_154 V148 V154 2.1715086195619526e-12
C148_154 V148 V154 -1.2265205501321098e-19

R148_155 V148 V155 -43.57286827089444
L148_155 V148 V155 -1.6629060384617887e-11
C148_155 V148 V155 -9.914706437418775e-20

R148_156 V148 V156 39.06111663165502
L148_156 V148 V156 7.628800245633636e-13
C148_156 V148 V156 7.06378807489421e-19

R148_157 V148 V157 -200.80350135771928
L148_157 V148 V157 -7.049601117041309e-13
C148_157 V148 V157 -3.255570152816457e-19

R148_158 V148 V158 -51.8649825490568
L148_158 V148 V158 -3.520137202874635e-12
C148_158 V148 V158 1.0363930272573572e-19

R148_159 V148 V159 -31.385790658404233
L148_159 V148 V159 4.5854610642640115e-12
C148_159 V148 V159 2.0014295265908495e-19

R148_160 V148 V160 13.92856305661233
L148_160 V148 V160 -1.7070687845658155e-11
C148_160 V148 V160 -5.527567662881226e-19

R148_161 V148 V161 415.32949826863836
L148_161 V148 V161 1.4754363638677134e-12
C148_161 V148 V161 1.9319368102642812e-19

R148_162 V148 V162 -142.46634100036724
L148_162 V148 V162 1.952172502172894e-12
C148_162 V148 V162 9.172811609925164e-20

R148_163 V148 V163 63.622397922570784
L148_163 V148 V163 2.6370254026144158e-11
C148_163 V148 V163 -8.627116386743135e-20

R148_164 V148 V164 -17.445306698251052
L148_164 V148 V164 -1.3499492790332419e-12
C148_164 V148 V164 3.7259738840039443e-19

R148_165 V148 V165 -114.73259050400652
L148_165 V148 V165 -2.164272507700146e-12
C148_165 V148 V165 -2.1390653172001359e-19

R148_166 V148 V166 51.31465087979698
L148_166 V148 V166 -2.7295979310192225e-12
C148_166 V148 V166 -2.725486284634495e-19

R148_167 V148 V167 284.58185044379996
L148_167 V148 V167 -1.5938420374833296e-11
C148_167 V148 V167 8.372767117409181e-20

R148_168 V148 V168 -52.027656429577895
L148_168 V148 V168 1.413504386187403e-12
C148_168 V148 V168 -4.034296119275223e-20

R148_169 V148 V169 -691.4964714646306
L148_169 V148 V169 -1.163950784186014e-10
C148_169 V148 V169 -2.7482972611979266e-19

R148_170 V148 V170 -108.75270612537787
L148_170 V148 V170 3.078118283104932e-12
C148_170 V148 V170 3.7207094196755476e-20

R148_171 V148 V171 -88.09068387122834
L148_171 V148 V171 1.4689788012664478e-12
C148_171 V148 V171 -9.709265474679022e-20

R148_172 V148 V172 29.019783772221675
L148_172 V148 V172 -9.63297544344543e-13
C148_172 V148 V172 -1.533516727385459e-19

R148_173 V148 V173 -2926.2413964250936
L148_173 V148 V173 2.1511096265327858e-12
C148_173 V148 V173 2.8164684540367164e-19

R148_174 V148 V174 -70.65346431088814
L148_174 V148 V174 -1.7964469537632818e-11
C148_174 V148 V174 1.6649708252518654e-20

R148_175 V148 V175 269.4483308819681
L148_175 V148 V175 -1.4119473641612924e-12
C148_175 V148 V175 -7.26721629087626e-20

R148_176 V148 V176 399.19995933755945
L148_176 V148 V176 5.90651305413022e-13
C148_176 V148 V176 7.556278966400878e-19

R148_177 V148 V177 -171.57558597252088
L148_177 V148 V177 -2.5419552129317268e-12
C148_177 V148 V177 -1.2562716149035946e-19

R148_178 V148 V178 97.5169743745219
L148_178 V148 V178 -3.9023358273354985e-12
C148_178 V148 V178 2.3919780802747917e-20

R148_179 V148 V179 -1496.1959405906732
L148_179 V148 V179 -2.606946043635992e-12
C148_179 V148 V179 1.7806936335608536e-20

R148_180 V148 V180 -98.44366884640293
L148_180 V148 V180 -1.2350055999366733e-12
C148_180 V148 V180 -5.585176871917208e-19

R148_181 V148 V181 259.09175863940555
L148_181 V148 V181 -2.6112776110441017e-11
C148_181 V148 V181 -6.716715781997192e-20

R148_182 V148 V182 92.38930634872052
L148_182 V148 V182 6.536163078287567e-12
C148_182 V148 V182 -8.246539725968083e-20

R148_183 V148 V183 160.81991135179126
L148_183 V148 V183 -7.042859188071657e-12
C148_183 V148 V183 -1.3514587940559662e-19

R148_184 V148 V184 691.3307098404266
L148_184 V148 V184 -1.229456470699296e-12
C148_184 V148 V184 1.5895459925032347e-19

R148_185 V148 V185 801.8870950841762
L148_185 V148 V185 6.891253094799673e-12
C148_185 V148 V185 1.3432361414591345e-19

R148_186 V148 V186 3709.344477684852
L148_186 V148 V186 -1.9152213074286594e-12
C148_186 V148 V186 4.08667618244067e-20

R148_187 V148 V187 182.07474435949882
L148_187 V148 V187 -3.324584164614788e-12
C148_187 V148 V187 1.231996354501405e-19

R148_188 V148 V188 -183.75873973469345
L148_188 V148 V188 4.796018369720582e-13
C148_188 V148 V188 1.4455879992128278e-19

R148_189 V148 V189 -657.9760647384675
L148_189 V148 V189 -2.117469685140106e-11
C148_189 V148 V189 -1.1251010500429182e-19

R148_190 V148 V190 -87.12030014133839
L148_190 V148 V190 7.082630474480796e-12
C148_190 V148 V190 -1.0183516116823107e-20

R148_191 V148 V191 -75.60179826205281
L148_191 V148 V191 8.92816738703134e-13
C148_191 V148 V191 1.2715146670980972e-19

R148_192 V148 V192 93.52812323879031
L148_192 V148 V192 -8.534341597886649e-13
C148_192 V148 V192 -4.683244722278628e-19

R148_193 V148 V193 339.11079698793424
L148_193 V148 V193 -1.3595582822746736e-11
C148_193 V148 V193 -5.055729046905787e-20

R148_194 V148 V194 -739.4358540627693
L148_194 V148 V194 -2.5672799340727564e-12
C148_194 V148 V194 -3.579194863609656e-19

R148_195 V148 V195 491.17923962353717
L148_195 V148 V195 -5.943427623296105e-13
C148_195 V148 V195 -5.897677696819087e-19

R148_196 V148 V196 -210.47393311786774
L148_196 V148 V196 6.290460134915988e-13
C148_196 V148 V196 1.1059540728073068e-18

R148_197 V148 V197 155.5266492570774
L148_197 V148 V197 -2.8975617153374016e-11
C148_197 V148 V197 1.6082632329350477e-19

R148_198 V148 V198 813.2122960779084
L148_198 V148 V198 7.939444736378007e-11
C148_198 V148 V198 -1.3219206440246233e-19

R148_199 V148 V199 -102.4681227709471
L148_199 V148 V199 3.0946775313914918e-12
C148_199 V148 V199 1.2307431582635868e-19

R148_200 V148 V200 165.19671966907072
L148_200 V148 V200 -1.4077747169549166e-12
C148_200 V148 V200 -1.8308641349032e-19

R149_149 V149 0 400.1856255529641
L149_149 V149 0 -1.1306339666119227e-13
C149_149 V149 0 -5.214585708057275e-18

R149_150 V149 V150 -28.378238477836952
L149_150 V149 V150 -1.767135971804358e-11
C149_150 V149 V150 1.6975328745357715e-18

R149_151 V149 V151 -76.15000847140318
L149_151 V149 V151 -1.4298839380805598e-12
C149_151 V149 V151 -5.868639893671364e-19

R149_152 V149 V152 -94.81765790150676
L149_152 V149 V152 -2.1913800291786752e-12
C149_152 V149 V152 8.754880605800226e-20

R149_153 V149 V153 -605.6415209560106
L149_153 V149 V153 -1.183395794543416e-12
C149_153 V149 V153 -2.686484518457404e-19

R149_154 V149 V154 127.8673882914488
L149_154 V149 V154 -1.3871392857322567e-12
C149_154 V149 V154 -1.453840752925659e-18

R149_155 V149 V155 85.98125835818834
L149_155 V149 V155 -4.964096440241753e-13
C149_155 V149 V155 -6.636929369946962e-19

R149_156 V149 V156 168.6486363467331
L149_156 V149 V156 -2.3997227990304096e-12
C149_156 V149 V156 -4.391143302934217e-19

R149_157 V149 V157 37.48473177764513
L149_157 V149 V157 1.5420882825716536e-13
C149_157 V149 V157 2.9741347768764735e-18

R149_158 V149 V158 48.49426679044157
L149_158 V149 V158 -1.8439504105723423e-12
C149_158 V149 V158 2.782975178050418e-20

R149_159 V149 V159 210.31842124028046
L149_159 V149 V159 1.2958074629475094e-12
C149_159 V149 V159 2.371227339176839e-20

R149_160 V149 V160 121.4203131366684
L149_160 V149 V160 -1.5257457053785854e-12
C149_160 V149 V160 -2.756453668171866e-19

R149_161 V149 V161 2169.921669881271
L149_161 V149 V161 3.2467386074295743e-12
C149_161 V149 V161 4.60051729108521e-19

R149_162 V149 V162 -75.90515787110922
L149_162 V149 V162 -9.271538764211722e-13
C149_162 V149 V162 -2.380615437041125e-19

R149_163 V149 V163 -73.4187804506724
L149_163 V149 V163 8.413936734968221e-13
C149_163 V149 V163 5.709038258370411e-19

R149_164 V149 V164 -55.24591590531199
L149_164 V149 V164 9.881076132556763e-13
C149_164 V149 V164 1.500312794482553e-19

R149_165 V149 V165 -75.02937828469572
L149_165 V149 V165 -3.672563489760051e-13
C149_165 V149 V165 -1.6650720719384293e-18

R149_166 V149 V166 -32.09717080004667
L149_166 V149 V166 1.8566129471334235e-12
C149_166 V149 V166 3.198748181431519e-19

R149_167 V149 V167 -349.000998777727
L149_167 V149 V167 3.3420113254734496e-12
C149_167 V149 V167 1.4392976550500575e-19

R149_168 V149 V168 149.71516114011146
L149_168 V149 V168 2.7522225862979164e-12
C149_168 V149 V168 5.736539000476695e-19

R149_169 V149 V169 147.2323240484411
L149_169 V149 V169 -2.2785286684652857e-12
C149_169 V149 V169 -2.119757515530913e-21

R149_170 V149 V170 29.196535977679137
L149_170 V149 V170 -2.821282878654545e-12
C149_170 V149 V170 -8.392627331250262e-19

R149_171 V149 V171 58.554163099790166
L149_171 V149 V171 -3.873853464947473e-13
C149_171 V149 V171 -1.2285715585092512e-18

R149_172 V149 V172 68.88736082008698
L149_172 V149 V172 -7.10901292875797e-13
C149_172 V149 V172 -8.460199215173328e-19

R149_173 V149 V173 67.54399917887622
L149_173 V149 V173 8.290436668822684e-13
C149_173 V149 V173 5.4708413399489625e-19

R149_174 V149 V174 189.12207093156965
L149_174 V149 V174 -2.1384464358280883e-12
C149_174 V149 V174 6.504124185106924e-19

R149_175 V149 V175 -165.3970933447859
L149_175 V149 V175 -1.375191271434624e-12
C149_175 V149 V175 -3.67663181523429e-19

R149_176 V149 V176 -76.43005544958673
L149_176 V149 V176 -1.5160996325043228e-12
C149_176 V149 V176 -2.670711266713653e-19

R149_177 V149 V177 -74.46071802014353
L149_177 V149 V177 4.4009210915789225e-12
C149_177 V149 V177 -3.082124974198461e-19

R149_178 V149 V178 -49.49367818096507
L149_178 V149 V178 8.806581713005028e-13
C149_178 V149 V178 5.844348849758951e-19

R149_179 V149 V179 -304.5186894021264
L149_179 V149 V179 3.8374921842765387e-13
C149_179 V149 V179 1.475984621121148e-18

R149_180 V149 V180 -398.1591444267112
L149_180 V149 V180 3.831389202724035e-13
C149_180 V149 V180 1.1117108301262434e-18

R149_181 V149 V181 -128.63233368060745
L149_181 V149 V181 -1.8504037941950606e-12
C149_181 V149 V181 4.827149018677151e-19

R149_182 V149 V182 271.45341071746526
L149_182 V149 V182 -3.680388434273715e-13
C149_182 V149 V182 -9.528301072420844e-19

R149_183 V149 V183 311.9087803557577
L149_183 V149 V183 7.3780021808607e-13
C149_183 V149 V183 1.9632477817662796e-19

R149_184 V149 V184 103.87466596631911
L149_184 V149 V184 1.4693422160381865e-12
C149_184 V149 V184 -6.25864723394525e-21

R149_185 V149 V185 37.2051471068156
L149_185 V149 V185 1.4974652003434538e-12
C149_185 V149 V185 -1.1063748833032764e-19

R149_186 V149 V186 5523.744111090474
L149_186 V149 V186 4.522775572292895e-12
C149_186 V149 V186 1.7977034525473979e-19

R149_187 V149 V187 -929.3783211778448
L149_187 V149 V187 -4.31940595036872e-13
C149_187 V149 V187 -1.0133191316803048e-18

R149_188 V149 V188 -163.4368752496586
L149_188 V149 V188 -3.6596212892944905e-13
C149_188 V149 V188 -7.879480092356166e-19

R149_189 V149 V189 -89.34725312474399
L149_189 V149 V189 -9.222256872715852e-13
C149_189 V149 V189 -8.144304478977363e-19

R149_190 V149 V190 -118.6662901107449
L149_190 V149 V190 1.413146725220128e-12
C149_190 V149 V190 8.338878201907578e-19

R149_191 V149 V191 1080.9499134098535
L149_191 V149 V191 -4.475258056117343e-13
C149_191 V149 V191 -6.910863793151804e-19

R149_192 V149 V192 522.5958244364261
L149_192 V149 V192 -1.045181104734691e-12
C149_192 V149 V192 -6.448061182336234e-19

R149_193 V149 V193 -43.250319283342954
L149_193 V149 V193 1.2502596777828823e-11
C149_193 V149 V193 4.42815064554595e-19

R149_194 V149 V194 55.22533728928878
L149_194 V149 V194 -5.622077454539853e-12
C149_194 V149 V194 -7.408083535414228e-20

R149_195 V149 V195 143.53484974070082
L149_195 V149 V195 2.870332530884137e-13
C149_195 V149 V195 1.2835824736475537e-18

R149_196 V149 V196 153.89941618654626
L149_196 V149 V196 3.0632089194995206e-13
C149_196 V149 V196 1.4682379370418069e-18

R149_197 V149 V197 50.94702464083753
L149_197 V149 V197 6.258022977063429e-13
C149_197 V149 V197 6.895351933349166e-19

R149_198 V149 V198 -93.36965285959499
L149_198 V149 V198 -2.2071876898503084e-12
C149_198 V149 V198 -2.3516421897004857e-19

R149_199 V149 V199 -59.50517381785216
L149_199 V149 V199 8.955946720130158e-13
C149_199 V149 V199 5.042795269484458e-19

R149_200 V149 V200 -141.6711455577396
L149_200 V149 V200 2.0113612878209056e-12
C149_200 V149 V200 2.4260095252817136e-19

R150_150 V150 0 51.74888528389878
L150_150 V150 0 7.450505634032385e-13
C150_150 V150 0 3.621203371996849e-18

R150_151 V150 V151 985.1059368357969
L150_151 V150 V151 -1.8217777038794602e-11
C150_151 V150 V151 1.1723986232827924e-19

R150_152 V150 V152 48.54247700116889
L150_152 V150 V152 6.358711575706503e-12
C150_152 V150 V152 -7.632155320345115e-21

R150_153 V150 V153 -14.906793197524314
L150_153 V150 V153 -3.770057448067615e-12
C150_153 V150 V153 3.303117872047195e-19

R150_154 V150 V154 29.119713504696396
L150_154 V150 V154 3.955729820671054e-12
C150_154 V150 V154 9.325408319664849e-19

R150_155 V150 V155 78.62723262045553
L150_155 V150 V155 8.281689307687977e-12
C150_155 V150 V155 3.5451127222987995e-19

R150_156 V150 V156 -30.11290974656873
L150_156 V150 V156 -1.053119164189575e-11
C150_156 V150 V156 2.6189784553294e-19

R150_157 V150 V157 41059.561758328455
L150_157 V150 V157 -6.841900705127904e-12
C150_157 V150 V157 -1.6802646371056697e-18

R150_158 V150 V158 7.594187648475383
L150_158 V150 V158 9.674632227684035e-13
C150_158 V150 V158 -4.910111050682709e-20

R150_159 V150 V159 -24.663916510389473
L150_159 V150 V159 5.784871645822685e-11
C150_159 V150 V159 1.1191162685370467e-19

R150_160 V150 V160 -40.016277408896364
L150_160 V150 V160 2.2524473741619044e-11
C150_160 V150 V160 2.2042765489084883e-19

R150_161 V150 V161 17.28449719116041
L150_161 V150 V161 4.741977383761766e-12
C150_161 V150 V161 -2.6417473190851943e-19

R150_162 V150 V162 51.94773420795072
L150_162 V150 V162 -2.4723962278270463e-10
C150_162 V150 V162 5.674898724633944e-20

R150_163 V150 V163 31.711044283729223
L150_163 V150 V163 1.3060952835268364e-11
C150_163 V150 V163 -3.966515170471334e-19

R150_164 V150 V164 22.782992413404695
L150_164 V150 V164 5.77655317501382e-11
C150_164 V150 V164 -1.2718371135340944e-19

R150_165 V150 V165 -145.62208276078388
L150_165 V150 V165 -4.515539700468827e-12
C150_165 V150 V165 9.249485661104776e-19

R150_166 V150 V166 -4.814832768188761
L150_166 V150 V166 -7.360033581012968e-13
C150_166 V150 V166 -2.1051727069752274e-19

R150_167 V150 V167 23.697440672828527
L150_167 V150 V167 2.192914836147813e-11
C150_167 V150 V167 -1.816075998773259e-19

R150_168 V150 V168 16.80367353272214
L150_168 V150 V168 7.436527645735227e-12
C150_168 V150 V168 -3.8216698477789134e-19

R150_169 V150 V169 -15.5189863531597
L150_169 V150 V169 1.466507635145164e-11
C150_169 V150 V169 3.4914270644549994e-20

R150_170 V150 V170 10.158338002371309
L150_170 V150 V170 1.3362924811828346e-12
C150_170 V150 V170 4.2744525664163267e-19

R150_171 V150 V171 -28.176400650602282
L150_171 V150 V171 -1.1016302325879185e-11
C150_171 V150 V171 7.209393344300187e-19

R150_172 V150 V172 -21.360270692397343
L150_172 V150 V172 -3.7333037951962314e-12
C150_172 V150 V172 5.450869261973636e-19

R150_173 V150 V173 17.865400085584692
L150_173 V150 V173 3.93248625425113e-12
C150_173 V150 V173 -2.9451878552386824e-19

R150_174 V150 V174 7.441925876546776
L150_174 V150 V174 1.0788511926875708e-12
C150_174 V150 V174 -3.2610895617353253e-19

R150_175 V150 V175 -35.99882118921969
L150_175 V150 V175 9.41779698076084e-12
C150_175 V150 V175 1.3585115496838638e-19

R150_176 V150 V176 -29.834724280123776
L150_176 V150 V176 3.651788139621558e-12
C150_176 V150 V176 2.4088116973684647e-19

R150_177 V150 V177 43.587877043289815
L150_177 V150 V177 -6.093058949178701e-12
C150_177 V150 V177 6.380996895656586e-20

R150_178 V150 V178 -9.812688103864062
L150_178 V150 V178 -1.169618554472372e-12
C150_178 V150 V178 -2.940282823223732e-19

R150_179 V150 V179 30.522090078224355
L150_179 V150 V179 -5.721283929435261e-12
C150_179 V150 V179 -7.044956058687762e-19

R150_180 V150 V180 20.472243942575137
L150_180 V150 V180 -8.265590129241085e-12
C150_180 V150 V180 -6.420768576115504e-19

R150_181 V150 V181 -23.84734669753487
L150_181 V150 V181 -6.384328014844656e-12
C150_181 V150 V181 -2.8290576963547087e-19

R150_182 V150 V182 -14.014560041358404
L150_182 V150 V182 -7.538121543322465e-12
C150_182 V150 V182 4.857196975869781e-19

R150_183 V150 V183 259.0990303552616
L150_183 V150 V183 -6.9529307956641216e-12
C150_183 V150 V183 -1.0328070749864907e-19

R150_184 V150 V184 688.3882258572181
L150_184 V150 V184 -2.6631876398035812e-12
C150_184 V150 V184 7.148034424601948e-20

R150_185 V150 V185 718.4761929217924
L150_185 V150 V185 3.810476140723174e-11
C150_185 V150 V185 1.3219785433136141e-19

R150_186 V150 V186 32.22125639675747
L150_186 V150 V186 4.977416130591179e-12
C150_186 V150 V186 -1.0034610803320073e-19

R150_187 V150 V187 -220.80491545438514
L150_187 V150 V187 1.824369991584886e-11
C150_187 V150 V187 4.720489559396347e-19

R150_188 V150 V188 -117.08752559249588
L150_188 V150 V188 2.2311785485436554e-12
C150_188 V150 V188 3.3173757942661935e-19

R150_189 V150 V189 80.77707326314463
L150_189 V150 V189 8.484002706878448e-12
C150_189 V150 V189 5.34208981509135e-19

R150_190 V150 V190 59.037289351900924
L150_190 V150 V190 -5.356996473029309e-11
C150_190 V150 V190 -5.5703135535153665e-19

R150_191 V150 V191 -115.74504423293604
L150_191 V150 V191 4.077735381842489e-11
C150_191 V150 V191 4.0712768127224995e-19

R150_192 V150 V192 -825.0264787129998
L150_192 V150 V192 -4.9811890329494124e-12
C150_192 V150 V192 3.4830169254845957e-19

R150_193 V150 V193 4741.7802621346855
L150_193 V150 V193 -6.267774078790259e-12
C150_193 V150 V193 -2.7224079333660926e-19

R150_194 V150 V194 -283.26719291455834
L150_194 V150 V194 3.1357980921186386e-12
C150_194 V150 V194 8.782354265912068e-20

R150_195 V150 V195 791.3023205261583
L150_195 V150 V195 -7.294134167997597e-12
C150_195 V150 V195 -8.605762968637012e-19

R150_196 V150 V196 -643.0926189300098
L150_196 V150 V196 5.895582856458061e-12
C150_196 V150 V196 -6.704974484559938e-19

R150_197 V150 V197 238.964423370934
L150_197 V150 V197 3.625077243141748e-11
C150_197 V150 V197 -4.880612788446263e-19

R150_198 V150 V198 -20.364786316231378
L150_198 V150 V198 -4.267192320975003e-12
C150_198 V150 V198 3.3649307951765596e-20

R150_199 V150 V199 -235.866040930466
L150_199 V150 V199 5.156523716658138e-10
C150_199 V150 V199 -3.858639930541881e-19

R150_200 V150 V200 38.83659347833558
L150_200 V150 V200 -1.2292823342470091e-11
C150_200 V150 V200 -1.4355740006478623e-19

R151_151 V151 0 88.08316302740114
L151_151 V151 0 1.4397283529046878e-12
C151_151 V151 0 -5.291838574019413e-19

R151_152 V151 V152 -63.87648555374038
L151_152 V151 V152 -1.0505466598065365e-11
C151_152 V151 V152 3.8118613179375e-20

R151_153 V151 V153 -42.73799484644736
L151_153 V151 V153 -1.3567870027201745e-11
C151_153 V151 V153 1.3845290315195829e-19

R151_154 V151 V154 -35.20666701426782
L151_154 V151 V154 -3.3081742690871507e-12
C151_154 V151 V154 -9.244605722743144e-20

R151_155 V151 V155 9.795788486139928
L151_155 V151 V155 -6.066221703716556e-12
C151_155 V151 V155 5.711408693477938e-21

R151_156 V151 V156 -408.6608140762014
L151_156 V151 V156 -7.90722321061569e-12
C151_156 V151 V156 2.2042858529045704e-20

R151_157 V151 V157 -167.58573884024764
L151_157 V151 V157 1.945820951926188e-12
C151_157 V151 V157 4.529206541700214e-19

R151_158 V151 V158 -81.9638047754775
L151_158 V151 V158 -7.940698303555752e-12
C151_158 V151 V158 -6.979003462041279e-20

R151_159 V151 V159 14.704329187588968
L151_159 V151 V159 5.057622147197411e-13
C151_159 V151 V159 2.2268982432974623e-19

R151_160 V151 V160 -606.3788782260625
L151_160 V151 V160 -5.953706647506318e-11
C151_160 V151 V160 -6.382979294596382e-20

R151_161 V151 V161 609.2528669474241
L151_161 V151 V161 -5.282557911948409e-12
C151_161 V151 V161 -1.524983144982088e-19

R151_162 V151 V162 193.60352409419173
L151_162 V151 V162 -1.6191544641796694e-11
C151_162 V151 V162 -9.777056158139036e-20

R151_163 V151 V163 -19.63040899192734
L151_163 V151 V163 -2.9752830670733842e-12
C151_163 V151 V163 -1.530361138270317e-21

R151_164 V151 V164 -112.76253218646171
L151_164 V151 V164 4.7872834463477675e-12
C151_164 V151 V164 -1.1931897791908507e-20

R151_165 V151 V165 116.28295692037881
L151_165 V151 V165 -1.5778039973043671e-12
C151_165 V151 V165 -2.232351118915902e-19

R151_166 V151 V166 37.239585510877056
L151_166 V151 V166 -4.4449217171248184e-11
C151_166 V151 V166 2.3567471898603325e-20

R151_167 V151 V167 -13.498722510170241
L151_167 V151 V167 -8.513820741947876e-13
C151_167 V151 V167 -1.814802817362535e-19

R151_168 V151 V168 81.27348551735429
L151_168 V151 V168 -5.575473774276552e-12
C151_168 V151 V168 5.517519297073965e-21

R151_169 V151 V169 238.0134305561701
L151_169 V151 V169 1.796501715380339e-12
C151_169 V151 V169 2.118492706643466e-19

R151_170 V151 V170 -89.67006242313421
L151_170 V151 V170 7.190072383419883e-10
C151_170 V151 V170 -9.478083156176383e-20

R151_171 V151 V171 11.80491793040454
L151_171 V151 V171 3.119715508700227e-12
C151_171 V151 V171 3.743805301753699e-20

R151_172 V151 V172 100.45007760845863
L151_172 V151 V172 -3.543072047817174e-10
C151_172 V151 V172 -2.784960132909481e-20

R151_173 V151 V173 -86.67060967909627
L151_173 V151 V173 7.254556234939995e-12
C151_173 V151 V173 1.1462189279839218e-20

R151_174 V151 V174 -40.071747930918264
L151_174 V151 V174 6.042880815963349e-12
C151_174 V151 V174 1.5974849831729711e-19

R151_175 V151 V175 351.038503213541
L151_175 V151 V175 2.5391108022182324e-12
C151_175 V151 V175 -2.8345939956266756e-19

R151_176 V151 V176 -675.3400953388239
L151_176 V151 V176 3.5329691540622702e-12
C151_176 V151 V176 1.2257893755798277e-19

R151_177 V151 V177 -105.57201176458636
L151_177 V151 V177 -4.4306638695026544e-12
C151_177 V151 V177 -7.67865733920671e-20

R151_178 V151 V178 80.38267218919344
L151_178 V151 V178 6.755335100785056e-12
C151_178 V151 V178 8.692595934754505e-20

R151_179 V151 V179 -44.092623622842716
L151_179 V151 V179 -1.2444315217584678e-11
C151_179 V151 V179 4.74299457522988e-19

R151_180 V151 V180 -85.44044122577036
L151_180 V151 V180 7.805309329394845e-12
C151_180 V151 V180 6.389051458276462e-20

R151_181 V151 V181 88.2963893398501
L151_181 V151 V181 6.30982614302278e-11
C151_181 V151 V181 -6.801740019887329e-20

R151_182 V151 V182 47.23689415176286
L151_182 V151 V182 -2.3364820699135167e-12
C151_182 V151 V182 -2.1026113355320338e-19

R151_183 V151 V183 -223.48190755846989
L151_183 V151 V183 5.0904931262506396e-12
C151_183 V151 V183 -1.3222428378848592e-20

R151_184 V151 V184 231.714299205516
L151_184 V151 V184 1.4215960759855143e-11
C151_184 V151 V184 7.333839548420295e-20

R151_185 V151 V185 827.1487443149633
L151_185 V151 V185 -4.180890792899736e-12
C151_185 V151 V185 5.760692392998583e-20

R151_186 V151 V186 -358.99408008928134
L151_186 V151 V186 -4.145820616281042e-12
C151_186 V151 V186 2.5823829967730093e-20

R151_187 V151 V187 515.3355536207686
L151_187 V151 V187 -1.9990897940914493e-12
C151_187 V151 V187 -3.735023984952559e-19

R151_188 V151 V188 141.25562076661342
L151_188 V151 V188 -1.2095376529098315e-12
C151_188 V151 V188 -1.6940750430885296e-19

R151_189 V151 V189 -139.38558576425763
L151_189 V151 V189 2.495753062179178e-12
C151_189 V151 V189 1.531845371448228e-20

R151_190 V151 V190 -82.74644035484292
L151_190 V151 V190 4.750385315147148e-12
C151_190 V151 V190 1.1102751406425772e-19

R151_191 V151 V191 -6088.490873520562
L151_191 V151 V191 -5.38605239289056e-12
C151_191 V151 V191 8.274177041363508e-20

R151_192 V151 V192 -116.8409527227311
L151_192 V151 V192 3.57470158764596e-12
C151_192 V151 V192 -7.253933773606414e-20

R151_193 V151 V193 -392.8016242168312
L151_193 V151 V193 4.806964052591434e-12
C151_193 V151 V193 5.239065807715597e-20

R151_194 V151 V194 807.7667635540487
L151_194 V151 V194 2.2745192291633045e-12
C151_194 V151 V194 1.356638849221114e-19

R151_195 V151 V195 83.45429929930579
L151_195 V151 V195 1.867211359718156e-12
C151_195 V151 V195 -1.27840442460478e-19

R151_196 V151 V196 -106.75236851859536
L151_196 V151 V196 1.6273964316171035e-12
C151_196 V151 V196 3.5308284330525137e-19

R151_197 V151 V197 -837.2872236864561
L151_197 V151 V197 -5.424062869979923e-12
C151_197 V151 V197 -5.287580629146619e-20

R151_198 V151 V198 133.81085483334985
L151_198 V151 V198 -6.221998976204574e-12
C151_198 V151 V198 -7.530081460456159e-20

R151_199 V151 V199 -192.24581705228474
L151_199 V151 V199 -2.3688884964275023e-11
C151_199 V151 V199 7.942233093281407e-20

R151_200 V151 V200 668.7483013263509
L151_200 V151 V200 -2.9113671737571756e-12
C151_200 V151 V200 -1.0521531079301887e-19

R152_152 V152 0 906.4952598910014
L152_152 V152 0 -3.152346696371677e-13
C152_152 V152 0 -5.043698269095232e-19

R152_153 V152 V153 -123.38685129166714
L152_153 V152 V153 -1.688056690614177e-12
C152_153 V152 V153 -6.637451428135086e-20

R152_154 V152 V154 -35.33297078005107
L152_154 V152 V154 -1.8032326340548567e-12
C152_154 V152 V154 6.98899427211526e-20

R152_155 V152 V155 237.4513224175347
L152_155 V152 V155 -1.5649993958296567e-09
C152_155 V152 V155 1.456711708226797e-19

R152_156 V152 V156 25.143069415860026
L152_156 V152 V156 3.3579901467354384e-12
C152_156 V152 V156 -2.707599692765951e-19

R152_157 V152 V157 444.6799479953638
L152_157 V152 V157 1.4022051096892717e-12
C152_157 V152 V157 -1.1448856646020317e-20

R152_158 V152 V158 -44.01342802838587
L152_158 V152 V158 1.5991128066969427e-11
C152_158 V152 V158 -4.361301227913442e-20

R152_159 V152 V159 217.17800162218154
L152_159 V152 V159 -1.8845103150039413e-12
C152_159 V152 V159 -1.7929886710987365e-19

R152_160 V152 V160 12.6788188773185
L152_160 V152 V160 5.700489311256213e-13
C152_160 V152 V160 2.5271020094439843e-19

R152_161 V152 V161 -77.52286689699727
L152_161 V152 V161 -1.9861658888847975e-12
C152_161 V152 V161 -3.8462409238783055e-20

R152_162 V152 V162 278.62789005633533
L152_162 V152 V162 -6.79537485786445e-12
C152_162 V152 V162 -3.3926810551815286e-20

R152_163 V152 V163 -64.57162571276166
L152_163 V152 V163 5.876058134425888e-12
C152_163 V152 V163 4.062574689480496e-20

R152_164 V152 V164 -16.399704056872004
L152_164 V152 V164 -1.1093752580819778e-12
C152_164 V152 V164 -1.4251657677237136e-19

R152_165 V152 V165 181.2397949337833
L152_165 V152 V165 3.4604403011749736e-12
C152_165 V152 V165 1.4567102499909862e-19

R152_166 V152 V166 25.848769617830154
L152_166 V152 V166 3.0680335951316162e-12
C152_166 V152 V166 1.0842736075380848e-19

R152_167 V152 V167 -314.4574208693288
L152_167 V152 V167 7.249881003384167e-12
C152_167 V152 V167 -3.6892797116309295e-20

R152_168 V152 V168 -22.971485490261447
L152_168 V152 V168 -9.111042857166877e-13
C152_168 V152 V168 4.361743899569356e-20

R152_169 V152 V169 56.068714925913966
L152_169 V152 V169 4.405219640352284e-12
C152_169 V152 V169 7.964070867820778e-21

R152_170 V152 V170 -51.789647261739276
L152_170 V152 V170 -5.01593017811675e-12
C152_170 V152 V170 1.4507870693503302e-20

R152_171 V152 V171 68.26353718980405
L152_171 V152 V171 -2.2727881598887554e-12
C152_171 V152 V171 8.138185903503141e-20

R152_172 V152 V172 16.828777306437328
L152_172 V152 V172 6.623764251164698e-13
C152_172 V152 V172 8.207280331178773e-20

R152_173 V152 V173 -61.06370024833889
L152_173 V152 V173 -2.6134385574279674e-12
C152_173 V152 V173 -9.782523005204e-20

R152_174 V152 V174 -32.086339330090844
L152_174 V152 V174 -2.9674630300749536e-11
C152_174 V152 V174 -7.115378292576511e-20

R152_175 V152 V175 955.0611603727247
L152_175 V152 V175 2.013930377643004e-12
C152_175 V152 V175 5.506549728910717e-20

R152_176 V152 V176 301.4939405191294
L152_176 V152 V176 -1.0902088298679868e-12
C152_176 V152 V176 -3.2741595766976035e-19

R152_177 V152 V177 -104.27006906733206
L152_177 V152 V177 6.8163593366164744e-12
C152_177 V152 V177 8.574442045892157e-20

R152_178 V152 V178 43.85633147107106
L152_178 V152 V178 4.232431613350953e-12
C152_178 V152 V178 -9.400524279094714e-21

R152_179 V152 V179 -2611.1012325345787
L152_179 V152 V179 4.264032681095099e-12
C152_179 V152 V179 -7.048845254284534e-20

R152_180 V152 V180 -28.670496211160486
L152_180 V152 V180 1.3121124028501561e-11
C152_180 V152 V180 1.9075984847923243e-19

R152_181 V152 V181 67.88924057254769
L152_181 V152 V181 1.150428377782306e-11
C152_181 V152 V181 3.0450007888957344e-20

R152_182 V152 V182 46.224427251821076
L152_182 V152 V182 1.3957818132475941e-11
C152_182 V152 V182 6.912667397958237e-20

R152_183 V152 V183 -1808.6403612274717
L152_183 V152 V183 1.3307595269517435e-11
C152_183 V152 V183 4.258776927329554e-20

R152_184 V152 V184 48.22143260386261
L152_184 V152 V184 1.4926129734058795e-12
C152_184 V152 V184 -5.1389117166544006e-20

R152_185 V152 V185 344.1016334658809
L152_185 V152 V185 -7.197930824493492e-12
C152_185 V152 V185 -8.420714502918738e-20

R152_186 V152 V186 7367.524717940558
L152_186 V152 V186 3.736430049751223e-12
C152_186 V152 V186 -1.986388912043144e-20

R152_187 V152 V187 361.5802866189602
L152_187 V152 V187 3.573300125664618e-12
C152_187 V152 V187 2.784569095103582e-20

R152_188 V152 V188 -61.685683224945734
L152_188 V152 V188 -5.568199439034831e-13
C152_188 V152 V188 -2.603689679044139e-21

R152_189 V152 V189 -154.57530145519067
L152_189 V152 V189 4.477831167293059e-12
C152_189 V152 V189 6.553245194696257e-20

R152_190 V152 V190 -79.69780641896185
L152_190 V152 V190 -7.578071862553952e-12
C152_190 V152 V190 -2.6982039624625824e-20

R152_191 V152 V191 -133.9808269708966
L152_191 V152 V191 -1.2038462683002535e-12
C152_191 V152 V191 -6.47800779768081e-20

R152_192 V152 V192 795.0965201039487
L152_192 V152 V192 9.419942269977132e-13
C152_192 V152 V192 1.7019931547260497e-19

R152_193 V152 V193 -219.865010284291
L152_193 V152 V193 -2.3751690681236958e-11
C152_193 V152 V193 -1.1004622431797351e-20

R152_194 V152 V194 325.32850014305535
L152_194 V152 V194 2.621250920956162e-12
C152_194 V152 V194 8.128232691703277e-20

R152_195 V152 V195 239.2741549429659
L152_195 V152 V195 9.418849137467722e-13
C152_195 V152 V195 2.2194299699005254e-19

R152_196 V152 V196 77.41313994668583
L152_196 V152 V196 -1.0199374746471913e-12
C152_196 V152 V196 -5.142637476956102e-19

R152_197 V152 V197 223.36588322019352
L152_197 V152 V197 -1.7239050090071972e-11
C152_197 V152 V197 -4.8209742324677054e-20

R152_198 V152 V198 134.3978535673356
L152_198 V152 V198 7.699715809308485e-12
C152_198 V152 V198 6.183362134966638e-20

R152_199 V152 V199 -226.05147302361223
L152_199 V152 V199 -1.1672347889500939e-11
C152_199 V152 V199 -9.393498169314673e-20

R152_200 V152 V200 -114.52819600724584
L152_200 V152 V200 2.0061565397149864e-11
C152_200 V152 V200 1.3533024069426377e-19

R153_153 V153 0 44.74550811829922
L153_153 V153 0 -2.1276258532569742e-13
C153_153 V153 0 -1.0528782807684972e-18

R153_154 V153 V154 -100.77335680032947
L153_154 V153 V154 -1.6800543546891936e-12
C153_154 V153 V154 -2.860044420533165e-19

R153_155 V153 V155 79.32667497656617
L153_155 V153 V155 -5.8291569605477754e-12
C153_155 V153 V155 3.466996075736492e-20

R153_156 V153 V156 -61.21490204759935
L153_156 V153 V156 -2.4616472554756082e-12
C153_156 V153 V156 -1.2646460344069105e-19

R153_157 V153 V157 -64.49587472779977
L153_157 V153 V157 6.6935676050099635e-12
C153_157 V153 V157 2.851286641780976e-19

R153_158 V153 V158 20.428753051976255
L153_158 V153 V158 2.2203586417586405e-12
C153_158 V153 V158 5.8877980387542574e-21

R153_159 V153 V159 1136.324307037882
L153_159 V153 V159 -5.483552195252552e-12
C153_159 V153 V159 -3.022912742845215e-19

R153_160 V153 V160 49.04931917198333
L153_160 V153 V160 2.3451884193277692e-12
C153_160 V153 V160 -6.417494837569117e-20

R153_161 V153 V161 32.95373377085268
L153_161 V153 V161 8.30954479822432e-13
C153_161 V153 V161 5.748823540933518e-19

R153_162 V153 V162 56.384942950615155
L153_162 V153 V162 9.009831200053892e-12
C153_162 V153 V162 -6.663625062224255e-20

R153_163 V153 V163 90.08901366317761
L153_163 V153 V163 2.3982814698001248e-11
C153_163 V153 V163 4.667271794819637e-20

R153_164 V153 V164 67.24258498399298
L153_164 V153 V164 4.1183006273336234e-12
C153_164 V153 V164 5.848531592698878e-20

R153_165 V153 V165 105.4077560790617
L153_165 V153 V165 1.6199228749526712e-12
C153_165 V153 V165 -8.161994748332714e-20

R153_166 V153 V166 -14.868315882927915
L153_166 V153 V166 2.6000632725387738e-11
C153_166 V153 V166 2.5227445412605508e-19

R153_167 V153 V167 -368.7094740347796
L153_167 V153 V167 3.900496258091677e-12
C153_167 V153 V167 2.261836900934041e-19

R153_168 V153 V168 -2356.26989343481
L153_168 V153 V168 -7.1878152304058156e-12
C153_168 V153 V168 3.4875950922058437e-19

R153_169 V153 V169 -30.433385246017718
L153_169 V153 V169 -1.0538733234425634e-12
C153_169 V153 V169 -5.070319130923832e-19

R153_170 V153 V170 40.476850628844595
L153_170 V153 V170 7.610633039452355e-12
C153_170 V153 V170 -7.170593004778079e-20

R153_171 V153 V171 -409.69895497117216
L153_171 V153 V171 -2.3766763719210465e-10
C153_171 V153 V171 -7.616242211533734e-20

R153_172 V153 V172 -211.90227348052835
L153_172 V153 V172 6.270963515518851e-12
C153_172 V153 V172 -2.0919375674388125e-19

R153_173 V153 V173 109.35552542653457
L153_173 V153 V173 -6.827375657296849e-12
C153_173 V153 V173 -1.56832362442163e-20

R153_174 V153 V174 22.852233055930036
L153_174 V153 V174 -1.4602270840246435e-12
C153_174 V153 V174 -3.5151282189694444e-19

R153_175 V153 V175 -216.307493780734
L153_175 V153 V175 -2.4353038661184933e-12
C153_175 V153 V175 -1.583873540330472e-19

R153_176 V153 V176 -836.9110531028356
L153_176 V153 V176 -1.1820371148119351e-12
C153_176 V153 V176 -3.355501256819717e-19

R153_177 V153 V177 66.26251155201652
L153_177 V153 V177 4.200347370205537e-12
C153_177 V153 V177 2.201547388799208e-19

R153_178 V153 V178 -34.31883131750662
L153_178 V153 V178 7.737802187315547e-12
C153_178 V153 V178 1.4488696392448043e-19

R153_179 V153 V179 155.89134767250067
L153_179 V153 V179 5.761614549415412e-12
C153_179 V153 V179 5.1572366541317065e-20

R153_180 V153 V180 304.7404545870699
L153_180 V153 V180 2.4336309860796955e-12
C153_180 V153 V180 2.3723118562723927e-19

R153_181 V153 V181 -119.01959961797418
L153_181 V153 V181 5.391505500388926e-12
C153_181 V153 V181 3.338325606450203e-19

R153_182 V153 V182 -48.40774170363486
L153_182 V153 V182 5.455986823245497e-12
C153_182 V153 V182 1.1292455854284143e-20

R153_183 V153 V183 639.4173635501446
L153_183 V153 V183 1.458036867670416e-11
C153_183 V153 V183 -1.874316628658308e-20

R153_184 V153 V184 240.2719699899237
L153_184 V153 V184 2.864271169110141e-12
C153_184 V153 V184 -1.334352912967687e-20

R153_185 V153 V185 -60.98456239882801
L153_185 V153 V185 3.5671841661146687e-12
C153_185 V153 V185 -2.8581061583803147e-19

R153_186 V153 V186 61.38387294280944
L153_186 V153 V186 2.462953525071775e-12
C153_186 V153 V186 1.2954739096522974e-19

R153_187 V153 V187 857.2086764556811
L153_187 V153 V187 2.5494647770441796e-12
C153_187 V153 V187 1.2602828137634385e-19

R153_188 V153 V188 -346.2954885818081
L153_188 V153 V188 -1.0813976505692908e-11
C153_188 V153 V188 1.8024609669793456e-19

R153_189 V153 V189 105.13002347821538
L153_189 V153 V189 -1.5113035494397227e-12
C153_189 V153 V189 -1.5122354214362583e-19

R153_190 V153 V190 265.0294851955056
L153_190 V153 V190 -5.413447535513374e-12
C153_190 V153 V190 9.135068535881385e-20

R153_191 V153 V191 -87.050237153427
L153_191 V153 V191 -2.7903832849505804e-12
C153_191 V153 V191 -8.084659905795659e-20

R153_192 V153 V192 -185.61859494699792
L153_192 V153 V192 -4.295741628072753e-12
C153_192 V153 V192 -2.4749811628399323e-19

R153_193 V153 V193 70.46745538177761
L153_193 V153 V193 8.333083440490174e-12
C153_193 V153 V193 -7.731455158765682e-20

R153_194 V153 V194 -86.1986064142041
L153_194 V153 V194 -1.343062729942708e-12
C153_194 V153 V194 -4.0804226915759195e-19

R153_195 V153 V195 258.5272793683332
L153_195 V153 V195 3.64218967166077e-12
C153_195 V153 V195 1.5774664815369951e-19

R153_196 V153 V196 -1547.3588199694127
L153_196 V153 V196 -1.756161576669857e-12
C153_196 V153 V196 -9.397242881859616e-20

R153_197 V153 V197 -107.13849382917645
L153_197 V153 V197 4.21328583057169e-12
C153_197 V153 V197 3.248864808893406e-19

R153_198 V153 V198 -97.62358694949704
L153_198 V153 V198 3.56481435515784e-12
C153_198 V153 V198 4.1087458732924566e-20

R153_199 V153 V199 185.59501466843477
L153_199 V153 V199 9.358817313924264e-12
C153_199 V153 V199 -5.690467652742638e-20

R153_200 V153 V200 67.68566740583798
L153_200 V153 V200 1.6384132421667633e-12
C153_200 V153 V200 2.605890696978047e-19

R154_154 V154 0 -65.2060964068682
L154_154 V154 0 -4.3265203307500387e-13
C154_154 V154 0 -2.3755944285144693e-18

R154_155 V154 V155 248.87577843051787
L154_155 V154 V155 -1.2019872646593134e-11
C154_155 V154 V155 -1.3209381359925614e-19

R154_156 V154 V156 147.61620758137468
L154_156 V154 V156 -4.574210909482624e-12
C154_156 V154 V156 -1.0851626319691278e-19

R154_157 V154 V157 -43.691370213504165
L154_157 V154 V157 4.4679059504007696e-12
C154_157 V154 V157 1.3799933581742064e-18

R154_158 V154 V158 180.76051684946233
L154_158 V154 V158 8.509495859102941e-12
C154_158 V154 V158 1.0771841928078116e-19

R154_159 V154 V159 33.562753646384664
L154_159 V154 V159 2.3878923305980727e-11
C154_159 V154 V159 -2.2638991149126265e-19

R154_160 V154 V160 31.223791337577573
L154_160 V154 V160 2.6624513332172908e-12
C154_160 V154 V160 -2.550493424612193e-19

R154_161 V154 V161 -212.86415900628137
L154_161 V154 V161 3.04852106256618e-12
C154_161 V154 V161 3.295216702269253e-19

R154_162 V154 V162 24.59600738804507
L154_162 V154 V162 1.5997503498136442e-12
C154_162 V154 V162 1.450541621343661e-20

R154_163 V154 V163 -63.1379481350201
L154_163 V154 V163 5.944714130874028e-12
C154_163 V154 V163 4.353663102070334e-19

R154_164 V154 V164 -43.50042282078282
L154_164 V154 V164 1.3563696686778483e-11
C154_164 V154 V164 2.0667854718680623e-19

R154_165 V154 V165 35.05864359570639
L154_165 V154 V165 6.129685937985457e-12
C154_165 V154 V165 -9.67925523465423e-19

R154_166 V154 V166 -342.0304289913747
L154_166 V154 V166 -1.1454471501856188e-11
C154_166 V154 V166 1.037822716818832e-19

R154_167 V154 V167 -127.05726397899419
L154_167 V154 V167 1.490353236402941e-11
C154_167 V154 V167 1.3407199292008755e-19

R154_168 V154 V168 -770.1100108538619
L154_168 V154 V168 1.6011030215710562e-11
C154_168 V154 V168 3.5150883578216983e-19

R154_169 V154 V169 96.38376016623471
L154_169 V154 V169 -2.3712185353566652e-12
C154_169 V154 V169 -1.3329542480243758e-19

R154_170 V154 V170 -35.52604815762113
L154_170 V154 V170 -2.5703224772611658e-12
C154_170 V154 V170 -3.977144248042272e-19

R154_171 V154 V171 69.94158298496212
L154_171 V154 V171 -2.6195704520147096e-12
C154_171 V154 V171 -6.952638728322471e-19

R154_172 V154 V172 92.89529670362393
L154_172 V154 V172 -7.229900369662788e-12
C154_172 V154 V172 -5.391000121315777e-19

R154_173 V154 V173 -30.194907348392537
L154_173 V154 V173 -1.2414012084576393e-11
C154_173 V154 V173 4.2439249822814063e-19

R154_174 V154 V174 50.30532425269133
L154_174 V154 V174 -7.105137689471193e-12
C154_174 V154 V174 2.6848779575777538e-19

R154_175 V154 V175 19356.257380200685
L154_175 V154 V175 -1.1395684903986766e-11
C154_175 V154 V175 -1.634999904047645e-20

R154_176 V154 V176 -136.17298760989323
L154_176 V154 V176 -2.3178081210183006e-12
C154_176 V154 V176 -4.9541564253054775e-20

R154_177 V154 V177 -3188.6969103762763
L154_177 V154 V177 3.5762913899503116e-12
C154_177 V154 V177 -1.0590306588107977e-19

R154_178 V154 V178 79.51314951573787
L154_178 V154 V178 1.820674581474577e-12
C154_178 V154 V178 2.80340237130817e-19

R154_179 V154 V179 -212.19051742631694
L154_179 V154 V179 2.7455327224654248e-12
C154_179 V154 V179 5.703558251551773e-19

R154_180 V154 V180 -1499.6026509219596
L154_180 V154 V180 1.8104156654957994e-12
C154_180 V154 V180 4.5386670637812655e-19

R154_181 V154 V181 56.91444303661228
L154_181 V154 V181 3.831186878449173e-11
C154_181 V154 V181 1.9979348400493944e-19

R154_182 V154 V182 -725.3883532319588
L154_182 V154 V182 -2.076895655018962e-12
C154_182 V154 V182 -4.3084906146727157e-19

R154_183 V154 V183 -420.95468218338596
L154_183 V154 V183 1.1414977580573963e-10
C154_183 V154 V183 6.13791187037405e-20

R154_184 V154 V184 -5207.518740977615
L154_184 V154 V184 7.630633708871402e-12
C154_184 V154 V184 -4.451021432125795e-20

R154_185 V154 V185 -95.97980750476978
L154_185 V154 V185 -6.890350330183227e-12
C154_185 V154 V185 -8.537918077806234e-20

R154_186 V154 V186 255.02540547600694
L154_186 V154 V186 -6.283437293340493e-11
C154_186 V154 V186 6.317001169954425e-20

R154_187 V154 V187 240.06699538952913
L154_187 V154 V187 -4.1872827342755267e-11
C154_187 V154 V187 -3.1219503742972e-19

R154_188 V154 V188 -138.95516765606152
L154_188 V154 V188 -1.4481154768756154e-12
C154_188 V154 V188 -2.337384346985697e-19

R154_189 V154 V189 -4577.923711196527
L154_189 V154 V189 -9.272657992935335e-12
C154_189 V154 V189 -4.957261552158989e-19

R154_190 V154 V190 65.54507022158424
L154_190 V154 V190 2.3188014031868056e-12
C154_190 V154 V190 4.621881472045445e-19

R154_191 V154 V191 272.82429667903995
L154_191 V154 V191 -3.795539695115546e-12
C154_191 V154 V191 -4.537891023229455e-19

R154_192 V154 V192 263.4912640720384
L154_192 V154 V192 7.331064901764888e-12
C154_192 V154 V192 -4.447962292625677e-19

R154_193 V154 V193 183.05753875563101
L154_193 V154 V193 8.565984137134984e-12
C154_193 V154 V193 2.3743413246863623e-19

R154_194 V154 V194 -127.09841893099342
L154_194 V154 V194 -2.2769682363106705e-12
C154_194 V154 V194 -2.1444997329603978e-19

R154_195 V154 V195 -326.502626964822
L154_195 V154 V195 2.541178370507358e-12
C154_195 V154 V195 7.967574962024506e-19

R154_196 V154 V196 9911.792462550888
L154_196 V154 V196 -2.1527074943817066e-11
C154_196 V154 V196 8.0211032900881815e-19

R154_197 V154 V197 -80.87673397214284
L154_197 V154 V197 9.396007542634506e-12
C154_197 V154 V197 4.88652730878358e-19

R154_198 V154 V198 -234.2694944758329
L154_198 V154 V198 -4.949516264887711e-12
C154_198 V154 V198 -6.514935849724978e-20

R154_199 V154 V199 -297.5441106406643
L154_199 V154 V199 2.685134738159083e-11
C154_199 V154 V199 3.5869524073813773e-19

R154_200 V154 V200 -78.48048508248336
L154_200 V154 V200 1.0294513833054395e-11
C154_200 V154 V200 1.819928135240757e-19

R155_155 V155 0 -37.27081217243093
L155_155 V155 0 -3.26252155434439e-13
C155_155 V155 0 -9.518347885637537e-19

R155_156 V155 V156 108.65422077771504
L155_156 V155 V156 -1.0286873622152855e-11
C155_156 V155 V156 2.821073119297329e-20

R155_157 V155 V157 -154.838241719188
L155_157 V155 V157 7.059035646562744e-13
C155_157 V155 V157 5.475678695641602e-19

R155_158 V155 V158 90.34185600343069
L155_158 V155 V158 -1.3313430723515045e-11
C155_158 V155 V158 -8.474845493590217e-20

R155_159 V155 V159 -48.65845816385856
L155_159 V155 V159 9.375063666525804e-13
C155_159 V155 V159 7.476019093933608e-19

R155_160 V155 V160 68.03453761933467
L155_160 V155 V160 4.448559654560993e-11
C155_160 V155 V160 -1.8485636924044116e-19

R155_161 V155 V161 338.6003847645713
L155_161 V155 V161 -1.555953519749845e-11
C155_161 V155 V161 -9.678823059085629e-20

R155_162 V155 V162 223.82466282040915
L155_162 V155 V162 -1.832556157266225e-12
C155_162 V155 V162 -8.889463851291882e-20

R155_163 V155 V163 14.285646785652766
L155_163 V155 V163 1.0380964473754607e-12
C155_163 V155 V163 -3.2223462771169824e-19

R155_164 V155 V164 173.6944675520147
L155_164 V155 V164 3.523444290642267e-12
C155_164 V155 V164 1.5387911083934834e-20

R155_165 V155 V165 138.23627312336856
L155_165 V155 V165 -8.520781797609714e-12
C155_165 V155 V165 -2.0193671447492581e-19

R155_166 V155 V166 -71.25848286751962
L155_166 V155 V166 3.2662161415815507e-12
C155_166 V155 V166 1.0872770298134713e-19

R155_167 V155 V167 33.98498329651739
L155_167 V155 V167 -1.5702210367011874e-12
C155_167 V155 V167 2.168659064593623e-19

R155_168 V155 V168 -54.7919253480848
L155_168 V155 V168 -5.603305356243679e-12
C155_168 V155 V168 -3.669844256202844e-20

R155_169 V155 V169 1109.6792717866313
L155_169 V155 V169 9.802841988573767e-12
C155_169 V155 V169 2.2616501092280117e-19

R155_170 V155 V170 112.5016303964283
L155_170 V155 V170 7.312875338132943e-11
C155_170 V155 V170 -1.8705702272676902e-19

R155_171 V155 V171 -11.746491461760353
L155_171 V155 V171 -2.5788112764622844e-12
C155_171 V155 V171 -2.1471068791872973e-19

R155_172 V155 V172 -221.63975391848746
L155_172 V155 V172 -7.140347195121264e-12
C155_172 V155 V172 -5.0312881429029906e-20

R155_173 V155 V173 -228.11558272453615
L155_173 V155 V173 -3.46772106764568e-12
C155_173 V155 V173 -5.325560230733974e-20

R155_174 V155 V174 142.77706402940774
L155_174 V155 V174 -3.0922391390844326e-12
C155_174 V155 V174 2.130336758142675e-19

R155_175 V155 V175 29.632838265741363
L155_175 V155 V175 -1.572984458157255e-12
C155_175 V155 V175 -3.119227719799209e-19

R155_176 V155 V176 642.0854275975415
L155_176 V155 V176 -1.109699667169616e-11
C155_176 V155 V176 6.029503531075857e-20

R155_177 V155 V177 90.38497499584585
L155_177 V155 V177 1.977561597056143e-12
C155_177 V155 V177 1.6755655169411285e-20

R155_178 V155 V178 -190.38081780184473
L155_178 V155 V178 2.467482462382624e-12
C155_178 V155 V178 5.11402767189693e-20

R155_179 V155 V179 -39533.87507431534
L155_179 V155 V179 1.2628924251821325e-12
C155_179 V155 V179 2.718560541779202e-19

R155_180 V155 V180 103.13136824194007
L155_180 V155 V180 1.7330123313363742e-12
C155_180 V155 V180 1.0853736216292005e-19

R155_181 V155 V181 -269.7866556519067
L155_181 V155 V181 -3.691746207168899e-12
C155_181 V155 V181 4.460928607569644e-20

R155_182 V155 V182 -82.66798419694265
L155_182 V155 V182 -1.438882731394261e-12
C155_182 V155 V182 -1.6930003847531076e-19

R155_183 V155 V183 1162.9699683314157
L155_183 V155 V183 1.5262556705659926e-12
C155_183 V155 V183 2.6620275892950442e-20

R155_184 V155 V184 -169.00138574610375
L155_184 V155 V184 3.760329494159735e-12
C155_184 V155 V184 -1.106686093481726e-20

R155_185 V155 V185 -142.58580964256336
L155_185 V155 V185 -3.928776754610826e-12
C155_185 V155 V185 -5.2818505580772205e-20

R155_186 V155 V186 371.64743847017684
L155_186 V155 V186 5.089569049459351e-12
C155_186 V155 V186 1.2565722970438433e-19

R155_187 V155 V187 108.26533707476403
L155_187 V155 V187 -7.989001401547581e-13
C155_187 V155 V187 -3.562859369374007e-19

R155_188 V155 V188 -71.46130892120895
L155_188 V155 V188 -1.2301536999258452e-12
C155_188 V155 V188 -2.0962031085461438e-19

R155_189 V155 V189 124.69067442469768
L155_189 V155 V189 6.317112607554105e-12
C155_189 V155 V189 -4.607659967146025e-20

R155_190 V155 V190 100.94729345348486
L155_190 V155 V190 5.562266693102144e-12
C155_190 V155 V190 1.2015536841631696e-19

R155_191 V155 V191 282.42557423969686
L155_191 V155 V191 -3.1604713004939626e-12
C155_191 V155 V191 3.2865504426067215e-19

R155_192 V155 V192 70.71982353219133
L155_192 V155 V192 -3.0271502377957977e-12
C155_192 V155 V192 9.872139961038739e-21

R155_193 V155 V193 184.9056314603566
L155_193 V155 V193 2.1106747999353014e-11
C155_193 V155 V193 7.984530935165759e-20

R155_194 V155 V194 -307.0966864547798
L155_194 V155 V194 2.8303123684540517e-11
C155_194 V155 V194 1.0444410006136949e-19

R155_195 V155 V195 -54.06481080846346
L155_195 V155 V195 2.2889817844936484e-12
C155_195 V155 V195 -4.1990549028982304e-19

R155_196 V155 V196 75.19681929182227
L155_196 V155 V196 8.651983941817996e-13
C155_196 V155 V196 5.42604960817123e-19

R155_197 V155 V197 -1200.351762701138
L155_197 V155 V197 7.470173996523825e-12
C155_197 V155 V197 1.0292070269234567e-19

R155_198 V155 V198 2101.877986549243
L155_198 V155 V198 -7.464628524365168e-12
C155_198 V155 V198 -4.402684478144892e-20

R155_199 V155 V199 -2311.6721740032685
L155_199 V155 V199 8.934538463314434e-12
C155_199 V155 V199 -2.4701737980776396e-20

R155_200 V155 V200 -113.14030194500297
L155_200 V155 V200 -5.183954849121728e-12
C155_200 V155 V200 -2.3028079910192265e-19

R156_156 V156 0 32.2349739696506
L156_156 V156 0 1.2248799368422612e-11
C156_156 V156 0 -1.9420664092804012e-18

R156_157 V156 V157 -56.38725403145255
L156_157 V156 V157 1.3459669840265531e-10
C156_157 V156 V157 5.463657065498587e-19

R156_158 V156 V158 30.888711746490788
L156_158 V156 V158 6.627502184891869e-12
C156_158 V156 V158 -7.495107630040749e-20

R156_159 V156 V159 -111.23143214347
L156_159 V156 V159 -1.4349622336957222e-11
C156_159 V156 V159 -2.379402211715729e-19

R156_160 V156 V160 -37.936859608071686
L156_160 V156 V160 -8.930662751224106e-12
C156_160 V156 V160 3.7693849701883303e-19

R156_161 V156 V161 40.88795396157943
L156_161 V156 V161 3.767687283160262e-12
C156_161 V156 V161 -4.349329292369539e-20

R156_162 V156 V162 195.92254533854427
L156_162 V156 V162 -1.3588139674217535e-11
C156_162 V156 V162 -7.659705647372289e-20

R156_163 V156 V163 130.53233948592015
L156_163 V156 V163 -8.81278666439241e-12
C156_163 V156 V163 1.5416782234151384e-19

R156_164 V156 V164 13.447200160083419
L156_164 V156 V164 6.504641182507352e-13
C156_164 V156 V164 -2.164905620476643e-19

R156_165 V156 V165 156.2368694452375
L156_165 V156 V165 4.53401300754216e-12
C156_165 V156 V165 -1.0720310208038806e-19

R156_166 V156 V166 -21.57317983353865
L156_166 V156 V166 3.3726302783766523e-11
C156_166 V156 V166 2.0872380634860746e-19

R156_167 V156 V167 73.78376358121297
L156_167 V156 V167 2.7746939047825014e-12
C156_167 V156 V167 -2.953078735900638e-20

R156_168 V156 V168 -88.00317687705235
L156_168 V156 V168 -1.0755918366454355e-12
C156_168 V156 V168 1.2031079716240518e-19

R156_169 V156 V169 -47.70354460674576
L156_169 V156 V169 -2.555634752437372e-12
C156_169 V156 V169 1.4993024807755185e-19

R156_170 V156 V170 39.38242289681674
L156_170 V156 V170 -2.4763041089790382e-11
C156_170 V156 V170 -1.214943093622408e-19

R156_171 V156 V171 -159.0142334674652
L156_171 V156 V171 -3.714234921496358e-12
C156_171 V156 V171 -1.1569963769994274e-19

R156_172 V156 V172 -18.76241673859913
L156_172 V156 V172 -2.895356030365929e-12
C156_172 V156 V172 3.9168063220768694e-20

R156_173 V156 V173 127.14183630264097
L156_173 V156 V173 -1.6571983601089205e-11
C156_173 V156 V173 -1.1730014197861754e-19

R156_174 V156 V174 38.18582664164697
L156_174 V156 V174 -6.086722195844112e-12
C156_174 V156 V174 1.445284799577185e-20

R156_175 V156 V175 -59.737735835747955
L156_175 V156 V175 -4.037345184847714e-12
C156_175 V156 V175 6.623353553434261e-20

R156_176 V156 V176 30.991438090191128
L156_176 V156 V176 1.7660454164343185e-12
C156_176 V156 V176 -5.900963377398259e-19

R156_177 V156 V177 114.06210938699537
L156_177 V156 V177 5.4176354254158934e-12
C156_177 V156 V177 7.772575026332215e-20

R156_178 V156 V178 -39.66214768227148
L156_178 V156 V178 1.3198701567907567e-11
C156_178 V156 V178 8.40436989258178e-20

R156_179 V156 V179 218.11399902986025
L156_179 V156 V179 5.947737614715103e-12
C156_179 V156 V179 1.1373273569580088e-19

R156_180 V156 V180 37.69331648201363
L156_180 V156 V180 3.6816579703044886e-12
C156_180 V156 V180 5.116440019066436e-19

R156_181 V156 V181 -95.46217111727036
L156_181 V156 V181 1.6730401178318458e-11
C156_181 V156 V181 1.0388537093994335e-19

R156_182 V156 V182 -62.06627236806655
L156_182 V156 V182 -9.507806739329236e-12
C156_182 V156 V182 -5.151852330116212e-20

R156_183 V156 V183 354.1946691418071
L156_183 V156 V183 5.584985804650518e-12
C156_183 V156 V183 1.2233908122208145e-19

R156_184 V156 V184 -25.886954953886676
L156_184 V156 V184 -1.8565011494376592e-12
C156_184 V156 V184 -7.101749028728183e-20

R156_185 V156 V185 -213.31861336096074
L156_185 V156 V185 -5.569294123149232e-12
C156_185 V156 V185 -1.327324327610016e-19

R156_186 V156 V186 -443.548645888229
L156_186 V156 V186 1.029860124113716e-10
C156_186 V156 V186 1.2954789010820619e-20

R156_187 V156 V187 -118.5929425158717
L156_187 V156 V187 -5.177708712404111e-12
C156_187 V156 V187 -1.0202867623503236e-19

R156_188 V156 V188 33.687834703233364
L156_188 V156 V188 2.906133729075955e-12
C156_188 V156 V188 -2.6933407892328466e-19

R156_189 V156 V189 297.72697733563524
L156_189 V156 V189 -5.94477867672516e-12
C156_189 V156 V189 -1.6507095288436063e-20

R156_190 V156 V190 123.05428383404796
L156_190 V156 V190 -1.0911805007628336e-11
C156_190 V156 V190 7.510935579173788e-20

R156_191 V156 V191 127.87622369315768
L156_191 V156 V191 -5.432575561581414e-12
C156_191 V156 V191 -2.5811287084757315e-19

R156_192 V156 V192 125.59985202504717
L156_192 V156 V192 2.1456920746153672e-11
C156_192 V156 V192 3.244333765832919e-19

R156_193 V156 V193 158.99018219866485
L156_193 V156 V193 5.997463772456975e-12
C156_193 V156 V193 9.952234908219096e-20

R156_194 V156 V194 -5783.1889248034595
L156_194 V156 V194 -1.0220384147911513e-11
C156_194 V156 V194 2.0107152769902845e-19

R156_195 V156 V195 -616.1668138693066
L156_195 V156 V195 3.653807018706258e-12
C156_195 V156 V195 6.556092882872204e-19

R156_196 V156 V196 -38.82395589232296
L156_196 V156 V196 -1.9171240879739448e-12
C156_196 V156 V196 -7.035806662692073e-19

R156_197 V156 V197 -239.87011709745974
L156_197 V156 V197 8.9485745583432e-12
C156_197 V156 V197 2.3150828180309894e-20

R156_198 V156 V198 -165.78319883246024
L156_198 V156 V198 -6.39351659085291e-11
C156_198 V156 V198 5.586129305228136e-20

R156_199 V156 V199 426.5752455247226
L156_199 V156 V199 -8.98740603057005e-12
C156_199 V156 V199 -7.713820619013945e-20

R156_200 V156 V200 -1641.8743436016039
L156_200 V156 V200 2.493034478293497e-12
C156_200 V156 V200 2.293630933059746e-19

R157_157 V157 0 34.75553966687975
L157_157 V157 0 1.3383515867729183e-13
C157_157 V157 0 5.27601277405586e-18

R157_158 V157 V158 276.0033636901951
L157_158 V157 V158 1.8720310257855815e-12
C157_158 V157 V158 -2.147853279946081e-20

R157_159 V157 V159 238.8722374083252
L157_159 V157 V159 -3.737372008903123e-12
C157_159 V157 V159 2.4534617186244614e-20

R157_160 V157 V160 82.58459627555487
L157_160 V157 V160 1.93244074516856e-12
C157_160 V157 V160 1.8452248545861527e-19

R157_161 V157 V161 49.47227532653218
L157_161 V157 V161 1.9460090317387714e-12
C157_161 V157 V161 -2.331542174201693e-20

R157_162 V157 V162 33.3036099123799
L157_162 V157 V162 7.842124722791591e-13
C157_162 V157 V162 5.721205611644764e-20

R157_163 V157 V163 46.4467154186625
L157_163 V157 V163 -9.581122199651533e-13
C157_163 V157 V163 -7.376369398067261e-19

R157_164 V157 V164 50.21101382348
L157_164 V157 V164 -1.8084352036103439e-12
C157_164 V157 V164 -1.0348578291603887e-19

R157_165 V157 V165 40.26244004067685
L157_165 V157 V165 3.3026597561677297e-13
C157_165 V157 V165 1.6882374018007768e-18

R157_166 V157 V166 -145.5512071656131
L157_166 V157 V166 -2.6861801986448656e-12
C157_166 V157 V166 -2.930671128540077e-19

R157_167 V157 V167 -99.4671841450933
L157_167 V157 V167 -3.0019202199722697e-12
C157_167 V157 V167 -8.675534304447029e-21

R157_168 V157 V168 -236.47248569159
L157_168 V157 V168 -1.2114955848815285e-11
C157_168 V157 V168 -4.1339287556293927e-19

R157_169 V157 V169 -52.09557054086097
L157_169 V157 V169 -7.333944196966329e-12
C157_169 V157 V169 -2.2194670997788447e-19

R157_170 V157 V170 -42.39882201105988
L157_170 V157 V170 4.587040217317492e-12
C157_170 V157 V170 8.432423113967924e-19

R157_171 V157 V171 -56.547497264503406
L157_171 V157 V171 4.126775933658473e-13
C157_171 V157 V171 1.2343730006591446e-18

R157_172 V157 V172 -48.47518556225159
L157_172 V157 V172 1.5143523186507333e-12
C157_172 V157 V172 8.028911750400382e-19

R157_173 V157 V173 -69.22532882376683
L157_173 V157 V173 -6.848729331027648e-13
C157_173 V157 V173 -6.780945664625189e-19

R157_174 V157 V174 58.09096718456726
L157_174 V157 V174 -4.692006469835286e-11
C157_174 V157 V174 -7.862736830900691e-19

R157_175 V157 V175 80.8418397014048
L157_175 V157 V175 4.595745111382186e-12
C157_175 V157 V175 6.337034618506354e-20

R157_176 V157 V176 75.70932592907415
L157_176 V157 V176 1.5033246183805073e-12
C157_176 V157 V176 2.1100450720385077e-19

R157_177 V157 V177 69.6999986372229
L157_177 V157 V177 -1.0322621062703466e-11
C157_177 V157 V177 3.7955336153792097e-19

R157_178 V157 V178 101.61591110350948
L157_178 V157 V178 -1.1926884827037303e-12
C157_178 V157 V178 -5.17845169068736e-19

R157_179 V157 V179 157.52332171425468
L157_179 V157 V179 -4.3288207617047587e-13
C157_179 V157 V179 -1.3077564297825736e-18

R157_180 V157 V180 73.22786911969044
L157_180 V157 V180 -4.815294179059211e-13
C157_180 V157 V180 -1.11111492024741e-18

R157_181 V157 V181 376.6562472279197
L157_181 V157 V181 3.101398767177775e-12
C157_181 V157 V181 -2.1167257192580757e-19

R157_182 V157 V182 -59.20559842327797
L157_182 V157 V182 4.1385705206894656e-13
C157_182 V157 V182 8.923338208184556e-19

R157_183 V157 V183 -89.69683806178325
L157_183 V157 V183 -7.913640747359898e-13
C157_183 V157 V183 -1.719330808827625e-19

R157_184 V157 V184 -53.55476874591127
L157_184 V157 V184 -1.183324369109185e-12
C157_184 V157 V184 1.7752307390301174e-19

R157_185 V157 V185 -46.93042583887313
L157_185 V157 V185 -5.652550889935582e-12
C157_185 V157 V185 -1.2316578556140858e-19

R157_186 V157 V186 -11791.879247816321
L157_186 V157 V186 -1.2327283999456772e-11
C157_186 V157 V186 3.8750909787418454e-20

R157_187 V157 V187 205.28809892731766
L157_187 V157 V187 4.798806099911404e-13
C157_187 V157 V187 9.920942843733045e-19

R157_188 V157 V188 139.93503750554433
L157_188 V157 V188 3.1149398980988747e-13
C157_188 V157 V188 7.753498030482947e-19

R157_189 V157 V189 91.93179031183348
L157_189 V157 V189 1.1925516515179057e-12
C157_189 V157 V189 7.587597168195294e-19

R157_190 V157 V190 65.9758126385307
L157_190 V157 V190 -1.4845956269758037e-12
C157_190 V157 V190 -9.10372498638927e-19

R157_191 V157 V191 119.70984333585477
L157_191 V157 V191 4.205267285415266e-13
C157_191 V157 V191 6.765944123692892e-19

R157_192 V157 V192 100.34725102760731
L157_192 V157 V192 3.821979720874407e-12
C157_192 V157 V192 3.060597398576595e-19

R157_193 V157 V193 58.838948345404205
L157_193 V157 V193 -2.2411952844110845e-12
C157_193 V157 V193 -5.420877486966083e-19

R157_194 V157 V194 -60.79749558217816
L157_194 V157 V194 -2.577362319805221e-12
C157_194 V157 V194 -1.571139240460005e-19

R157_195 V157 V195 -70.88790652813361
L157_195 V157 V195 -2.6830077206407925e-13
C157_195 V157 V195 -1.478005532850977e-18

R157_196 V157 V196 -67.36033068116059
L157_196 V157 V196 -3.6093116687761466e-13
C157_196 V157 V196 -1.0300474145740615e-18

R157_197 V157 V197 -62.86411688615813
L157_197 V157 V197 -7.192367558179465e-13
C157_197 V157 V197 -3.9922214151903056e-19

R157_198 V157 V198 -193.79724813348068
L157_198 V157 V198 2.3313927584441414e-12
C157_198 V157 V198 1.528002114236584e-19

R157_199 V157 V199 -2989.431092130499
L157_199 V157 V199 -8.568554214809725e-13
C157_199 V157 V199 -6.473159320931307e-19

R157_200 V157 V200 -27174.698953713072
L157_200 V157 V200 -2.567816511073901e-12
C157_200 V157 V200 -1.187230509575118e-19

R158_158 V158 0 49.990952427579415
L158_158 V158 0 1.9269607409453035e-12
C158_158 V158 0 1.2608258516235327e-19

R158_159 V158 V159 34.47942339551688
L158_159 V158 V159 3.1241200234462966e-12
C158_159 V158 V159 7.881108298165389e-20

R158_160 V158 V160 25.241446403859687
L158_160 V158 V160 6.391377879736543e-11
C158_160 V158 V160 8.175605734971923e-20

R158_161 V158 V161 -23.644431794031995
L158_161 V158 V161 -5.601618467645707e-12
C158_161 V158 V161 -7.824817512466882e-20

R158_162 V158 V162 -29.88562064955264
L158_162 V158 V162 4.346229258409424e-12
C158_162 V158 V162 1.570418244734049e-20

R158_163 V158 V163 -34.982117347633384
L158_163 V158 V163 -7.906013449437458e-12
C158_163 V158 V163 -7.89483941671156e-20

R158_164 V158 V164 -21.201681988414098
L158_164 V158 V164 -6.563373621513972e-12
C158_164 V158 V164 -5.0223097719648474e-20

R158_165 V158 V165 -163.33188170400155
L158_165 V158 V165 -2.0609659085195442e-12
C158_165 V158 V165 7.694027627328784e-20

R158_166 V158 V166 5.094585279613231
L158_166 V158 V166 6.376992905194146e-13
C158_166 V158 V166 6.936870438090432e-20

R158_167 V158 V167 -19.586222595764387
L158_167 V158 V167 -3.4818834138399814e-12
C158_167 V158 V167 -2.765527059186919e-20

R158_168 V158 V168 -15.966927557178204
L158_168 V158 V168 -4.490882867793102e-12
C158_168 V158 V168 -3.246082223496498e-20

R158_169 V158 V169 21.254793505751454
L158_169 V158 V169 5.564636249389406e-12
C158_169 V158 V169 1.0239222269766222e-20

R158_170 V158 V170 -12.257578000057094
L158_170 V158 V170 -9.07432673277572e-13
C158_170 V158 V170 1.9177879315728082e-20

R158_171 V158 V171 23.643022650528962
L158_171 V158 V171 -1.703229098740669e-11
C158_171 V158 V171 9.167624316246566e-20

R158_172 V158 V172 19.473762893660894
L158_172 V158 V172 -9.915440851197924e-12
C158_172 V158 V172 8.098078338268017e-20

R158_173 V158 V173 -29.959076287941304
L158_173 V158 V173 -1.0284285505136222e-11
C158_173 V158 V173 -1.4904721108061953e-20

R158_174 V158 V174 -7.0860959449107055
L158_174 V158 V174 -1.8585773814393693e-12
C158_174 V158 V174 -3.56691506201168e-20

R158_175 V158 V175 39.28130028589652
L158_175 V158 V175 -2.2049463566199127e-11
C158_175 V158 V175 -7.899317882578205e-20

R158_176 V158 V176 25.737032134549082
L158_176 V158 V176 3.3069539645295034e-12
C158_176 V158 V176 -7.129188670619833e-20

R158_177 V158 V177 -48.30945272497037
L158_177 V158 V177 -9.720357113683576e-12
C158_177 V158 V177 5.708758672072457e-20

R158_178 V158 V178 10.712856590903533
L158_178 V158 V178 1.2700721056076751e-12
C158_178 V158 V178 -1.3323427900072055e-20

R158_179 V158 V179 -32.237078099657005
L158_179 V158 V179 9.732369055407902e-10
C158_179 V158 V179 2.7952963795703646e-20

R158_180 V158 V180 -20.419632284979677
L158_180 V158 V180 -1.0707739804823064e-11
C158_180 V158 V180 4.442501975676509e-20

R158_181 V158 V181 34.653331335026984
L158_181 V158 V181 4.264385652693111e-12
C158_181 V158 V181 -7.786147739795101e-20

R158_182 V158 V182 15.200632112952713
L158_182 V158 V182 -3.786392385162472e-12
C158_182 V158 V182 -2.9023661237760726e-21

R158_183 V158 V183 -2177.988163064071
L158_183 V158 V183 6.5424743808377175e-12
C158_183 V158 V183 -9.684200763385024e-21

R158_184 V158 V184 -1245.4185164780006
L158_184 V158 V184 -2.3925507623816116e-11
C158_184 V158 V184 1.256939308399064e-20

R158_185 V158 V185 295.95257513706883
L158_185 V158 V185 -7.093775679264142e-12
C158_185 V158 V185 -1.7479962347874005e-20

R158_186 V158 V186 -31.75276358688639
L158_186 V158 V186 -1.9438765534292108e-11
C158_186 V158 V186 -1.359757175070952e-20

R158_187 V158 V187 290.8865931921937
L158_187 V158 V187 -3.875811581855895e-12
C158_187 V158 V187 -3.9094727886431546e-20

R158_188 V158 V188 82.56883223999822
L158_188 V158 V188 6.819925166663175e-11
C158_188 V158 V188 -3.663873243192112e-20

R158_189 V158 V189 -93.02709732970924
L158_189 V158 V189 -3.0511242049860586e-12
C158_189 V158 V189 1.2574566792735149e-19

R158_190 V158 V190 -32.27538405354164
L158_190 V158 V190 -1.0562345212088925e-11
C158_190 V158 V190 -2.1776449466173934e-20

R158_191 V158 V191 -3055.7858451906163
L158_191 V158 V191 -3.715357413125598e-12
C158_191 V158 V191 1.3539408937258234e-19

R158_192 V158 V192 491.1517833543695
L158_192 V158 V192 -2.4267720912289833e-12
C158_192 V158 V192 1.4468569497724416e-19

R158_193 V158 V193 -531.0105194489832
L158_193 V158 V193 3.804851984646735e-12
C158_193 V158 V193 -7.155630733852666e-21

R158_194 V158 V194 185.29927725658075
L158_194 V158 V194 -3.770638798791369e-12
C158_194 V158 V194 2.9791327010685214e-20

R158_195 V158 V195 178.0130421739018
L158_195 V158 V195 4.544685905335185e-12
C158_195 V158 V195 -1.764979447956467e-19

R158_196 V158 V196 -274.14527905623703
L158_196 V158 V196 1.7855516346856619e-12
C158_196 V158 V196 -1.9477697015868363e-19

R158_197 V158 V197 352.2335868537645
L158_197 V158 V197 5.511916769897466e-12
C158_197 V158 V197 -7.816886619362353e-20

R158_198 V158 V198 21.85303655423933
L158_198 V158 V198 2.303025246224699e-12
C158_198 V158 V198 4.6754081064574054e-20

R158_199 V158 V199 -1989.5797041638016
L158_199 V158 V199 4.083205854204983e-12
C158_199 V158 V199 -9.738536346508615e-20

R158_200 V158 V200 -80.54774402534639
L158_200 V158 V200 1.567999598579572e-11
C158_200 V158 V200 -1.3533547483731117e-20

R159_159 V159 0 32.23579929552827
L159_159 V159 0 -5.01723506214151e-13
C159_159 V159 0 -3.6060159018864875e-19

R159_160 V159 V160 35.71375455253625
L159_160 V159 V160 1.7911568783834563e-12
C159_160 V159 V160 1.6355598760728045e-19

R159_161 V159 V161 98.87364954370909
L159_161 V159 V161 2.7465903832564178e-12
C159_161 V159 V161 3.1289466113547707e-19

R159_162 V159 V162 -517.9558375914908
L159_162 V159 V162 3.912099967407972e-12
C159_162 V159 V162 3.058728900996158e-20

R159_163 V159 V163 29.710529661646095
L159_163 V159 V163 1.0244492124269327e-12
C159_163 V159 V163 4.130057905248713e-19

R159_164 V159 V164 -2212.9214009154693
L159_164 V159 V164 -7.596683607225766e-11
C159_164 V159 V164 1.1044766115264017e-20

R159_165 V159 V165 -70.02535479831245
L159_165 V159 V165 2.404140384965834e-12
C159_165 V159 V165 -1.067389635245867e-19

R159_166 V159 V166 -17.389884213057407
L159_166 V159 V166 -5.740498661796756e-12
C159_166 V159 V166 5.0656009551638285e-20

R159_167 V159 V167 11.210455679352474
L159_167 V159 V167 4.897463368491094e-13
C159_167 V159 V167 7.059769410951233e-21

R159_168 V159 V168 -63.331534249780205
L159_168 V159 V168 -3.1264421740355274e-12
C159_168 V159 V168 2.5733926966562798e-19

R159_169 V159 V169 -49.83126011037535
L159_169 V159 V169 -1.0455338755377265e-12
C159_169 V159 V169 -3.994495353599892e-19

R159_170 V159 V170 54.20636107094213
L159_170 V159 V170 -1.0499347334503727e-11
C159_170 V159 V170 -2.608981696589128e-21

R159_171 V159 V171 -16.740183109716394
L159_171 V159 V171 -8.095804634493456e-13
C159_171 V159 V171 -1.1214379021190027e-19

R159_172 V159 V172 -246.23428402869317
L159_172 V159 V172 2.793330339327696e-11
C159_172 V159 V172 -1.1739726025895572e-19

R159_173 V159 V173 41.08347747741403
L159_173 V159 V173 4.6460030240834034e-12
C159_173 V159 V173 1.5779419120085705e-19

R159_174 V159 V174 19.629376407060217
L159_174 V159 V174 -8.504001391889115e-11
C159_174 V159 V174 -2.1229526533498234e-19

R159_175 V159 V175 -26.855833357714136
L159_175 V159 V175 1.3659303979226726e-11
C159_175 V159 V175 2.894433803670156e-19

R159_176 V159 V176 156.34688760589228
L159_176 V159 V176 -3.0303387206284283e-12
C159_176 V159 V176 -3.4498381663173564e-19

R159_177 V159 V177 202.13745765479567
L159_177 V159 V177 6.526139911719923e-12
C159_177 V159 V177 5.269238409158094e-20

R159_178 V159 V178 -38.72546166531508
L159_178 V159 V178 -5.60291382168035e-12
C159_178 V159 V178 9.194294569268351e-20

R159_179 V159 V179 23.026857420996357
L159_179 V159 V179 3.657032845843293e-12
C159_179 V159 V179 -1.671746304949095e-19

R159_180 V159 V180 111.74079099630633
L159_180 V159 V180 1.3606655367410144e-11
C159_180 V159 V180 2.0629134477881972e-19

R159_181 V159 V181 -71.70456673725563
L159_181 V159 V181 7.37225926834944e-12
C159_181 V159 V181 1.7323685841327047e-19

R159_182 V159 V182 -37.02142369458807
L159_182 V159 V182 2.7763263256014597e-12
C159_182 V159 V182 4.669770343764476e-20

R159_183 V159 V183 751.8466770682536
L159_183 V159 V183 -1.6726006406535588e-12
C159_183 V159 V183 3.1233518182435714e-20

R159_184 V159 V184 -188.9280732867521
L159_184 V159 V184 -5.777967781839934e-12
C159_184 V159 V184 -8.861437958732614e-21

R159_185 V159 V185 420.9672170394933
L159_185 V159 V185 4.255585194967704e-12
C159_185 V159 V185 -1.46622077359386e-19

R159_186 V159 V186 151.14130906328205
L159_186 V159 V186 4.309605247000712e-12
C159_186 V159 V186 -2.950838493971575e-20

R159_187 V159 V187 -159.77553995678412
L159_187 V159 V187 8.257837313036309e-13
C159_187 V159 V187 3.1603637620273483e-19

R159_188 V159 V188 544.2228128478481
L159_188 V159 V188 2.269593156389341e-12
C159_188 V159 V188 7.269919126894983e-20

R159_189 V159 V189 322.2849891804626
L159_189 V159 V189 -1.4809813163021098e-12
C159_189 V159 V189 -1.6650838251670015e-19

R159_190 V159 V190 93.71380568961338
L159_190 V159 V190 -5.427454659941646e-12
C159_190 V159 V190 3.5189867510253937e-20

R159_191 V159 V191 -273.7798630824947
L159_191 V159 V191 -5.818925867209965e-12
C159_191 V159 V191 -4.782095895590127e-19

R159_192 V159 V192 120.54329231354866
L159_192 V159 V192 4.361689558171325e-12
C159_192 V159 V192 -8.249785505498362e-20

R159_193 V159 V193 263.4289315921247
L159_193 V159 V193 -4.1348452351011756e-11
C159_193 V159 V193 2.7370450779234804e-20

R159_194 V159 V194 4472.124770320723
L159_194 V159 V194 -2.168244791981354e-12
C159_194 V159 V194 -2.456404558616237e-19

R159_195 V159 V195 -128.35467998604864
L159_195 V159 V195 -8.624476141981393e-12
C159_195 V159 V195 7.22342323669865e-19

R159_196 V159 V196 -197.03987417455596
L159_196 V159 V196 -7.08582482430466e-13
C159_196 V159 V196 -4.556686350350999e-19

R159_197 V159 V197 673.5144505915199
L159_197 V159 V197 2.639499897956612e-12
C159_197 V159 V197 2.1130683150334846e-19

R159_198 V159 V198 -50.30079963165972
L159_198 V159 V198 4.597799579639358e-12
C159_198 V159 V198 2.2275921843442212e-20

R159_199 V159 V199 211.74423981273702
L159_199 V159 V199 3.205357326830972e-12
C159_199 V159 V199 1.48024532424594e-20

R159_200 V159 V200 165.6549621717326
L159_200 V159 V200 1.527958339235558e-12
C159_200 V159 V200 4.2315518175052106e-19

R160_160 V160 0 -14.378561576023595
L160_160 V160 0 -5.186616057946964e-13
C160_160 V160 0 -3.13958394370991e-20

R160_161 V160 V161 114.8673141641332
L160_161 V160 V161 2.9505229494198018e-12
C160_161 V160 V161 1.5635260035854778e-19

R160_162 V160 V162 -791.9978436263245
L160_162 V160 V162 -5.441078343427987e-12
C160_162 V160 V162 1.2184863201831878e-20

R160_163 V160 V163 148.81033987766526
L160_163 V160 V163 -6.542849367376651e-12
C160_163 V160 V163 -8.908729658881147e-21

R160_164 V160 V164 10.989100824894878
L160_164 V160 V164 8.774993766472956e-13
C160_164 V160 V164 2.8839927696544967e-19

R160_165 V160 V165 -219.62107903958085
L160_165 V160 V165 -3.5640814728285906e-12
C160_165 V160 V165 -2.411009503867301e-19

R160_166 V160 V166 -16.86700744452239
L160_166 V160 V166 -3.9160220331201846e-12
C160_166 V160 V166 -4.1849829554703843e-20

R160_167 V160 V167 -75.39392821993772
L160_167 V160 V167 -2.495001278418119e-12
C160_167 V160 V167 1.2819804268244757e-19

R160_168 V160 V168 10.603969012844242
L160_168 V160 V168 4.373836778933894e-13
C160_168 V160 V168 1.114055689350424e-19

R160_169 V160 V169 -50.17329996230086
L160_169 V160 V169 -1.660123874035656e-12
C160_169 V160 V169 -1.5475175132087156e-19

R160_170 V160 V170 37.62732858370337
L160_170 V160 V170 4.645389794277178e-12
C160_170 V160 V170 -5.928749446285995e-20

R160_171 V160 V171 -177.16041378021558
L160_171 V160 V171 6.21566137022009e-12
C160_171 V160 V171 -1.3099560745174678e-19

R160_172 V160 V172 -11.966316886268924
L160_172 V160 V172 -6.023503650444584e-13
C160_172 V160 V172 -2.7508284457087663e-19

R160_173 V160 V173 40.45179510190513
L160_173 V160 V173 2.4446385457292386e-12
C160_173 V160 V173 1.864317340853156e-19

R160_174 V160 V174 19.874736149267598
L160_174 V160 V174 -1.0871519203781014e-11
C160_174 V160 V174 4.01815168233997e-20

R160_175 V160 V175 137.26718165290913
L160_175 V160 V175 -3.06477353263719e-12
C160_175 V160 V175 -1.9008909741654906e-19

R160_176 V160 V176 -31.177145491643095
L160_176 V160 V176 -3.428406197030263e-12
C160_176 V160 V176 3.853195284065843e-19

R160_177 V160 V177 64.16998160641668
L160_177 V160 V177 4.2981889522643775e-12
C160_177 V160 V177 -4.4841920936951185e-20

R160_178 V160 V178 -31.231935835448674
L160_178 V160 V178 -1.3374804509108738e-11
C160_178 V160 V178 4.840948381151676e-20

R160_179 V160 V179 -726.5126981994973
L160_179 V160 V179 2.8733692335324767e-11
C160_179 V160 V179 1.8231865452141962e-19

R160_180 V160 V180 21.711316153223503
L160_180 V160 V180 1.929804298879777e-12
C160_180 V160 V180 -2.238967872514393e-19

R160_181 V160 V181 -44.29321303502305
L160_181 V160 V181 -5.711814428323127e-12
C160_181 V160 V181 8.856116327144425e-20

R160_182 V160 V182 -27.59818423929902
L160_182 V160 V182 -3.301486247822756e-12
C160_182 V160 V182 -1.234803447088627e-19

R160_183 V160 V183 -150.24102150785052
L160_183 V160 V183 -1.1064882253507424e-11
C160_183 V160 V183 -6.589207083505833e-20

R160_184 V160 V184 -246.32535411104593
L160_184 V160 V184 -6.328920293089205e-11
C160_184 V160 V184 5.544245621977631e-20

R160_185 V160 V185 -521.735933161069
L160_185 V160 V185 7.159525906441816e-12
C160_185 V160 V185 -3.335724929843501e-20

R160_186 V160 V186 259.2508887422548
L160_186 V160 V186 1.1489512857628042e-11
C160_186 V160 V186 7.145583520939616e-20

R160_187 V160 V187 -620.764652860804
L160_187 V160 V187 -6.948220737193056e-12
C160_187 V160 V187 -1.237344000624475e-19

R160_188 V160 V188 220.26125614221806
L160_188 V160 V188 1.5653064903459528e-12
C160_188 V160 V188 1.1384855296297865e-19

R160_189 V160 V189 101.82326357000034
L160_189 V160 V189 -1.976522798250743e-12
C160_189 V160 V189 -2.049615322438106e-19

R160_190 V160 V190 41.64245113330497
L160_190 V160 V190 6.336222056149326e-12
C160_190 V160 V190 1.3208078774132316e-19

R160_191 V160 V191 67.14761336767846
L160_191 V160 V191 3.5474789856927073e-12
C160_191 V160 V191 1.0808691250129491e-19

R160_192 V160 V192 -63.599945726976394
L160_192 V160 V192 -9.899358194093917e-13
C160_192 V160 V192 -4.1986025540160745e-19

R160_193 V160 V193 6565.701613772114
L160_193 V160 V193 -1.2883423060527176e-11
C160_193 V160 V193 2.882337119104684e-20

R160_194 V160 V194 -245.96725683382837
L160_194 V160 V194 -1.671662241010233e-12
C160_194 V160 V194 -2.2618704769646814e-19

R160_195 V160 V195 -184.54912971280817
L160_195 V160 V195 -2.5384645090036205e-12
C160_195 V160 V195 -2.648509560715361e-19

R160_196 V160 V196 336.5396123965226
L160_196 V160 V196 1.230194703837409e-12
C160_196 V160 V196 8.604658328948599e-19

R160_197 V160 V197 -105.17936650777645
L160_197 V160 V197 1.930508396700033e-12
C160_197 V160 V197 2.2492195621627563e-19

R160_198 V160 V198 -75.56900032560307
L160_198 V160 V198 2.117150486733526e-11
C160_198 V160 V198 -5.593273794364333e-20

R160_199 V160 V199 89.23549846918094
L160_199 V160 V199 4.35947575191898e-12
C160_199 V160 V199 2.1725130633485575e-19

R160_200 V160 V200 103.74383404981747
L160_200 V160 V200 2.9740024159675163e-12
C160_200 V160 V200 -1.747250806878433e-19

R161_161 V161 0 -47.43627957762754
L161_161 V161 0 3.876281889338726e-13
C161_161 V161 0 7.478946468324774e-19

R161_162 V161 V162 -57.88725151349286
L161_162 V161 V162 -1.729639474361527e-12
C161_162 V161 V162 8.264759798841541e-20

R161_163 V161 V163 -38.45369048209899
L161_163 V161 V163 -1.6592611100588981e-12
C161_163 V161 V163 -5.876935467791802e-20

R161_164 V161 V164 -29.29361233326833
L161_164 V161 V164 -1.4214201771708401e-12
C161_164 V161 V164 -1.712937266189022e-19

R161_165 V161 V165 -139.23016992828153
L161_165 V161 V165 1.96072215384038e-12
C161_165 V161 V165 2.773025348539077e-19

R161_166 V161 V166 15.085879744418014
L161_166 V161 V166 5.8680686320047985e-12
C161_166 V161 V166 -1.79613386009928e-19

R161_167 V161 V167 -527.8155673156008
L161_167 V161 V167 -4.1693361427235925e-12
C161_167 V161 V167 -2.883600847564393e-19

R161_168 V161 V168 -87.90916832702173
L161_168 V161 V168 -1.5569757464193828e-12
C161_168 V161 V168 -3.5909055568973377e-19

R161_169 V161 V169 27.3586091772416
L161_169 V161 V169 9.479949467074135e-13
C161_169 V161 V169 6.113311270054267e-19

R161_170 V161 V170 -52.205691664737536
L161_170 V161 V170 9.055225262886577e-11
C161_170 V161 V170 7.546212888435864e-20

R161_171 V161 V171 50.21972046069542
L161_171 V161 V171 3.729446056912684e-12
C161_171 V161 V171 1.2499502719095473e-19

R161_172 V161 V172 40.24215304198697
L161_172 V161 V172 1.0468954270688984e-12
C161_172 V161 V172 2.8673424373856146e-19

R161_173 V161 V173 -50.29350885463694
L161_173 V161 V173 -2.132547581046724e-12
C161_173 V161 V173 4.1187513337888303e-20

R161_174 V161 V174 -21.956351091065994
L161_174 V161 V174 1.7637880899205116e-12
C161_174 V161 V174 3.873123371806731e-19

R161_175 V161 V175 -5526.15054630803
L161_175 V161 V175 2.4952725317281825e-12
C161_175 V161 V175 1.984104587736456e-19

R161_176 V161 V176 667.5189345811605
L161_176 V161 V176 1.0367235848158287e-11
C161_176 V161 V176 2.107808584464003e-19

R161_177 V161 V177 -77.01144596847028
L161_177 V161 V177 1.0500538177470269e-11
C161_177 V161 V177 -2.7620239685400665e-19

R161_178 V161 V178 48.47665995753955
L161_178 V161 V178 -4.293942311434949e-12
C161_178 V161 V178 -1.8352877888217285e-19

R161_179 V161 V179 -81.57234004451084
L161_179 V161 V179 -3.6278807907111694e-12
C161_179 V161 V179 -3.742687052299087e-20

R161_180 V161 V180 -61.390069777453704
L161_180 V161 V180 -2.4581158435479642e-12
C161_180 V161 V180 -1.5124006623718925e-19

R161_181 V161 V181 69.82811966165906
L161_181 V161 V181 -3.5616786092370058e-12
C161_181 V161 V181 -3.452287709722256e-19

R161_182 V161 V182 31.108972998163523
L161_182 V161 V182 6.789121810322077e-12
C161_182 V161 V182 1.3491979839280501e-20

R161_183 V161 V183 193.68378842917375
L161_183 V161 V183 4.543970369057332e-12
C161_183 V161 V183 1.8323501378790585e-20

R161_184 V161 V184 190.31897018478372
L161_184 V161 V184 4.648138478327855e-12
C161_184 V161 V184 -4.2026861197054317e-20

R161_185 V161 V185 163.1846571501678
L161_185 V161 V185 -2.3359766245077193e-12
C161_185 V161 V185 2.936727642769329e-19

R161_186 V161 V186 -297.20634365166035
L161_186 V161 V186 1.0921769391185823e-11
C161_186 V161 V186 -1.9881016995035125e-19

R161_187 V161 V187 -1365.803077363472
L161_187 V161 V187 -3.034080765506276e-12
C161_187 V161 V187 -2.3874496632297157e-19

R161_188 V161 V188 -315.8862602246285
L161_188 V161 V188 -8.542160682583437e-13
C161_188 V161 V188 -2.5408693240750143e-19

R161_189 V161 V189 -184.46135692573375
L161_189 V161 V189 1.4159279837137308e-12
C161_189 V161 V189 1.216085514397871e-19

R161_190 V161 V190 -61.963088668352746
L161_190 V161 V190 -8.325037498385726e-12
C161_190 V161 V190 -3.240033696555806e-20

R161_191 V161 V191 -256.55766465165703
L161_191 V161 V191 -3.909037952198303e-12
C161_191 V161 V191 1.308558744569327e-19

R161_192 V161 V192 -426.61499611392406
L161_192 V161 V192 1.120537868204479e-12
C161_192 V161 V192 4.593894413681559e-19

R161_193 V161 V193 -118.2294505299644
L161_193 V161 V193 -8.602845500583842e-12
C161_193 V161 V193 2.461542816759802e-19

R161_194 V161 V194 136.12908666711127
L161_194 V161 V194 1.0129745221719855e-12
C161_194 V161 V194 5.643409722261922e-19

R161_195 V161 V195 156.67121795396696
L161_195 V161 V195 2.415253277529659e-12
C161_195 V161 V195 -7.418350722675022e-20

R161_196 V161 V196 194.78523578943577
L161_196 V161 V196 -3.4553040202354707e-12
C161_196 V161 V196 -2.4449771215061215e-19

R161_197 V161 V197 239.7842667139866
L161_197 V161 V197 -2.7006014163051213e-12
C161_197 V161 V197 -4.853352753497686e-19

R161_198 V161 V198 47.586376828951096
L161_198 V161 V198 -1.2015989807562248e-11
C161_198 V161 V198 -4.2252835443625906e-21

R161_199 V161 V199 202.01997252882504
L161_199 V161 V199 -2.868895836391438e-12
C161_199 V161 V199 3.799212141805619e-20

R161_200 V161 V200 -142.35375937561432
L161_200 V161 V200 -1.6130760786207884e-12
C161_200 V161 V200 -2.7898943962398644e-19

R162_162 V162 0 167.21330851077101
L162_162 V162 0 -4.419890793907956e-13
C162_162 V162 0 -7.69578220521908e-19

R162_163 V162 V163 -132.6755510161807
L162_163 V162 V163 -9.237120899415993e-12
C162_163 V162 V163 -1.083180462901196e-19

R162_164 V162 V164 -187.14192391401315
L162_164 V162 V164 1.1523586430024438e-11
C162_164 V162 V164 -7.114434701759203e-20

R162_165 V162 V165 -40.53775061269999
L162_165 V162 V165 -3.9751120373023846e-12
C162_165 V162 V165 1.097276799727139e-19

R162_166 V162 V166 17.266416910281176
L162_166 V162 V166 1.912359814467334e-12
C162_166 V162 V166 9.66099247799147e-20

R162_167 V162 V167 -66.56029694695593
L162_167 V162 V167 -9.81283501432065e-12
C162_167 V162 V167 5.606198295053534e-20

R162_168 V162 V168 -36.725436045818704
L162_168 V162 V168 -2.2262196165365315e-12
C162_168 V162 V168 1.0846563475063914e-19

R162_169 V162 V169 50.977155813947554
L162_169 V162 V169 2.4446939055183977e-12
C162_169 V162 V169 -1.5018226029931502e-20

R162_170 V162 V170 50.92745699705711
L162_170 V162 V170 1.1680529485193438e-12
C162_170 V162 V170 1.5624454111644796e-20

R162_171 V162 V171 67.9723732078095
L162_171 V162 V171 -1.3210042469201178e-11
C162_171 V162 V171 5.826185455853234e-20

R162_172 V162 V172 53.95661820083095
L162_172 V162 V172 2.8635861043981687e-12
C162_172 V162 V172 3.161746538428126e-20

R162_173 V162 V173 117.09564110682594
L162_173 V162 V173 -2.0049709663317957e-11
C162_173 V162 V173 -2.1585764665162354e-19

R162_174 V162 V174 -14.709697323907706
L162_174 V162 V174 -1.1989525775576353e-12
C162_174 V162 V174 -5.852901480673371e-20

R162_175 V162 V175 136.1441314119474
L162_175 V162 V175 -4.247380438873828e-12
C162_175 V162 V175 -2.0301137484684426e-19

R162_176 V162 V176 56.66209939010183
L162_176 V162 V176 -5.598725129225932e-12
C162_176 V162 V176 -1.8781698984887184e-19

R162_177 V162 V177 -74.89883578680826
L162_177 V162 V177 2.3940716230490572e-11
C162_177 V162 V177 5.664900701071294e-20

R162_178 V162 V178 366.1197079043676
L162_178 V162 V178 -1.80175431395068e-11
C162_178 V162 V178 2.1416412036068126e-20

R162_179 V162 V179 -109.68977614258759
L162_179 V162 V179 2.645066406644999e-12
C162_179 V162 V179 1.2724231335964197e-19

R162_180 V162 V180 -49.17007619417414
L162_180 V162 V180 4.132983408958493e-12
C162_180 V162 V180 9.318121335244148e-20

R162_181 V162 V181 1055.0741032115832
L162_181 V162 V181 -3.726684397701678e-12
C162_181 V162 V181 2.189918109151838e-19

R162_182 V162 V182 24.082315669286288
L162_182 V162 V182 2.883969414115013e-12
C162_182 V162 V182 -9.619568990723503e-21

R162_183 V162 V183 1871.7192065908955
L162_183 V162 V183 2.5889769677084025e-12
C162_183 V162 V183 3.81544943495639e-20

R162_184 V162 V184 563.639656180891
L162_184 V162 V184 3.384147126685778e-12
C162_184 V162 V184 7.369414774326028e-20

R162_185 V162 V185 67.41840558825491
L162_185 V162 V185 4.921561962816685e-12
C162_185 V162 V185 -1.3858249607977516e-19

R162_186 V162 V186 -144.04101809155375
L162_186 V162 V186 -6.494797792640588e-12
C162_186 V162 V186 1.159836341436523e-19

R162_187 V162 V187 -292.7480576402436
L162_187 V162 V187 -1.4668252768919794e-12
C162_187 V162 V187 -9.017765643850922e-20

R162_188 V162 V188 207.96148927383348
L162_188 V162 V188 -1.1335613290634967e-12
C162_188 V162 V188 -5.725979758198232e-20

R162_189 V162 V189 -111.7772116040206
L162_189 V162 V189 5.2093584510436e-12
C162_189 V162 V189 -4.886633102895445e-20

R162_190 V162 V190 -30.0078401218765
L162_190 V162 V190 -3.40113723448082e-12
C162_190 V162 V190 -1.6933853204429055e-20

R162_191 V162 V191 -429.93961979458675
L162_191 V162 V191 -2.7340501959208183e-12
C162_191 V162 V191 -4.951308262399845e-22

R162_192 V162 V192 -505.3243190184888
L162_192 V162 V192 5.102493188157112e-12
C162_192 V162 V192 -5.838133178588447e-20

R162_193 V162 V193 -88.53873436322563
L162_193 V162 V193 -4.384051847357238e-12
C162_193 V162 V193 -2.5328425673451863e-20

R162_194 V162 V194 56.00614202661271
L162_194 V162 V194 2.19984267241159e-12
C162_194 V162 V194 1.168107693352919e-20

R162_195 V162 V195 157.22655307643063
L162_195 V162 V195 1.460714997796559e-12
C162_195 V162 V195 -4.249987987159037e-21

R162_196 V162 V196 708.5633506411964
L162_196 V162 V196 4.746140197011112e-12
C162_196 V162 V196 -4.988361034279478e-22

R162_197 V162 V197 57.680210200680364
L162_197 V162 V197 4.680506751995636e-12
C162_197 V162 V197 9.061427498856729e-20

R162_198 V162 V198 40.385305509773644
L162_198 V162 V198 5.288597583990022e-12
C162_198 V162 V198 -3.1929012041267466e-20

R162_199 V162 V199 540.6675664665495
L162_199 V162 V199 8.12135454960303e-11
C162_199 V162 V199 -7.528532474616127e-20

R162_200 V162 V200 -1606.5258678561504
L162_200 V162 V200 -2.023689959597372e-11
C162_200 V162 V200 5.740627003808368e-20

R163_163 V163 0 -97.68973103262849
L163_163 V163 0 1.0465376730196502e-12
C163_163 V163 0 1.1137585183282541e-18

R163_164 V163 V164 -33.36512725848851
L163_164 V163 V164 -1.6244507110044062e-12
C163_164 V163 V164 -9.852173335085823e-20

R163_165 V163 V165 -123.8874521642742
L163_165 V163 V165 8.040242655663009e-13
C163_165 V163 V165 6.364275363608435e-19

R163_166 V163 V166 24.331578370903262
L163_166 V163 V166 7.095812139093185e-12
C163_166 V163 V166 9.971664370887833e-21

R163_167 V163 V167 -171.03798725041764
L163_167 V163 V167 1.1771636871964099e-12
C163_167 V163 V167 1.1237042437560798e-19

R163_168 V163 V168 -240.93413674844
L163_168 V163 V168 -9.33260149008077e-11
C163_168 V163 V168 -9.583678043382628e-20

R163_169 V163 V169 37.02772300948589
L163_169 V163 V169 3.5240833741214918e-12
C163_169 V163 V169 -2.951975237476088e-20

R163_170 V163 V170 -62.000401350589385
L163_170 V163 V170 5.525529683390213e-12
C163_170 V163 V170 2.232855204419578e-19

R163_171 V163 V171 14.392840450636697
L163_171 V163 V171 5.315669750495219e-13
C163_171 V163 V171 4.134707656757495e-19

R163_172 V163 V172 43.492624786212374
L163_172 V163 V172 1.3812898956428108e-12
C163_172 V163 V172 2.7935225016576757e-19

R163_173 V163 V173 -102.40066390542691
L163_173 V163 V173 -1.078489925740599e-12
C163_173 V163 V173 -3.9001253166340413e-19

R163_174 V163 V174 -37.43872432889669
L163_174 V163 V174 -4.379639403265819e-12
C163_174 V163 V174 -2.2666799406195444e-19

R163_175 V163 V175 -30.04691540654489
L163_175 V163 V175 -6.736829462298175e-13
C163_175 V163 V175 -2.8351873387946757e-19

R163_176 V163 V176 -608.7679491479047
L163_176 V163 V176 -3.8499582468489646e-12
C163_176 V163 V176 1.0471422400002099e-20

R163_177 V163 V177 -61.969130776248214
L163_177 V163 V177 1.0158891753108647e-11
C163_177 V163 V177 1.6302411933574142e-19

R163_178 V163 V178 55.84451378838756
L163_178 V163 V178 -4.123307273538293e-12
C163_178 V163 V178 -1.5885540891516138e-19

R163_179 V163 V179 -48.195760822586834
L163_179 V163 V179 -1.3753742701189343e-12
C163_179 V163 V179 -1.7366874649087558e-19

R163_180 V163 V180 -73.80781031730486
L163_180 V163 V180 -1.4970492202298846e-12
C163_180 V163 V180 -2.836807761297463e-19

R163_181 V163 V181 80.54377337042871
L163_181 V163 V181 9.062359537240423e-12
C163_181 V163 V181 8.75623669355489e-20

R163_182 V163 V182 45.0377162821281
L163_182 V163 V182 1.141343392493918e-12
C163_182 V163 V182 2.4242199644965576e-19

R163_183 V163 V183 41.72316067925528
L163_183 V163 V183 2.0044465296358865e-12
C163_183 V163 V183 -6.020445202482747e-20

R163_184 V163 V184 157.91101032205484
L163_184 V163 V184 5.092437796783562e-12
C163_184 V163 V184 1.0040766894614067e-19

R163_185 V163 V185 97.61690744093708
L163_185 V163 V185 5.753324712442577e-12
C163_185 V163 V185 -1.221545157756911e-19

R163_186 V163 V186 -188.62244496886373
L163_186 V163 V186 2.843909211841261e-12
C163_186 V163 V186 1.4280968200712657e-19

R163_187 V163 V187 -90.43565236056246
L163_187 V163 V187 1.8900254592261346e-11
C163_187 V163 V187 7.010437189568515e-20

R163_188 V163 V188 440.1808795053211
L163_188 V163 V188 1.5889960539161896e-12
C163_188 V163 V188 1.4511408379588754e-19

R163_189 V163 V189 -78.71741943935159
L163_189 V163 V189 -3.8821645980455995e-10
C163_189 V163 V189 2.045933520474337e-19

R163_190 V163 V190 -97.22315251456166
L163_190 V163 V190 -2.411631898309703e-12
C163_190 V163 V190 -2.8190815235366233e-19

R163_191 V163 V191 -62.54925087659268
L163_191 V163 V191 4.109817111714532e-12
C163_191 V163 V191 4.2962797318317034e-19

R163_192 V163 V192 -104.50831464311939
L163_192 V163 V192 -6.753577190245895e-12
C163_192 V163 V192 7.44436808034283e-20

R163_193 V163 V193 -105.824481809484
L163_193 V163 V193 -2.520252259648587e-12
C163_193 V163 V193 -1.6213404384981206e-19

R163_194 V163 V194 163.01000285050853
L163_194 V163 V194 -4.464375236709648e-12
C163_194 V163 V194 -1.8423586310069528e-20

R163_195 V163 V195 34.61985512930963
L163_195 V163 V195 -2.1982992497816797e-12
C163_195 V163 V195 -7.387040636221681e-19

R163_196 V163 V196 1974.126749184574
L163_196 V163 V196 -1.6183895450785355e-12
C163_196 V163 V196 -1.2158257040302915e-19

R163_197 V163 V197 130.97937575691014
L163_197 V163 V197 -4.426146525460383e-12
C163_197 V163 V197 -1.2205323715153628e-19

R163_198 V163 V198 108.08329532750822
L163_198 V163 V198 3.8345743574514994e-12
C163_198 V163 V198 4.018596972858792e-20

R163_199 V163 V199 399.7066215637174
L163_199 V163 V199 -1.9338498699375252e-12
C163_199 V163 V199 -3.110778059514855e-19

R163_200 V163 V200 -473.23777981219087
L163_200 V163 V200 -9.036357715048646e-12
C163_200 V163 V200 -1.5489353420133334e-19

R164_164 V164 0 179.37782006689847
L164_164 V164 0 9.882560790207992e-13
C164_164 V164 0 -1.6054963098215842e-19

R164_165 V164 V165 -78.77476520065322
L164_165 V164 V165 1.767883434959459e-12
C164_165 V164 V165 2.837428983451075e-19

R164_166 V164 V166 17.226707984931004
L164_166 V164 V166 1.0946492663692456e-11
C164_166 V164 V166 4.1617285265447955e-20

R164_167 V164 V167 -88.74075789845664
L164_167 V164 V167 3.8408246147344825e-11
C164_167 V164 V167 -6.183117820588201e-20

R164_168 V164 V168 212.60471710593254
L164_168 V164 V168 2.1884180651260987e-12
C164_168 V164 V168 -5.2091702112316174e-20

R164_169 V164 V169 25.595926571123826
L164_169 V164 V169 1.656339622103232e-12
C164_169 V164 V169 1.41662140853802e-19

R164_170 V164 V170 -40.085790389182236
L164_170 V164 V170 7.351437616948506e-12
C164_170 V164 V170 6.251947971062515e-20

R164_171 V164 V171 32.74739301180536
L164_171 V164 V171 1.3154691580492693e-12
C164_171 V164 V171 1.3977213290629e-19

R164_172 V164 V172 11.312186168013268
L164_172 V164 V172 7.436566110679275e-13
C164_172 V164 V172 2.021072540679344e-19

R164_173 V164 V173 -55.0986828774117
L164_173 V164 V173 -2.0416698021796803e-12
C164_173 V164 V173 -2.2830919846837105e-19

R164_174 V164 V174 -28.711224416947143
L164_174 V164 V174 1.0968196571130706e-11
C164_174 V164 V174 -1.2225449350843161e-20

R164_175 V164 V175 334.0853842474759
L164_175 V164 V175 6.661600930428674e-11
C164_175 V164 V175 1.3039817362087686e-20

R164_176 V164 V176 -25.214836146523933
L164_176 V164 V176 -9.280265740582372e-13
C164_176 V164 V176 -2.6112204885086006e-19

R164_177 V164 V177 -38.32909306810373
L164_177 V164 V177 -4.089468994662554e-12
C164_177 V164 V177 2.100596261128192e-20

R164_178 V164 V178 42.83488917927384
L164_178 V164 V178 -3.3472857891118018e-12
C164_178 V164 V178 -6.792301174518812e-20

R164_179 V164 V179 -107.93408174174716
L164_179 V164 V179 -1.8244494680291358e-12
C164_179 V164 V179 -6.281099299651779e-20

R164_180 V164 V180 -24.466604050714782
L164_180 V164 V180 -1.826417338545224e-12
C164_180 V164 V180 1.4111467478238856e-19

R164_181 V164 V181 39.150748356084236
L164_181 V164 V181 5.731875813985341e-12
C164_181 V164 V181 2.2566974524123115e-20

R164_182 V164 V182 24.802476708231175
L164_182 V164 V182 1.4593574311162596e-12
C164_182 V164 V182 1.0163337448554434e-19

R164_183 V164 V183 334.02597757492373
L164_183 V164 V183 -1.521306380531783e-11
C164_183 V164 V183 4.8460545819419114e-20

R164_184 V164 V184 24.635642011080193
L164_184 V164 V184 2.132933964065093e-12
C164_184 V164 V184 -2.627512380290344e-20

R164_185 V164 V185 77.18627400173206
L164_185 V164 V185 7.048622884872001e-12
C164_185 V164 V185 -1.349012576271816e-21

R164_186 V164 V186 321.4691488601252
L164_186 V164 V186 6.12323095853898e-12
C164_186 V164 V186 6.002643778240464e-21

R164_187 V164 V187 151.39808272114396
L164_187 V164 V187 3.161508011824996e-12
C164_187 V164 V187 -4.234414824498947e-21

R164_188 V164 V188 -51.722586416561875
L164_188 V164 V188 -4.846784658237762e-12
C164_188 V164 V188 -8.70705919485766e-20

R164_189 V164 V189 -60.31932292079983
L164_189 V164 V189 8.745537314207978e-12
C164_189 V164 V189 1.0179129194086274e-19

R164_190 V164 V190 -43.531168072029786
L164_190 V164 V190 -4.0662924935044e-12
C164_190 V164 V190 -1.0117810790445453e-19

R164_191 V164 V191 -88.80858471018207
L164_191 V164 V191 5.308646279559622e-12
C164_191 V164 V191 9.502631644252267e-22

R164_192 V164 V192 -124.51313428421273
L164_192 V164 V192 1.141112331674625e-11
C164_192 V164 V192 2.533709787703827e-19

R164_193 V164 V193 -121.87061444532522
L164_193 V164 V193 -5.385405611061718e-12
C164_193 V164 V193 -8.407372129420437e-21

R164_194 V164 V194 162.88273570037293
L164_194 V164 V194 4.612387041501667e-12
C164_194 V164 V194 1.8856686417124785e-19

R164_195 V164 V195 198.68893969156767
L164_195 V164 V195 -2.836177129967431e-12
C164_195 V164 V195 8.101612241856044e-20

R164_196 V164 V196 60.857202214987595
L164_196 V164 V196 -3.2674336283697517e-12
C164_196 V164 V196 -4.943764789262715e-19

R164_197 V164 V197 67.46641845543085
L164_197 V164 V197 -3.309187932781959e-12
C164_197 V164 V197 -1.674365205560977e-19

R164_198 V164 V198 93.63010784220963
L164_198 V164 V198 1.1628543626784298e-11
C164_198 V164 V198 2.6893155203098138e-20

R164_199 V164 V199 -67.05920006522172
L164_199 V164 V199 -3.7654145924275424e-12
C164_199 V164 V199 -1.61427690330639e-19

R164_200 V164 V200 161.26731118269575
L164_200 V164 V200 -4.645603999783842e-12
C164_200 V164 V200 5.532079918795181e-20

R165_165 V165 0 61.462835451905626
L165_165 V165 0 4.777505031889042e-13
C165_165 V165 0 -2.0592298447483364e-18

R165_166 V165 V166 156.7671287738101
L165_166 V165 V166 -1.7974159459699394e-12
C165_166 V165 V166 2.4791266137927986e-20

R165_167 V165 V167 125.06530986236517
L165_167 V165 V167 -4.0765228858961115e-12
C165_167 V165 V167 1.9782208906698523e-21

R165_168 V165 V168 277.27415117697734
L165_168 V165 V168 -2.0220910174825932e-11
C165_168 V165 V168 2.001056485459447e-19

R165_169 V165 V169 131.29234235771577
L165_169 V165 V169 7.702459277077309e-13
C165_169 V165 V169 2.9525324100336515e-19

R165_170 V165 V170 67.73954447248171
L165_170 V165 V170 -5.963054424723308e-12
C165_170 V165 V170 -6.0728303596819565e-19

R165_171 V165 V171 140.2937469636722
L165_171 V165 V171 -4.734767291593563e-13
C165_171 V165 V171 -9.529418190901048e-19

R165_172 V165 V172 93.7527082848155
L165_172 V165 V172 -7.491381069841558e-13
C165_172 V165 V172 -6.008072099043564e-19

R165_173 V165 V173 53.745654001904256
L165_173 V165 V173 3.6622327805993274e-13
C165_173 V165 V173 7.347976314303014e-19

R165_174 V165 V174 -79.7895289917297
L165_174 V165 V174 1.129423546350811e-12
C165_174 V165 V174 5.370597532333336e-19

R165_175 V165 V175 -117.32250637521823
L165_175 V165 V175 1.5397594005886038e-12
C165_175 V165 V175 1.9351463169821843e-19

R165_176 V165 V176 -204.0440038666392
L165_176 V165 V176 7.746661845173269e-13
C165_176 V165 V176 2.264470365969616e-19

R165_177 V165 V177 -74.83728800332578
L165_177 V165 V177 -8.253802044730307e-13
C165_177 V165 V177 -2.460402260144385e-19

R165_178 V165 V178 -202.041905716922
L165_178 V165 V178 1.942329471851846e-12
C165_178 V165 V178 4.053079729431654e-19

R165_179 V165 V179 -555.6589762939495
L165_179 V165 V179 7.032883518826862e-13
C165_179 V165 V179 6.963421642635907e-19

R165_180 V165 V180 -119.90178661681183
L165_180 V165 V180 1.0942388317806635e-12
C165_180 V165 V180 4.814307836905831e-19

R165_181 V165 V181 -517.90611309748
L165_181 V165 V181 -6.677430354773936e-12
C165_181 V165 V181 -2.5413985487358184e-19

R165_182 V165 V182 109.69558966859383
L165_182 V165 V182 -4.680471452146756e-13
C165_182 V165 V182 -6.241664008836811e-19

R165_183 V165 V183 141.71175147679818
L165_183 V165 V183 3.0924200356213358e-12
C165_183 V165 V183 3.957036350419966e-20

R165_184 V165 V184 117.03161514283354
L165_184 V165 V184 -1.7196121805564872e-12
C165_184 V165 V184 -1.2856550330372236e-19

R165_185 V165 V185 63.811091544783075
L165_185 V165 V185 -7.98935182199633e-12
C165_185 V165 V185 1.7901174188147188e-19

R165_186 V165 V186 -297.0985822276638
L165_186 V165 V186 -8.173903429511689e-13
C165_186 V165 V186 -1.4190914114890787e-19

R165_187 V165 V187 -217.23169057661494
L165_187 V165 V187 -5.811942742270015e-13
C165_187 V165 V187 -4.066355871539487e-19

R165_188 V165 V188 2472.5939363825114
L165_188 V165 V188 -7.510373724179383e-13
C165_188 V165 V188 -3.8672166831040057e-19

R165_189 V165 V189 -147.58200856187207
L165_189 V165 V189 5.326084012408907e-11
C165_189 V165 V189 -3.3020991331360717e-19

R165_190 V165 V190 -93.71422162640927
L165_190 V165 V190 8.987598202924763e-13
C165_190 V165 V190 5.817263480666921e-19

R165_191 V165 V191 -185.900527956481
L165_191 V165 V191 -9.625382029380947e-13
C165_191 V165 V191 -4.859629371409446e-19

R165_192 V165 V192 -195.05015160594985
L165_192 V165 V192 -1.0531831328135056e-11
C165_192 V165 V192 -2.6115159766627593e-19

R165_193 V165 V193 -84.03314153768773
L165_193 V165 V193 2.0398182272236233e-12
C165_193 V165 V193 3.077658319837417e-19

R165_194 V165 V194 84.70586079859555
L165_194 V165 V194 8.598041710419463e-13
C165_194 V165 V194 -4.6703735270749895e-20

R165_195 V165 V195 109.77966408372653
L165_195 V165 V195 4.86613531042732e-13
C165_195 V165 V195 8.661053024485818e-19

R165_196 V165 V196 173.9335787695916
L165_196 V165 V196 3.6910345060590887e-13
C165_196 V165 V196 9.70217554917375e-19

R165_197 V165 V197 78.44003078959824
L165_197 V165 V197 9.120851584625323e-13
C165_197 V165 V197 3.9289987352414646e-19

R165_198 V165 V198 850.725615817544
L165_198 V165 V198 -1.2517526464027825e-12
C165_198 V165 V198 -1.5455075970712714e-19

R165_199 V165 V199 -337.4252040667874
L165_199 V165 V199 1.1122795241063688e-12
C165_199 V165 V199 4.7814616486419645e-19

R165_200 V165 V200 288.2982381794561
L165_200 V165 V200 -2.8806614048263545e-12
C165_200 V165 V200 8.404475229092301e-20

R166_166 V166 0 -36.31654088289189
L166_166 V166 0 5.145808456709142e-13
C166_166 V166 0 1.3560052201948234e-18

R166_167 V166 V167 11.065464204117093
L166_167 V166 V167 2.6633478966361302e-12
C166_167 V166 V167 -7.949206396558743e-20

R166_168 V166 V168 8.757715570134526
L166_168 V166 V168 1.6559110337498785e-12
C166_168 V166 V168 -1.5841741970342013e-19

R166_169 V166 V169 -13.417727504629203
L166_169 V166 V169 5.977124071308967e-12
C166_169 V166 V169 1.5259193388087815e-19

R166_170 V166 V170 8.139393586394444
L166_170 V166 V170 8.144356428023476e-13
C166_170 V166 V170 1.2496099157915342e-19

R166_171 V166 V171 -14.804393164807957
L166_171 V166 V171 -3.1452848182039762e-12
C166_171 V166 V171 -2.576759405843694e-21

R166_172 V166 V172 -12.210513300893139
L166_172 V166 V172 -1.7463767621494966e-12
C166_172 V166 V172 7.401197806584328e-20

R166_173 V166 V173 17.742620198718917
L166_173 V166 V173 1.6872722829648392e-12
C166_173 V166 V173 2.0058587359626256e-20

R166_174 V166 V174 4.3072119306380445
L166_174 V166 V174 5.193858033361092e-13
C166_174 V166 V174 1.1419250298342737e-19

R166_175 V166 V175 -20.466775601937325
L166_175 V166 V175 -1.961271616543607e-11
C166_175 V166 V175 1.7588438737428491e-19

R166_176 V166 V176 -13.959060385112474
L166_176 V166 V176 4.504247990826248e-12
C166_176 V166 V176 2.973877098034011e-19

R166_177 V166 V177 33.07774618269337
L166_177 V166 V177 -2.876470874901893e-12
C166_177 V166 V177 -1.5825305555580902e-19

R166_178 V166 V178 -6.785143468743655
L166_178 V166 V178 -7.572988562517714e-13
C166_178 V166 V178 -7.867201813556984e-20

R166_179 V166 V179 19.41177199659228
L166_179 V166 V179 6.5513459067178246e-12
C166_179 V166 V179 -1.275698804198809e-19

R166_180 V166 V180 11.628576567331388
L166_180 V166 V180 1.0306787009596164e-11
C166_180 V166 V180 -2.502498419655495e-19

R166_181 V166 V181 -22.55683702177934
L166_181 V166 V181 4.863110086736269e-11
C166_181 V166 V181 -1.0404235918757684e-19

R166_182 V166 V182 -9.151778541378569
L166_182 V166 V182 -1.9459023078949346e-12
C166_182 V166 V182 1.3793615145221915e-20

R166_183 V166 V183 198.4871898303055
L166_183 V166 V183 -8.64551228846158e-12
C166_183 V166 V183 -1.1372955739780758e-20

R166_184 V166 V184 -3533.6506943603285
L166_184 V166 V184 -3.104174925473416e-12
C166_184 V166 V184 3.3155808825468645e-20

R166_185 V166 V185 -276.2446979315839
L166_185 V166 V185 -6.59873765720018e-12
C166_185 V166 V185 1.7919450014661572e-19

R166_186 V166 V186 20.16722666352232
L166_186 V166 V186 -1.3171671166605371e-11
C166_186 V166 V186 -7.98456026605342e-20

R166_187 V166 V187 -143.31472090618558
L166_187 V166 V187 -4.6296307260066606e-12
C166_187 V166 V187 9.180442987532286e-20

R166_188 V166 V188 -54.36908153399054
L166_188 V166 V188 1.0601579795830897e-11
C166_188 V166 V188 2.5490154964080886e-20

R166_189 V166 V189 82.28406997023902
L166_189 V166 V189 1.3737355009833172e-11
C166_189 V166 V189 -1.9200748458689478e-20

R166_190 V166 V190 19.778277512280518
L166_190 V166 V190 1.7391041908590748e-12
C166_190 V166 V190 -5.704307303353175e-20

R166_191 V166 V191 -854.6825392479992
L166_191 V166 V191 6.9192429280059755e-12
C166_191 V166 V191 -6.109975994285923e-20

R166_192 V166 V192 -560.0621355652373
L166_192 V166 V192 4.660039105744713e-11
C166_192 V166 V192 -5.1530957025151784e-20

R166_193 V166 V193 149.2934005613115
L166_193 V166 V193 4.088890235619944e-12
C166_193 V166 V193 2.897166363008292e-20

R166_194 V166 V194 -102.05406522491955
L166_194 V166 V194 2.6192305094925476e-12
C166_194 V166 V194 5.512172530886453e-20

R166_195 V166 V195 -122.98577344332814
L166_195 V166 V195 -5.6831138604477825e-12
C166_195 V166 V195 -5.666606749771816e-20

R166_196 V166 V196 466.71131009131784
L166_196 V166 V196 2.778683400618384e-12
C166_196 V166 V196 2.2351024409176655e-19

R166_197 V166 V197 -458.32976313917453
L166_197 V166 V197 -1.6070933640037786e-11
C166_197 V166 V197 -1.0505620973873647e-19

R166_198 V166 V198 -13.088948801074158
L166_198 V166 V198 -1.5541392583700484e-12
C166_198 V166 V198 -4.888095949828285e-20

R166_199 V166 V199 -333.4186427266251
L166_199 V166 V199 2.3624294201145227e-11
C166_199 V166 V199 6.088261162794354e-20

R166_200 V166 V200 41.61231692206425
L166_200 V166 V200 -4.149716091452776e-12
C166_200 V166 V200 -6.514549926288986e-20

R167_167 V167 0 114.75550538930052
L167_167 V167 0 3.908211397903762e-13
C167_167 V167 0 4.227136042119792e-19

R167_168 V167 V168 85.70729631792071
L167_168 V167 V168 3.5642199194130762e-12
C167_168 V167 V168 -1.6507557779773967e-19

R167_169 V167 V169 74.15022620870849
L167_169 V167 V169 1.776678948896107e-12
C167_169 V167 V169 2.307997027218012e-19

R167_170 V167 V170 -44.064828830864705
L167_170 V167 V170 1.9998979936072773e-11
C167_170 V167 V170 4.680190273387491e-21

R167_171 V167 V171 16.994048516689297
L167_171 V167 V171 1.760795427715575e-12
C167_171 V167 V171 1.2801187529332505e-19

R167_172 V167 V172 71.0908596804923
L167_172 V167 V172 -4.554710202269859e-11
C167_172 V167 V172 1.2137683449861257e-19

R167_173 V167 V173 -54.20704747417815
L167_173 V167 V173 -1.0856834157227177e-11
C167_173 V167 V173 3.765217562209225e-20

R167_174 V167 V174 -12.088573571072994
L167_174 V167 V174 -3.724512611016623e-12
C167_174 V167 V174 1.3870918885233608e-19

R167_175 V167 V175 15.844240783524777
L167_175 V167 V175 5.582644988335705e-13
C167_175 V167 V175 9.780588035992149e-20

R167_176 V167 V176 1036.021980406485
L167_176 V167 V176 4.1228202188768526e-12
C167_176 V167 V176 9.923231868435793e-20

R167_177 V167 V177 -95.63410688970374
L167_177 V167 V177 -4.26230728463977e-12
C167_177 V167 V177 -1.1067320507216101e-19

R167_178 V167 V178 27.53615705444376
L167_178 V167 V178 8.192857246598702e-12
C167_178 V167 V178 -1.962798810081218e-20

R167_179 V167 V179 -24.721903034419473
L167_179 V167 V179 -1.1173564400576313e-12
C167_179 V167 V179 2.1142969614874736e-20

R167_180 V167 V180 -47.03175873036028
L167_180 V167 V180 -3.5358474322565734e-12
C167_180 V167 V180 -2.6318616100368873e-20

R167_181 V167 V181 70.58121347767204
L167_181 V167 V181 -3.639715127194999e-11
C167_181 V167 V181 -2.292534540412982e-19

R167_182 V167 V182 22.333009756004515
L167_182 V167 V182 4.6406023338005676e-12
C167_182 V167 V182 -1.8963404981856825e-20

R167_183 V167 V183 -43.058275787984584
L167_183 V167 V183 -2.843440674794234e-12
C167_183 V167 V183 -2.9822283800233636e-21

R167_184 V167 V184 199.0912297793169
L167_184 V167 V184 -1.1844874456034227e-11
C167_184 V167 V184 -1.850357045942658e-20

R167_185 V167 V185 490.96512608735253
L167_185 V167 V185 -3.0487266921544255e-12
C167_185 V167 V185 1.906130837997022e-19

R167_186 V167 V186 -74.48742920734249
L167_186 V167 V186 -3.4036738472400218e-12
C167_186 V167 V186 -1.1611004894947628e-19

R167_187 V167 V187 57.243419103806794
L167_187 V167 V187 1.576495800257756e-11
C167_187 V167 V187 -8.145976899238677e-20

R167_188 V167 V188 127.32682003606233
L167_188 V167 V188 -2.4747193422602166e-12
C167_188 V167 V188 -9.03938120672083e-20

R167_189 V167 V189 -192.13941875185753
L167_189 V167 V189 1.862578887919604e-12
C167_189 V167 V189 1.3148637005698831e-19

R167_190 V167 V190 -40.443995704677214
L167_190 V167 V190 -1.7679250950537638e-11
C167_190 V167 V190 -2.3280362684788e-20

R167_191 V167 V191 66.11105985287082
L167_191 V167 V191 4.164304617567285e-12
C167_191 V167 V191 1.4321913039310358e-20

R167_192 V167 V192 -228.95533080579577
L167_192 V167 V192 3.5023108789583278e-12
C167_192 V167 V192 1.9442278400560306e-19

R167_193 V167 V193 -344.98218717668186
L167_193 V167 V193 5.973869167051961e-12
C167_193 V167 V193 3.718389664367478e-20

R167_194 V167 V194 321.8020566900152
L167_194 V167 V194 1.5829450911983979e-12
C167_194 V167 V194 2.436808553634391e-19

R167_195 V167 V195 -115.27475454666784
L167_195 V167 V195 -2.4005153329469015e-12
C167_195 V167 V195 -1.8017001278787152e-20

R167_196 V167 V196 -191.50902485533095
L167_196 V167 V196 5.811476708554092e-12
C167_196 V167 V196 -1.750694430703869e-19

R167_197 V167 V197 696.8668142251931
L167_197 V167 V197 -2.3916739625011236e-12
C167_197 V167 V197 -2.3654428482063695e-19

R167_198 V167 V198 37.50685601395977
L167_198 V167 V198 2.912237709276456e-11
C167_198 V167 V198 -2.9831324355788026e-20

R167_199 V167 V199 -73.89821012253235
L167_199 V167 V199 -4.680405637716198e-12
C167_199 V167 V199 5.893063558420538e-20

R167_200 V167 V200 -1143.6986347611864
L167_200 V167 V200 -2.209494978415975e-12
C167_200 V167 V200 -5.803146109375534e-20

R168_168 V168 0 22.242280422733604
L168_168 V168 0 3.7516528053983814e-13
C168_168 V168 0 1.2268367464502943e-18

R168_169 V168 V169 52.01960991792592
L168_169 V168 V169 1.482248089706898e-12
C168_169 V168 V169 3.044261885463744e-19

R168_170 V168 V170 -27.97415346292234
L168_170 V168 V170 -3.727692557539723e-12
C168_170 V168 V170 9.746014050724114e-20

R168_171 V168 V171 832.3026810363219
L168_171 V168 V171 -2.9756114183966286e-12
C168_171 V168 V171 1.6767404603248487e-19

R168_172 V168 V172 20.888762590899997
L168_172 V168 V172 7.491422202006115e-13
C168_172 V168 V172 2.4365645739175446e-19

R168_173 V168 V173 -52.43473764662516
L168_173 V168 V173 -2.730922909804827e-12
C168_173 V168 V173 -2.5620566500707225e-20

R168_174 V168 V174 -9.657168848363584
L168_174 V168 V174 -4.41059782384945e-12
C168_174 V168 V174 1.341383040349811e-19

R168_175 V168 V175 -260.4169260644381
L168_175 V168 V175 8.039927669878912e-12
C168_175 V168 V175 1.6037210298954816e-19

R168_176 V168 V176 11.477328996876718
L168_176 V168 V176 7.462822641416897e-13
C168_176 V168 V176 2.537927456395132e-19

R168_177 V168 V177 -128.69238241027907
L168_177 V168 V177 -1.1332396499149568e-11
C168_177 V168 V177 -1.0459612215839696e-19

R168_178 V168 V178 17.02531154782852
L168_178 V168 V178 2.407901710312922e-12
C168_178 V168 V178 -1.2123988221722637e-19

R168_179 V168 V179 -222.77916037910734
L168_179 V168 V179 8.524113851881157e-12
C168_179 V168 V179 -1.9995368828620926e-19

R168_180 V168 V180 -19.285805852002785
L168_180 V168 V180 -1.1197493068582653e-12
C168_180 V168 V180 -2.36990909032147e-19

R168_181 V168 V181 83.81265344126018
L168_181 V168 V181 -6.518059296992094e-12
C168_181 V168 V181 -3.3711479161278743e-19

R168_182 V168 V182 24.172329814224124
L168_182 V168 V182 6.034360142288173e-12
C168_182 V168 V182 9.033538964223169e-20

R168_183 V168 V183 131.9688802489372
L168_183 V168 V183 4.913283317776582e-12
C168_183 V168 V183 -3.708821063116773e-20

R168_184 V168 V184 -58.79526738025157
L168_184 V168 V184 -1.0665223499397006e-11
C168_184 V168 V184 -2.552886384753798e-20

R168_185 V168 V185 353.8776751200405
L168_185 V168 V185 -3.5316130665507934e-12
C168_185 V168 V185 2.6874112820359886e-19

R168_186 V168 V186 -43.50324962961002
L168_186 V168 V186 -5.48652426377828e-12
C168_186 V168 V186 -1.4541625413156517e-19

R168_187 V168 V187 -157.26262359053422
L168_187 V168 V187 -2.8830456974928982e-12
C168_187 V168 V187 5.149263873606319e-20

R168_188 V168 V188 86.46918202105648
L168_188 V168 V188 -1.2662491552284902e-12
C168_188 V168 V188 -1.7958242233267745e-20

R168_189 V168 V189 -193.85607740730003
L168_189 V168 V189 1.3607600993192435e-12
C168_189 V168 V189 2.5646810775187486e-19

R168_190 V168 V190 -42.48051466370829
L168_190 V168 V190 -9.769357167482518e-12
C168_190 V168 V190 -1.2372688054601915e-19

R168_191 V168 V191 -123.08243970822885
L168_191 V168 V191 -2.0845395764379045e-12
C168_191 V168 V191 1.9234668046390582e-19

R168_192 V168 V192 58.13671702345755
L168_192 V168 V192 9.106088928558091e-13
C168_192 V168 V192 3.045582583481702e-19

R168_193 V168 V193 -206.45638402113414
L168_193 V168 V193 1.663027633486281e-11
C168_193 V168 V193 -3.1984019917823066e-20

R168_194 V168 V194 119.00082232040062
L168_194 V168 V194 1.0714502040468817e-12
C168_194 V168 V194 2.7011450408609675e-19

R168_195 V168 V195 100.41151230955974
L168_195 V168 V195 1.6325882667070432e-12
C168_195 V168 V195 -3.1779230212953406e-19

R168_196 V168 V196 -182.9761223953278
L168_196 V168 V196 -1.307842162989849e-12
C168_196 V168 V196 -2.153913454820727e-19

R168_197 V168 V197 143.972992704327
L168_197 V168 V197 -1.9551800744951797e-12
C168_197 V168 V197 -3.5842301205698556e-19

R168_198 V168 V198 33.027100483811836
L168_198 V168 V198 -1.3431729073487574e-10
C168_198 V168 V198 1.0825424344040792e-20

R168_199 V168 V199 152.35625414701303
L168_199 V168 V199 -3.946149591842169e-12
C168_199 V168 V199 -2.0359542098002265e-20

R168_200 V168 V200 -38.64518835623582
L168_200 V168 V200 -1.949519745235799e-12
C168_200 V168 V200 -2.0972337190354273e-19

R169_169 V169 0 77.5573577250853
L169_169 V169 0 -5.005682747171857e-13
C169_169 V169 0 8.367393810901685e-19

R169_170 V169 V170 65.28087025200541
L169_170 V169 V170 -3.5146403292648805e-12
C169_170 V169 V170 6.158927851249398e-21

R169_171 V169 V171 -39.14165577489911
L169_171 V169 V171 -4.592832867060805e-12
C169_171 V169 V171 2.1482072764847656e-20

R169_172 V169 V172 -33.82447431538867
L169_172 V169 V172 -1.4637528829320846e-12
C169_172 V169 V172 -1.8360160884673142e-19

R169_173 V169 V173 43.26636615580904
L169_173 V169 V173 2.4894236154601807e-12
C169_173 V169 V173 2.026143819802992e-19

R169_174 V169 V174 17.064457970691205
L169_174 V169 V174 -1.5840993345028162e-12
C169_174 V169 V174 -4.664183256344766e-19

R169_175 V169 V175 -149.7410031016585
L169_175 V169 V175 -2.182709238902033e-12
C169_175 V169 V175 -8.559323789312496e-20

R169_176 V169 V176 -161.9430294636458
L169_176 V169 V176 -1.7053039306170096e-12
C169_176 V169 V176 -8.542820754596166e-20

R169_177 V169 V177 46.39482770302605
L169_177 V169 V177 1.3367599721526333e-12
C169_177 V169 V177 2.300059045145962e-19

R169_178 V169 V178 -45.95477694487345
L169_178 V169 V178 3.0055456086255908e-12
C169_178 V169 V178 1.0905131197099184e-19

R169_179 V169 V179 60.275041617314216
L169_179 V169 V179 1.1129979729651187e-11
C169_179 V169 V179 -1.5283216161003135e-19

R169_180 V169 V180 52.49022159885642
L169_180 V169 V180 2.4995214167290896e-12
C169_180 V169 V180 -5.163545978111686e-20

R169_181 V169 V181 -51.26117961254343
L169_181 V169 V181 -7.455107365222256e-12
C169_181 V169 V181 3.0971973355474773e-19

R169_182 V169 V182 -23.934351516505068
L169_182 V169 V182 4.363562457235154e-12
C169_182 V169 V182 1.2720648550742203e-19

R169_183 V169 V183 -966.5626588415221
L169_183 V169 V183 -5.465537507383492e-12
C169_183 V169 V183 -9.621900433878562e-20

R169_184 V169 V184 -1180.6177371887254
L169_184 V169 V184 -6.640737679209494e-11
C169_184 V169 V184 5.254310778758893e-20

R169_185 V169 V185 -71.03582435496824
L169_185 V169 V185 3.740576351994995e-12
C169_185 V169 V185 -2.0314895616790654e-19

R169_186 V169 V186 148.61399358274636
L169_186 V169 V186 5.243003597727135e-11
C169_186 V169 V186 1.0289485679072529e-19

R169_187 V169 V187 -2448.2210101526334
L169_187 V169 V187 1.840950450497444e-12
C169_187 V169 V187 3.5463089473283735e-19

R169_188 V169 V188 3836.3293884278473
L169_188 V169 V188 1.2464880827738119e-12
C169_188 V169 V188 3.3992401265625975e-19

R169_189 V169 V189 84.7499931168639
L169_189 V169 V189 -1.0407899260019706e-12
C169_189 V169 V189 -1.7388124258181648e-19

R169_190 V169 V190 47.260028986839636
L169_190 V169 V190 1.0581546686402335e-11
C169_190 V169 V190 -4.1960619888898674e-20

R169_191 V169 V191 -343.63584354701607
L169_191 V169 V191 7.429506275080132e-12
C169_191 V169 V191 -1.393481376339829e-20

R169_192 V169 V192 -359.10697508518075
L169_192 V169 V192 -1.6388457698985409e-12
C169_192 V169 V192 -3.8955000544781735e-19

R169_193 V169 V193 68.74422962387152
L169_193 V169 V193 3.362624238566091e-12
C169_193 V169 V193 -1.8930185157490203e-19

R169_194 V169 V194 -73.17912303265967
L169_194 V169 V194 -7.341238945740934e-13
C169_194 V169 V194 -6.585897391724421e-19

R169_195 V169 V195 -335.3409270874967
L169_195 V169 V195 -2.5814604634078994e-12
C169_195 V169 V195 -1.4012493901609763e-19

R169_196 V169 V196 -436.1931300335891
L169_196 V169 V196 -2.374351779411649e-12
C169_196 V169 V196 7.515701704448662e-20

R169_197 V169 V197 -91.82596634037861
L169_197 V169 V197 7.940456831603147e-12
C169_197 V169 V197 2.393871613507167e-19

R169_198 V169 V198 -43.18874819464656
L169_198 V169 V198 4.735032322326126e-12
C169_198 V169 V198 3.1204756504886387e-20

R169_199 V169 V199 294.607049958054
L169_199 V169 V199 7.451841176156324e-12
C169_199 V169 V199 -1.686135778919414e-19

R169_200 V169 V200 69.87542903584952
L169_200 V169 V200 1.497061975455701e-12
C169_200 V169 V200 2.4155073261827454e-19

R170_170 V170 0 35.86453347745478
L170_170 V170 0 8.680414529417709e-13
C170_170 V170 0 -1.0241070906153007e-18

R170_171 V170 V171 50.857932649835874
L170_171 V170 V171 -1.9100910157786945e-12
C170_171 V170 V171 -4.0790581384714256e-19

R170_172 V170 V172 35.60289301269799
L170_172 V170 V172 -1.4358433066392923e-11
C170_172 V170 V172 -2.5819136479020194e-19

R170_173 V170 V173 -31.30383574816453
L170_173 V170 V173 8.481917678240197e-11
C170_173 V170 V173 3.757832845576465e-19

R170_174 V170 V174 -18.68098946220735
L170_174 V170 V174 2.2562216457607082e-12
C170_174 V170 V174 2.5029092700949804e-19

R170_175 V170 V175 85.20075810920518
L170_175 V170 V175 2.7416817289379826e-12
C170_175 V170 V175 5.704874953991821e-20

R170_176 V170 V176 44.90822449064374
L170_176 V170 V176 1.1039528998839132e-11
C170_176 V170 V176 2.4517714121651078e-20

R170_177 V170 V177 -454.4648177975961
L170_177 V170 V177 4.4900925740901124e-12
C170_177 V170 V177 -9.483463682870483e-20

R170_178 V170 V178 10.08011697014394
L170_178 V170 V178 7.459267200611874e-13
C170_178 V170 V178 1.9007351819650017e-19

R170_179 V170 V179 -55.98233263275314
L170_179 V170 V179 -6.284411652429788e-10
C170_179 V170 V179 3.254110432531509e-19

R170_180 V170 V180 -30.453711921457725
L170_180 V170 V180 2.0895669120995764e-11
C170_180 V170 V180 2.8143190737550284e-19

R170_181 V170 V181 57.55873116798738
L170_181 V170 V181 -3.997958274853677e-12
C170_181 V170 V181 -1.0861441001270581e-19

R170_182 V170 V182 339.45396669961656
L170_182 V170 V182 -1.0063518708745646e-12
C170_182 V170 V182 -2.176062125660413e-19

R170_183 V170 V183 415.94063507502204
L170_183 V170 V183 3.168273128060196e-11
C170_183 V170 V183 4.3672648086131955e-21

R170_184 V170 V184 216.31183232906315
L170_184 V170 V184 -1.1088462303677678e-08
C170_184 V170 V184 -9.748411269823067e-20

R170_185 V170 V185 -96.79503823001204
L170_185 V170 V185 -7.623876704783202e-12
C170_185 V170 V185 7.170534306190811e-20

R170_186 V170 V186 -36.16844428520263
L170_186 V170 V186 6.185293694144896e-12
C170_186 V170 V186 -1.1245220327047038e-20

R170_187 V170 V187 142.45947925057752
L170_187 V170 V187 3.3988098215997077e-12
C170_187 V170 V187 -2.348867763924531e-19

R170_188 V170 V188 153.5477943658219
L170_188 V170 V188 -8.062095510003083e-12
C170_188 V170 V188 -2.0370678044434184e-19

R170_189 V170 V189 145.1923742031899
L170_189 V170 V189 2.90155371211637e-12
C170_189 V170 V189 -1.1421109317368255e-19

R170_190 V170 V190 53.0653045826826
L170_190 V170 V190 4.25020292911879e-12
C170_190 V170 V190 2.1468983785650104e-19

R170_191 V170 V191 -707.8834967531935
L170_191 V170 V191 -2.5976539137677898e-12
C170_191 V170 V191 -1.5345118153675906e-19

R170_192 V170 V192 -4893.798083878475
L170_192 V170 V192 6.477541465401414e-12
C170_192 V170 V192 -3.5389952565659426e-20

R170_193 V170 V193 321.91046391636735
L170_193 V170 V193 -1.6922803579978295e-11
C170_193 V170 V193 1.1435212005722424e-19

R170_194 V170 V194 -53.493876867058134
L170_194 V170 V194 -4.994893183327811e-12
C170_194 V170 V194 2.7487573906620014e-20

R170_195 V170 V195 331.2497304213388
L170_195 V170 V195 2.2660886372052088e-12
C170_195 V170 V195 3.6470814002341206e-19

R170_196 V170 V196 981.7072524787303
L170_196 V170 V196 -2.6741670277204154e-11
C170_196 V170 V196 2.9771961716841284e-19

R170_197 V170 V197 -56.22831347167092
L170_197 V170 V197 -3.2253211202466697e-12
C170_197 V170 V197 1.0693417900834238e-19

R170_198 V170 V198 127.71232304552689
L170_198 V170 V198 -1.1992328782805176e-11
C170_198 V170 V198 -1.0554948463401939e-19

R170_199 V170 V199 -24952.653373672238
L170_199 V170 V199 -7.41789696255326e-11
C170_199 V170 V199 1.3195143021061176e-19

R170_200 V170 V200 -94.09563885896348
L170_200 V170 V200 -1.1488576547316185e-10
C170_200 V170 V200 7.450235119726804e-21

R171_171 V171 0 796.884161560911
L171_171 V171 0 -8.282541960147861e-13
C171_171 V171 0 -1.4376525349695837e-18

R171_172 V171 V172 -39.930824053216554
L171_172 V171 V172 -1.0614509213465747e-12
C171_172 V171 V172 -4.538899286654417e-19

R171_173 V171 V173 99.47859761603011
L171_173 V171 V173 7.232256548271097e-13
C171_173 V171 V173 5.378804588647966e-19

R171_174 V171 V174 18.1972685294336
L171_174 V171 V174 1.3527249469935456e-12
C171_174 V171 V174 4.204213887733607e-19

R171_175 V171 V175 73.66838589601959
L171_175 V171 V175 1.1089012350276585e-12
C171_175 V171 V175 2.817733084832072e-19

R171_176 V171 V176 -346.21600873406777
L171_176 V171 V176 4.666952418762687e-12
C171_176 V171 V176 8.513049317399898e-20

R171_177 V171 V177 46.929923348537294
L171_177 V171 V177 -5.997390436077575e-12
C171_177 V171 V177 -2.6450674125953923e-19

R171_178 V171 V178 -35.086869459755704
L171_178 V171 V178 2.155939412773634e-12
C171_178 V171 V178 2.310560103526587e-19

R171_179 V171 V179 25.053625267335345
L171_179 V171 V179 5.488487627175062e-13
C171_179 V171 V179 4.011716426736687e-19

R171_180 V171 V180 53.305899336905355
L171_180 V171 V180 8.46819311270055e-13
C171_180 V171 V180 3.883463696787138e-19

R171_181 V171 V181 -62.6173993009307
L171_181 V171 V181 -2.662301585709436e-12
C171_181 V171 V181 -3.5136386967932384e-21

R171_182 V171 V182 -26.65976161902116
L171_182 V171 V182 -5.936242530598634e-13
C171_182 V171 V182 -4.0790497529287493e-19

R171_183 V171 V183 -50.765980942467024
L171_183 V171 V183 -3.695750169276546e-12
C171_183 V171 V183 8.723079026128426e-20

R171_184 V171 V184 -287.93123549431436
L171_184 V171 V184 -4.995419495602574e-12
C171_184 V171 V184 -1.0106564299920198e-19

R171_185 V171 V185 -81.93557881203499
L171_185 V171 V185 -1.7075030491670577e-11
C171_185 V171 V185 1.4433516101164688e-19

R171_186 V171 V186 87.35683196167138
L171_186 V171 V186 -2.4889825086385424e-12
C171_186 V171 V186 -1.0329015728095167e-19

R171_187 V171 V187 366.06784177411356
L171_187 V171 V187 -1.5539142037289138e-12
C171_187 V171 V187 -2.061610203120416e-19

R171_188 V171 V188 -108.3538013845011
L171_188 V171 V188 -6.824367696386689e-13
C171_188 V171 V188 -3.132523836006424e-19

R171_189 V171 V189 59.53831112133611
L171_189 V171 V189 -1.2125708182915352e-11
C171_189 V171 V189 -3.968858094793609e-19

R171_190 V171 V190 50.82265931377657
L171_190 V171 V190 1.1991538440022442e-12
C171_190 V171 V190 4.300994005532384e-19

R171_191 V171 V191 67.23208481512613
L171_191 V171 V191 -8.416798509824974e-13
C171_191 V171 V191 -5.381708748758472e-19

R171_192 V171 V192 107.2959980293981
L171_192 V171 V192 6.1258560845813636e-12
C171_192 V171 V192 -2.357348221597832e-19

R171_193 V171 V193 115.9213760200477
L171_193 V171 V193 2.2208502631762265e-12
C171_193 V171 V193 2.5359701567744893e-19

R171_194 V171 V194 -143.3764550211029
L171_194 V171 V194 4.379751506744886e-12
C171_194 V171 V194 -7.236148767142786e-20

R171_195 V171 V195 -35.01895311536795
L171_195 V171 V195 5.395818551496453e-13
C171_195 V171 V195 9.046052618637634e-19

R171_196 V171 V196 130.8459830746044
L171_196 V171 V196 9.281533400513652e-13
C171_196 V171 V196 6.665160317172666e-19

R171_197 V171 V197 -105.63885260641817
L171_197 V171 V197 2.4109003654708987e-12
C171_197 V171 V197 2.6474895240660433e-19

R171_198 V171 V198 -58.70701493192059
L171_198 V171 V198 -1.939377666487599e-12
C171_198 V171 V198 -9.275747206013432e-20

R171_199 V171 V199 727.9226342735157
L171_199 V171 V199 1.7370808761791753e-12
C171_199 V171 V199 2.889000887597231e-19

R171_200 V171 V200 -1975.0008385456722
L171_200 V171 V200 7.99346204070839e-12
C171_200 V171 V200 1.103348129991452e-19

R172_172 V172 0 -2833.0227989450564
L172_172 V172 0 9.260939419420271e-13
C172_172 V172 0 -1.2867448229310502e-18

R172_173 V172 V173 94.23755201327444
L172_173 V172 V173 9.383773030657987e-13
C172_173 V172 V173 3.6233025269565043e-19

R172_174 V172 V174 15.369899159314642
L172_174 V172 V174 3.9327573451786235e-12
C172_174 V172 V174 1.3443373714576074e-19

R172_175 V172 V175 -117.16107903556349
L172_175 V172 V175 -4.088090067300334e-12
C172_175 V172 V175 1.0076361381562765e-22

R172_176 V172 V176 167.56272557165917
L172_176 V172 V176 8.805784842902323e-13
C172_176 V172 V176 9.318917394023587e-20

R172_177 V172 V177 49.61016527662754
L172_177 V172 V177 -6.69071397984541e-12
C172_177 V172 V177 -7.727038290352251e-20

R172_178 V172 V178 -24.230697495522517
L172_178 V172 V178 2.1110454013013786e-11
C172_178 V172 V178 1.6943951075134444e-19

R172_179 V172 V179 162.01996817166338
L172_179 V172 V179 1.885250901241655e-12
C172_179 V172 V179 3.154765338202754e-19

R172_180 V172 V180 14.714625431987864
L172_180 V172 V180 9.225509892171255e-13
C172_180 V172 V180 2.0956561142254138e-19

R172_181 V172 V181 -53.80606099814084
L172_181 V172 V181 -4.485677568764433e-12
C172_181 V172 V181 1.112373272059685e-19

R172_182 V172 V182 -23.754598388534408
L172_182 V172 V182 -9.772932876140655e-13
C172_182 V172 V182 -2.5720569937266495e-19

R172_183 V172 V183 416.1160841419914
L172_183 V172 V183 -1.4392386421894977e-11
C172_183 V172 V183 1.7198910583458046e-20

R172_184 V172 V184 -21.97785229139033
L172_184 V172 V184 -9.441188501116035e-13
C172_184 V172 V184 -5.676441632079083e-20

R172_185 V172 V185 -79.34429137119692
L172_185 V172 V185 7.528241449606902e-12
C172_185 V172 V185 -2.9077445910508687e-20

R172_186 V172 V186 171.33820100137078
L172_186 V172 V186 -2.320628865767252e-12
C172_186 V172 V186 4.277482384047632e-21

R172_187 V172 V187 -296.6362711791843
L172_187 V172 V187 -2.126520444327617e-12
C172_187 V172 V187 -1.7383797834788027e-19

R172_188 V172 V188 87.69203440172193
L172_188 V172 V188 1.0601259432882261e-12
C172_188 V172 V188 -2.7620762356963384e-20

R172_189 V172 V189 69.82145226205672
L172_189 V172 V189 -2.18001047104533e-12
C172_189 V172 V189 -3.142386294240906e-19

R172_190 V172 V190 42.42997995988628
L172_190 V172 V190 1.6845031483558496e-12
C172_190 V172 V190 3.080957923974603e-19

R172_191 V172 V191 129.78340164858972
L172_191 V172 V191 3.6348304505482175e-11
C172_191 V172 V191 -2.433898344830968e-19

R172_192 V172 V192 69.69103418389614
L172_192 V172 V192 -1.0475181160202435e-12
C172_192 V172 V192 -3.79753343327695e-19

R172_193 V172 V193 98.50804602072988
L172_193 V172 V193 4.099484694944698e-12
C172_193 V172 V193 1.0461879831498366e-19

R172_194 V172 V194 -197.89501535119237
L172_194 V172 V194 -1.5923365781876597e-12
C172_194 V172 V194 -2.1925144716684336e-19

R172_195 V172 V195 -187.19807473727354
L172_195 V172 V195 -9.209145552736046e-11
C172_195 V172 V195 4.2955802312343926e-19

R172_196 V172 V196 -43.01349571024478
L172_196 V172 V196 6.169264716822159e-13
C172_196 V172 V196 6.485963097276911e-19

R172_197 V172 V197 -64.07138679486533
L172_197 V172 V197 2.1616516313805836e-12
C172_197 V172 V197 2.9888800653491853e-19

R172_198 V172 V198 -54.71628397939857
L172_198 V172 V198 -4.034056318733326e-12
C172_198 V172 V198 -3.4988319050070516e-20

R172_199 V172 V199 156.39020121108302
L172_199 V172 V199 1.8629411201242836e-12
C172_199 V172 V199 2.8043431186942027e-19

R172_200 V172 V200 -681.2729022974034
L172_200 V172 V200 -1.3920376843229375e-11
C172_200 V172 V200 2.0517453536662746e-20

R173_173 V173 0 -249.47859035876272
L173_173 V173 0 -3.860702314728344e-13
C173_173 V173 0 -4.1905784115857023e-19

R173_174 V173 V174 -30.915843878242786
L173_174 V173 V174 -1.9527943973780595e-12
C173_174 V173 V174 -2.413976292046708e-19

R173_175 V173 V175 68.49593643269718
L173_175 V173 V175 -2.0200095728838407e-12
C173_175 V173 V175 -3.3599972688773413e-19

R173_176 V173 V176 72.86491512447813
L173_176 V173 V176 -1.347623970890772e-12
C173_176 V173 V176 -3.8959178391427953e-19

R173_177 V173 V177 676.3980101877704
L173_177 V173 V177 1.0893518988521884e-12
C173_177 V173 V177 2.4017027768664687e-19

R173_178 V173 V178 42.93577488382122
L173_178 V173 V178 -4.554328326094145e-12
C173_178 V173 V178 -2.0809588174492366e-19

R173_179 V173 V179 -89.93970976265794
L173_179 V173 V179 -1.2337590508568788e-12
C173_179 V173 V179 -1.6916070893723004e-19

R173_180 V173 V180 -138.6419919090316
L173_180 V173 V180 -1.8970510317969625e-12
C173_180 V173 V180 -5.826139210893389e-20

R173_181 V173 V181 54.02140702618344
L173_181 V173 V181 1.3134285158283593e-11
C173_181 V173 V181 3.7828417472757216e-19

R173_182 V173 V182 42.864419314230716
L173_182 V173 V182 9.20689435506385e-13
C173_182 V173 V182 2.496430820758712e-19

R173_183 V173 V183 -193.74048798157267
L173_183 V173 V183 -7.060885712628725e-11
C173_183 V173 V183 7.266474371010139e-20

R173_184 V173 V184 -99.95236986992738
L173_184 V173 V184 2.2090229279679025e-12
C173_184 V173 V184 1.381499964271527e-19

R173_185 V173 V185 -66.72331441076199
L173_185 V173 V185 -7.562446576873618e-12
C173_185 V173 V185 -2.3915987370836766e-19

R173_186 V173 V186 1507.6945168094753
L173_186 V173 V186 8.060569785050361e-13
C173_186 V173 V186 2.3973341779117066e-19

R173_187 V173 V187 178.44013149216372
L173_187 V173 V187 1.277304090305761e-12
C173_187 V173 V187 5.404431442105645e-20

R173_188 V173 V188 622.8112545684004
L173_188 V173 V188 3.1647748030583428e-12
C173_188 V173 V188 7.956132928078236e-20

R173_189 V173 V189 257.62394473699106
L173_189 V173 V189 1.5297245534081813e-12
C173_189 V173 V189 1.1151460687300275e-19

R173_190 V173 V190 -129.7750374398048
L173_190 V173 V190 -1.0806157312776082e-12
C173_190 V173 V190 -3.004725551981427e-19

R173_191 V173 V191 440.1357910519965
L173_191 V173 V191 2.631097212862717e-12
C173_191 V173 V191 1.91429461280066e-19

R173_192 V173 V192 182.7982150146459
L173_192 V173 V192 3.6148107874014428e-12
C173_192 V173 V192 1.0324249033361633e-19

R173_193 V173 V193 145.96571221358576
L173_193 V173 V193 -1.4050019814908139e-12
C173_193 V173 V193 -1.9780998970457103e-19

R173_194 V173 V194 -191.93684305971993
L173_194 V173 V194 -3.1845975867970267e-12
C173_194 V173 V194 1.821080493080643e-19

R173_195 V173 V195 -199.35564213307205
L173_195 V173 V195 -9.482422620628412e-13
C173_195 V173 V195 -3.071845063081397e-19

R173_196 V173 V196 -164.52695774952903
L173_196 V173 V196 -6.255982657828295e-13
C173_196 V173 V196 -4.966676188788554e-19

R173_197 V173 V197 -98.80003732995165
L173_197 V173 V197 -1.7611626106840318e-12
C173_197 V173 V197 -1.5318180084613597e-20

R173_198 V173 V198 49.09496291278436
L173_198 V173 V198 1.4095627868710912e-12
C173_198 V173 V198 7.848671124239635e-20

R173_199 V173 V199 215.52478249694772
L173_199 V173 V199 -2.0157201884955393e-12
C173_199 V173 V199 -2.255597829268167e-19

R173_200 V173 V200 -113.73842458246003
L173_200 V173 V200 2.52808705311632e-11
C173_200 V173 V200 2.7852362970860184e-20

R174_174 V174 0 45.24465020816437
L174_174 V174 0 -2.4495710823705044e-13
C174_174 V174 0 6.048603702847939e-19

R174_175 V174 V175 22.21262898929312
L174_175 V174 V175 -1.6119221656775979e-12
C174_175 V174 V175 -1.9955745297414566e-19

R174_176 V174 V176 15.260805123608087
L174_176 V174 V176 -2.2202457666831173e-12
C174_176 V174 V176 -2.553460828419458e-19

R174_177 V174 V177 -36.30794470814985
L174_177 V174 V177 2.6511771358910073e-12
C174_177 V174 V177 3.319092803712369e-19

R174_178 V174 V178 10.895836133996752
L174_178 V174 V178 9.971841583717376e-13
C174_178 V174 V178 -7.511271270600999e-21

R174_179 V174 V179 -24.76498340213947
L174_179 V174 V179 2.7858432142432525e-11
C174_179 V174 V179 -3.209277890277173e-19

R174_180 V174 V180 -14.8891616136875
L174_180 V174 V180 1.1670875912175861e-11
C174_180 V174 V180 -1.3308646776425797e-19

R174_181 V174 V181 33.88089116110011
L174_181 V174 V181 4.728120613130909e-12
C174_181 V174 V181 2.1156268845668944e-19

R174_182 V174 V182 9.616869803051083
L174_182 V174 V182 6.892217481383086e-13
C174_182 V174 V182 2.7924660893783275e-19

R174_183 V174 V183 -129.46336136665323
L174_183 V174 V183 -1.861580356645417e-11
C174_183 V174 V183 -6.170986788770385e-20

R174_184 V174 V184 -228.71850234223467
L174_184 V174 V184 3.4604144201394568e-12
C174_184 V174 V184 8.346249829785919e-20

R174_185 V174 V185 77.8781073901733
L174_185 V174 V185 1.9333152528990865e-12
C174_185 V174 V185 -3.1309243179282013e-19

R174_186 V174 V186 -25.140117651358562
L174_186 V174 V186 -4.353143718096961e-12
C174_186 V174 V186 1.2915285914870316e-19

R174_187 V174 V187 509.21020846070184
L174_187 V174 V187 8.757141369761773e-12
C174_187 V174 V187 3.6317591636742907e-19

R174_188 V174 V188 68.6422826124845
L174_188 V174 V188 2.5523743434658698e-12
C174_188 V174 V188 3.3416021840259704e-19

R174_189 V174 V189 -66.47378947753481
L174_189 V174 V189 -1.428610830939573e-12
C174_189 V174 V189 1.564606236656178e-19

R174_190 V174 V190 -16.793168781126038
L174_190 V174 V190 -1.8641832290170533e-12
C174_190 V174 V190 -2.3199791769916126e-19

R174_191 V174 V191 215.80796798079083
L174_191 V174 V191 2.7343308230521094e-12
C174_191 V174 V191 2.0609580712370125e-19

R174_192 V174 V192 164.3671314908962
L174_192 V174 V192 -3.320836049135454e-12
C174_192 V174 V192 -4.514415649357959e-20

R174_193 V174 V193 -91.10074353761375
L174_193 V174 V193 -2.642229379321528e-12
C174_193 V174 V193 -2.314940933023291e-19

R174_194 V174 V194 42.79885607799605
L174_194 V174 V194 -1.3577334831533542e-12
C174_194 V174 V194 -3.7698432687649007e-19

R174_195 V174 V195 157.48644628057008
L174_195 V174 V195 -2.469027914816585e-12
C174_195 V174 V195 -4.2288866807070095e-19

R174_196 V174 V196 -318.56026968660495
L174_196 V174 V196 -2.056303649928463e-12
C174_196 V174 V196 -4.673790147570183e-19

R174_197 V174 V197 79.97968804743851
L174_197 V174 V197 1.7090693099076585e-12
C174_197 V174 V197 9.634840736778697e-20

R174_198 V174 V198 15.162001862439912
L174_198 V174 V198 2.2805242869936937e-12
C174_198 V174 V198 1.0593952463515691e-19

R174_199 V174 V199 -356.9572356760484
L174_199 V174 V199 -1.0653155119106322e-11
C174_199 V174 V199 -2.7618237378150106e-19

R174_200 V174 V200 -45.601530198193664
L174_200 V174 V200 3.2380465870915707e-12
C174_200 V174 V200 1.577430927790481e-19

R175_175 V175 0 -247.5815374896194
L175_175 V175 0 -2.36924724604731e-13
C175_175 V175 0 -1.133360111903481e-18

R175_176 V175 V176 471.56696283742076
L175_176 V175 V176 -3.6133396674314366e-12
C175_176 V175 V176 -1.3549393999417162e-19

R175_177 V175 V177 17379.255955363424
L175_177 V175 V177 2.441770541958488e-12
C175_177 V175 V177 2.1428061504111045e-19

R175_178 V175 V178 -54.70821624597912
L175_178 V175 V178 7.632527629351214e-12
C175_178 V175 V178 2.5841558291961435e-20

R175_179 V175 V179 96.8509623961193
L175_179 V175 V179 1.5230071230368687e-12
C175_179 V175 V179 3.472768578435185e-19

R175_180 V175 V180 64.1456103424675
L175_180 V175 V180 3.943769374908574e-12
C175_180 V175 V180 2.4805936057179598e-20

R175_181 V175 V181 -181.68263404778776
L175_181 V175 V181 5.595476281128092e-12
C175_181 V175 V181 3.150002746168865e-19

R175_182 V175 V182 -46.383292373074696
L175_182 V175 V182 -1.942924932432816e-11
C175_182 V175 V182 -4.121921639033437e-20

R175_183 V175 V183 29.982734164406512
L175_183 V175 V183 9.207353550587062e-13
C175_183 V175 V183 -1.8990197905969517e-20

R175_184 V175 V184 -124.60536322239302
L175_184 V175 V184 3.754196126404509e-12
C175_184 V175 V184 1.3937774240952388e-19

R175_185 V175 V185 601.1736974817504
L175_185 V175 V185 5.238166676334907e-12
C175_185 V175 V185 -3.0128323491283294e-19

R175_186 V175 V186 240.6103736278988
L175_186 V175 V186 2.198129106397906e-12
C175_186 V175 V186 2.8571390420891394e-19

R175_187 V175 V187 -55.990505666947044
L175_187 V175 V187 -8.740522639654426e-13
C175_187 V175 V187 -2.8913166825632048e-19

R175_188 V175 V188 538.5551473787431
L175_188 V175 V188 1.8114306060261843e-12
C175_188 V175 V188 5.646662268328545e-20

R175_189 V175 V189 -211.80218677337095
L175_189 V175 V189 -1.6733057999703928e-12
C175_189 V175 V189 -2.362583951407074e-21

R175_190 V175 V190 81.65461846093719
L175_190 V175 V190 1.4782676069344383e-11
C175_190 V175 V190 -2.726004089010727e-20

R175_191 V175 V191 -42.80063909468242
L175_191 V175 V191 7.847536540436566e-11
C175_191 V175 V191 3.6418007339524176e-19

R175_192 V175 V192 -1075.5131466015214
L175_192 V175 V192 -9.493538916454484e-13
C175_192 V175 V192 -2.3031403878914355e-19

R175_193 V175 V193 313.94405136114335
L175_193 V175 V193 -5.20050758551089e-12
C175_193 V175 V193 -1.0856365243602594e-19

R175_194 V175 V194 -784.5610575815858
L175_194 V175 V194 -1.0259453821934882e-12
C175_194 V175 V194 -1.1100320526492948e-19

R175_195 V175 V195 37.55548852504162
L175_195 V175 V195 -4.427833033099635e-12
C175_195 V175 V195 -5.591163016014185e-19

R175_196 V175 V196 -173.2828119267541
L175_196 V175 V196 1.5029358776973123e-12
C175_196 V175 V196 3.051734723135242e-19

R175_197 V175 V197 638.901470868055
L175_197 V175 V197 2.181677712494275e-12
C175_197 V175 V197 2.0040023575888184e-19

R175_198 V175 V198 -62.3700903060984
L175_198 V175 V198 1.1163749881121178e-11
C175_198 V175 V198 4.246646965292617e-21

R175_199 V175 V199 89.86288184469261
L175_199 V175 V199 4.455022367358184e-12
C175_199 V175 V199 -5.3269346956203615e-20

R175_200 V175 V200 210.4254151195894
L175_200 V175 V200 5.854762810377494e-12
C175_200 V175 V200 -6.03913951879878e-20

R176_176 V176 0 -20.138785538946927
L176_176 V176 0 -1.333678242374714e-13
C176_176 V176 0 -2.227009481910998e-18

R176_177 V176 V177 3064.6662936294947
L176_177 V176 V177 1.8493580395920494e-12
C176_177 V176 V177 2.710214991295687e-19

R176_178 V176 V178 -29.280563137926414
L176_178 V176 V178 8.965703721550356e-11
C176_178 V176 V178 4.1686975153209824e-20

R176_179 V176 V179 143.25919112600002
L176_179 V176 V179 3.533842843244212e-11
C176_179 V176 V179 1.5716864597160658e-20

R176_180 V176 V180 92.76107764388864
L176_180 V176 V180 9.252244635762409e-13
C176_180 V176 V180 5.623082198166428e-19

R176_181 V176 V181 -273.79453843171734
L176_181 V176 V181 3.1078371749930556e-12
C176_181 V176 V181 3.9107491239244797e-19

R176_182 V176 V182 -46.25524124381753
L176_182 V176 V182 2.732350253148507e-12
C176_182 V176 V182 6.97051704242093e-20

R176_183 V176 V183 -203.1960973696428
L176_183 V176 V183 6.504233037905627e-12
C176_183 V176 V183 1.3394521049770286e-19

R176_184 V176 V184 25.742222570853514
L176_184 V176 V184 7.232900947018647e-13
C176_184 V176 V184 -3.1398472289540697e-21

R176_185 V176 V185 362.1105954322567
L176_185 V176 V185 3.908966606123317e-12
C176_185 V176 V185 -3.796070312035364e-19

R176_186 V176 V186 53.27690469964822
L176_186 V176 V186 1.0948115363361665e-12
C176_186 V176 V186 1.7578394060436038e-19

R176_187 V176 V187 194.92348243780987
L176_187 V176 V187 1.806394932383875e-12
C176_187 V176 V187 1.6687569719971874e-20

R176_188 V176 V188 -47.579053655221806
L176_188 V176 V188 -7.876039065741265e-13
C176_188 V176 V188 -1.2185865214920597e-19

R176_189 V176 V189 -373.96471964091927
L176_189 V176 V189 -1.6129756252373035e-12
C176_189 V176 V189 -3.080307459971131e-20

R176_190 V176 V190 76.3245482983114
L176_190 V176 V190 -5.544282302923531e-12
C176_190 V176 V190 -2.5771103499916554e-20

R176_191 V176 V191 789.2590096880905
L176_191 V176 V191 -1.9922054690979515e-12
C176_191 V176 V191 -1.9239261786112617e-19

R176_192 V176 V192 -49.02372955953998
L176_192 V176 V192 -5.952229086247622e-11
C176_192 V176 V192 1.9909971468818592e-19

R176_193 V176 V193 891.3492476126753
L176_193 V176 V193 -5.0915064340720476e-12
C176_193 V176 V193 -2.948932485261235e-20

R176_194 V176 V194 -172.4491957367755
L176_194 V176 V194 -1.4132540980359624e-12
C176_194 V176 V194 1.7943194708804193e-20

R176_195 V176 V195 -182.55160107928623
L176_195 V176 V195 1.9910478062436615e-12
C176_195 V176 V195 5.069734066222427e-19

R176_196 V176 V196 47.92361066131216
L176_196 V176 V196 -8.418190936032861e-13
C176_196 V176 V196 -8.54481391186589e-19

R176_197 V176 V197 574.2729703889612
L176_197 V176 V197 2.909349140647086e-12
C176_197 V176 V197 1.884420619372893e-19

R176_198 V176 V198 -49.01062133194857
L176_198 V176 V198 5.184146661745439e-12
C176_198 V176 V198 1.1397965255578075e-19

R176_199 V176 V199 -158.71094497647942
L176_199 V176 V199 -4.3782419759494814e-12
C176_199 V176 V199 -1.994515951453862e-19

R176_200 V176 V200 50.29197587893856
L176_200 V176 V200 9.675306788841128e-13
C176_200 V176 V200 3.623768937957594e-19

R177_177 V177 0 65.53635841185108
L177_177 V177 0 2.411473798568656e-13
C177_177 V177 0 3.5525040377678094e-19

R177_178 V177 V178 98.33449893818403
L177_178 V177 V178 -3.966904713675644e-12
C177_178 V177 V178 -2.370415279064255e-21

R177_179 V177 V179 -123.4006468633263
L177_179 V177 V179 -1.1383651439849793e-11
C177_179 V177 V179 1.2733234736822662e-19

R177_180 V177 V180 -79.40045544211524
L177_180 V177 V180 -4.606742290614382e-12
C177_180 V177 V180 -2.0913805435344095e-20

R177_181 V177 V181 98.33961546336838
L177_181 V177 V181 1.0187216493664684e-12
C177_181 V177 V181 -7.557518535263516e-20

R177_182 V177 V182 49.72409595060636
L177_182 V177 V182 -1.2699688609144648e-11
C177_182 V177 V182 -1.4100253353478643e-19

R177_183 V177 V183 -754.6924368377623
L177_183 V177 V183 -5.747835732369739e-12
C177_183 V177 V183 2.977708030807596e-20

R177_184 V177 V184 417.94888834852185
L177_184 V177 V184 -2.9014135338266576e-12
C177_184 V177 V184 -3.232204108073036e-20

R177_185 V177 V185 39.77952257723669
L177_185 V177 V185 1.1316370781414112e-12
C177_185 V177 V185 2.5264174416744143e-19

R177_186 V177 V186 -133.77083667012963
L177_186 V177 V186 -1.9830064025291124e-12
C177_186 V177 V186 -1.424965485971372e-19

R177_187 V177 V187 2180.9624846856987
L177_187 V177 V187 -6.887766149267228e-12
C177_187 V177 V187 -1.5065776706897995e-19

R177_188 V177 V188 387.6017589500871
L177_188 V177 V188 8.272220830633222e-12
C177_188 V177 V188 -1.7429191056651091e-19

R177_189 V177 V189 -60.58483661845656
L177_189 V177 V189 -1.309523076235416e-12
C177_189 V177 V189 -1.2302637974502894e-19

R177_190 V177 V190 -98.80042778728513
L177_190 V177 V190 1.877836667081902e-11
C177_190 V177 V190 1.1673370434043372e-19

R177_191 V177 V191 159.79752705740233
L177_191 V177 V191 1.738590964376939e-11
C177_191 V177 V191 -1.9363772260928673e-19

R177_192 V177 V192 262.8611174366764
L177_192 V177 V192 -2.15622885901558e-11
C177_192 V177 V192 -3.4259580709033297e-20

R177_193 V177 V193 -54.57503475989963
L177_193 V177 V193 5.5959169376447074e-12
C177_193 V177 V193 1.7856621253256288e-19

R177_194 V177 V194 80.33553924691937
L177_194 V177 V194 1.4993171348221495e-12
C177_194 V177 V194 1.696100269666417e-19

R177_195 V177 V195 1224.1326653719482
L177_195 V177 V195 7.755509355240646e-12
C177_195 V177 V195 2.541458767300923e-19

R177_196 V177 V196 -1101.9543163399987
L177_196 V177 V196 2.244172598063439e-12
C177_196 V177 V196 3.3389891405392e-19

R177_197 V177 V197 58.453082407368065
L177_197 V177 V197 -5.927763486713918e-12
C177_197 V177 V197 -1.594117923719425e-19

R177_198 V177 V198 253.91077394515526
L177_198 V177 V198 -3.0005725984768126e-12
C177_198 V177 V198 -1.0374376224078775e-19

R177_199 V177 V199 -82.66243160965924
L177_199 V177 V199 -4.766232590990589e-12
C177_199 V177 V199 1.731511694214165e-19

R177_200 V177 V200 -97.22929327095457
L177_200 V177 V200 -2.1555981481167565e-12
C177_200 V177 V200 -8.11970948649097e-20

R178_178 V178 0 -28.291779895296727
L178_178 V178 0 7.218355791082021e-13
C178_178 V178 0 8.393723399023726e-19

R178_179 V178 V179 41.191931662383645
L178_179 V178 V179 -2.1307140792488967e-12
C178_179 V178 V179 -2.3372897303955734e-19

R178_180 V178 V180 21.27115188477531
L178_180 V178 V180 -3.2980090580680033e-12
C178_180 V178 V180 -2.0168047584486977e-19

R178_181 V178 V181 -66.96561135426619
L178_181 V178 V181 3.0011382543222732e-12
C178_181 V178 V181 -8.096403462462006e-22

R178_182 V178 V182 -52.467794025477495
L178_182 V178 V182 1.320851354468233e-12
C178_182 V178 V182 1.7586259984888102e-19

R178_183 V178 V183 -329.33561975199717
L178_183 V178 V183 -3.912270458428217e-12
C178_183 V178 V183 -2.768146001977455e-21

R178_184 V178 V184 -126.74164487917558
L178_184 V178 V184 -4.216023828147406e-12
C178_184 V178 V184 8.518437339593588e-21

R178_185 V178 V185 -299.23695447098555
L178_185 V178 V185 -7.003545862303221e-12
C178_185 V178 V185 1.8377232657173206e-20

R178_186 V178 V186 24.959355829541874
L178_186 V178 V186 1.6429990177625118e-12
C178_186 V178 V186 8.329447568151828e-21

R178_187 V178 V187 -230.13242536780092
L178_187 V178 V187 2.2641798706723587e-12
C178_187 V178 V187 9.724373701565561e-20

R178_188 V178 V188 -127.65507963443977
L178_188 V178 V188 1.4287629374571053e-12
C178_188 V178 V188 1.0689130384847564e-19

R178_189 V178 V189 -1093.260319996717
L178_189 V178 V189 -5.705809451509449e-12
C178_189 V178 V189 1.0095786979706429e-19

R178_190 V178 V190 -112.07138012827087
L178_190 V178 V190 -1.5550990297539822e-12
C178_190 V178 V190 -1.7420532720262083e-19

R178_191 V178 V191 -1073.0503310384504
L178_191 V178 V191 3.5118768911319792e-12
C178_191 V178 V191 1.2315783791190568e-19

R178_192 V178 V192 -774.2935059964123
L178_192 V178 V192 -6.4491464923170465e-12
C178_192 V178 V192 9.446124887446124e-20

R178_193 V178 V193 132.2173198597878
L178_193 V178 V193 5.114184482870322e-12
C178_193 V178 V193 -5.666405202701335e-20

R178_194 V178 V194 128.51696397934919
L178_194 V178 V194 3.764566297394871e-12
C178_194 V178 V194 1.1528733259568431e-19

R178_195 V178 V195 -141.25608895423463
L178_195 V178 V195 -1.6621797395549892e-12
C178_195 V178 V195 -2.1169271311822877e-19

R178_196 V178 V196 -209.04043079081947
L178_196 V178 V196 -3.214182293632367e-12
C178_196 V178 V196 -1.9033135713887738e-19

R178_197 V178 V197 146.81851538232962
L178_197 V178 V197 -6.735368519119394e-12
C178_197 V178 V197 -1.503867946797572e-19

R178_198 V178 V198 -82.78242618983124
L178_198 V178 V198 3.2819730156043023e-12
C178_198 V178 V198 4.180754136466777e-20

R178_199 V178 V199 147.4252830572422
L178_199 V178 V199 1.3085662009754756e-10
C178_199 V178 V199 -7.969139443059893e-20

R178_200 V178 V200 58.579922530939925
L178_200 V178 V200 8.112462565091396e-12
C178_200 V178 V200 -9.988969224450276e-20

R179_179 V179 0 -453.47564950060627
L179_179 V179 0 2.740559989968286e-13
C179_179 V179 0 2.4001462881840292e-18

R179_180 V179 V180 -245.63037035516192
L179_180 V179 V180 -9.262953019089763e-13
C179_180 V179 V180 -4.120177689381324e-19

R179_181 V179 V181 119.32490473041736
L179_181 V179 V181 8.381644283604014e-12
C179_181 V179 V181 -1.3074413322967965e-19

R179_182 V179 V182 51.68879229855436
L179_182 V179 V182 7.408367484959332e-13
C179_182 V179 V182 4.557130890309962e-19

R179_183 V179 V183 57.1584085916584
L179_183 V179 V183 -3.165895917352309e-12
C179_183 V179 V183 -5.0289000095313693e-20

R179_184 V179 V184 -169.3696201804659
L179_184 V179 V184 -2.6433888001772996e-12
C179_184 V179 V184 -3.344858691011477e-20

R179_185 V179 V185 366.3647612821085
L179_185 V179 V185 -2.140212265820378e-11
C179_185 V179 V185 1.0191117323655337e-20

R179_186 V179 V186 -118.29135200149517
L179_186 V179 V186 5.325040564164861e-12
C179_186 V179 V186 -9.759285860753378e-20

R179_187 V179 V187 218.67265588602496
L179_187 V179 V187 7.329088527920318e-13
C179_187 V179 V187 6.271918814067581e-19

R179_188 V179 V188 362.659309883679
L179_188 V179 V188 7.511761051592838e-13
C179_188 V179 V188 3.4497203848901563e-19

R179_189 V179 V189 -218.75478499584116
L179_189 V179 V189 3.2004861919124464e-12
C179_189 V179 V189 2.8987866423331065e-19

R179_190 V179 V190 -108.81624642547165
L179_190 V179 V190 -1.4376241378010496e-12
C179_190 V179 V190 -3.7551150205074076e-19

R179_191 V179 V191 -80.83688616866463
L179_191 V179 V191 1.4201413954383817e-12
C179_191 V179 V191 1.3574848149713471e-19

R179_192 V179 V192 4537.186725322441
L179_192 V179 V192 5.1228032468144e-12
C179_192 V179 V192 2.7875500507138596e-19

R179_193 V179 V193 -259.79603838582796
L179_193 V179 V193 -2.8203097172433618e-12
C179_193 V179 V193 -1.9407892101016492e-19

R179_194 V179 V194 1422.2166150243813
L179_194 V179 V194 6.618262300278663e-12
C179_194 V179 V194 -4.988717056583023e-20

R179_195 V179 V195 64.12204094471466
L179_195 V179 V195 -7.089286932909191e-13
C179_195 V179 V195 -3.319602800728886e-19

R179_196 V179 V196 -338.87135894824536
L179_196 V179 V196 -6.580138032375984e-13
C179_196 V179 V196 -7.4882751279308525e-19

R179_197 V179 V197 249.72943563122553
L179_197 V179 V197 -1.6871263010058082e-12
C179_197 V179 V197 -2.3322498020078123e-19

R179_198 V179 V198 68.63723953457166
L179_198 V179 V198 2.0191500385254886e-12
C179_198 V179 V198 9.965398236653841e-20

R179_199 V179 V199 1139.649408286747
L179_199 V179 V199 -1.7764937426471265e-12
C179_199 V179 V199 -2.6703416372052446e-19

R179_200 V179 V200 -404.0709974645997
L179_200 V179 V200 -1.2010324041648244e-11
C179_200 V179 V200 -1.3231776399387984e-21

R180_180 V180 0 651.0058236889641
L180_180 V180 0 2.1104867167959194e-13
C180_180 V180 0 2.876891370415238e-18

R180_181 V180 V181 78.69167018038185
L180_181 V180 V181 7.351207944219473e-12
C180_181 V180 V181 -1.7498499356950742e-19

R180_182 V180 V182 28.92998741393789
L180_182 V180 V182 8.599114637849189e-13
C180_182 V180 V182 2.6819774062430474e-19

R180_183 V180 V183 -89.46052597789283
L180_183 V180 V183 -1.5274946632741918e-12
C180_183 V180 V183 -1.3960237420091834e-19

R180_184 V180 V184 25.19105616942124
L180_184 V180 V184 5.435974438521068e-12
C180_184 V180 V184 9.285268204370487e-20

R180_185 V180 V185 146.58006449651722
L180_185 V180 V185 -5.777541436188739e-12
C180_185 V180 V185 1.0996977885011758e-19

R180_186 V180 V186 -96.03211933916748
L180_186 V180 V186 8.274412149879201e-11
C180_186 V180 V186 -4.548875663744154e-20

R180_187 V180 V187 380.1315872403202
L180_187 V180 V187 1.5492210734363986e-12
C180_187 V180 V187 2.8580564035027487e-19

R180_188 V180 V188 222.61414000342666
L180_188 V180 V188 6.820259540863499e-13
C180_188 V180 V188 3.445966375023566e-19

R180_189 V180 V189 -126.30304635075117
L180_189 V180 V189 2.639341700356872e-12
C180_189 V180 V189 2.0213230113739725e-19

R180_190 V180 V190 -59.159694131489516
L180_190 V180 V190 -1.7844501947178272e-12
C180_190 V180 V190 -2.8642574507989795e-19

R180_191 V180 V191 636.072232331944
L180_191 V180 V191 1.0480261493539242e-12
C180_191 V180 V191 3.588341639683702e-19

R180_192 V180 V192 -47.022770250197915
L180_192 V180 V192 -4.528900621719728e-12
C180_192 V180 V192 -6.360322816246194e-20

R180_193 V180 V193 -124.03155384894137
L180_193 V180 V193 -4.168404258875648e-12
C180_193 V180 V193 -1.4505171446816362e-19

R180_194 V180 V194 2311.1474998986655
L180_194 V180 V194 2.5774925592470024e-12
C180_194 V180 V194 -6.955359593692935e-20

R180_195 V180 V195 -1100.9001982425211
L180_195 V180 V195 -6.548452623405142e-13
C180_195 V180 V195 -8.083576170005708e-19

R180_196 V180 V196 48.933433602437226
L180_196 V180 V196 -1.612563947890846e-12
C180_196 V180 V196 1.965749401420655e-19

R180_197 V180 V197 103.62420938587077
L180_197 V180 V197 -1.6915436912180349e-12
C180_197 V180 V197 -2.0255966673559882e-19

R180_198 V180 V198 47.567931389363416
L180_198 V180 V198 2.1395337146380983e-12
C180_198 V180 V198 -2.461850012724869e-20

R180_199 V180 V199 2521.483078042208
L180_199 V180 V199 -3.020525178406891e-12
C180_199 V180 V199 -1.0029867137178797e-19

R180_200 V180 V200 278.909176860945
L180_200 V180 V200 -2.12309028113486e-12
C180_200 V180 V200 -2.543509726741542e-19

R181_181 V181 0 364.187702622977
L181_181 V181 0 2.447026906940803e-12
C181_181 V181 0 1.3191899004823215e-18

R181_182 V181 V182 -42.115943633556874
L181_182 V181 V182 -2.6965962197671123e-12
C181_182 V181 V182 -1.422095340298216e-20

R181_183 V181 V183 535.3250016995762
L181_183 V181 V183 1.31032929490414e-11
C181_183 V181 V183 -8.956963681982178e-20

R181_184 V181 V184 -9530.241636473362
L181_184 V181 V184 -2.4212749852164844e-11
C181_184 V181 V184 -1.2297582074342544e-19

R181_185 V181 V185 188.0399098112601
L181_185 V181 V185 -4.76386404123137e-11
C181_185 V181 V185 3.9320985681310597e-19

R181_186 V181 V186 1848.3080704288548
L181_186 V181 V186 -3.411088098993749e-12
C181_186 V181 V186 -2.698780458638473e-19

R181_187 V181 V187 -562.5202252776828
L181_187 V181 V187 -4.158799558575583e-12
C181_187 V181 V187 4.012086164822264e-20

R181_188 V181 V188 -1017.7814690865292
L181_188 V181 V188 -3.1002529782477356e-12
C181_188 V181 V188 -4.405916821416375e-20

R181_189 V181 V189 117.01902308997835
L181_189 V181 V189 7.412496176447324e-13
C181_189 V181 V189 3.7633816670783944e-19

R181_190 V181 V190 95.14530171037148
L181_190 V181 V190 2.2385597315623267e-12
C181_190 V181 V190 3.2045308965189375e-21

R181_191 V181 V191 7136.326768547993
L181_191 V181 V191 -8.790787683732493e-10
C181_191 V181 V191 1.7662981467032713e-19

R181_192 V181 V192 1327.4673301490902
L181_192 V181 V192 4.776418915155954e-12
C181_192 V181 V192 3.8973181420834426e-19

R181_193 V181 V193 -154.80188933104094
L181_193 V181 V193 -1.4600061699466718e-12
C181_193 V181 V193 2.163309954830957e-20

R181_194 V181 V194 6194.460943670464
L181_194 V181 V194 5.9487262634638065e-12
C181_194 V181 V194 2.184701515149876e-19

R181_195 V181 V195 861.6250542691641
L181_195 V181 V195 1.5311696530759694e-11
C181_195 V181 V195 -2.356268070560215e-19

R181_196 V181 V196 537.56129382812
L181_196 V181 V196 4.28561777952737e-12
C181_196 V181 V196 -1.762062238982588e-19

R181_197 V181 V197 -1689.8242995974388
L181_197 V181 V197 -4.2527710704300405e-12
C181_197 V181 V197 -3.343085327673317e-19

R181_198 V181 V198 -62.4723047060862
L181_198 V181 V198 -3.224007650734228e-12
C181_198 V181 V198 3.3592291958240352e-21

R181_199 V181 V199 -398.0689125170911
L181_199 V181 V199 -1.5359169249237433e-11
C181_199 V181 V199 4.786822792479592e-20

R181_200 V181 V200 452.699096161054
L181_200 V181 V200 -3.4080269583965515e-12
C181_200 V181 V200 -2.0509081827228688e-19

R182_182 V182 0 370.86828371402504
L182_182 V182 0 -8.746644779501813e-13
C182_182 V182 0 -1.3969149888677589e-18

R182_183 V182 V183 113.21650261495375
L182_183 V182 V183 1.5397742759351576e-12
C182_183 V182 V183 5.43770017150902e-20

R182_184 V182 V184 1910.914179391647
L182_184 V182 V184 1.3523088158296763e-11
C182_184 V182 V184 1.0127706174881761e-21

R182_185 V182 V185 -170.66747938948262
L182_185 V182 V185 -4.3543965098632836e-12
C182_185 V182 V185 6.969236432529735e-20

R182_186 V182 V186 122.49304178515271
L182_186 V182 V186 -2.4300825195799823e-11
C182_186 V182 V186 -2.875530174270544e-20

R182_187 V182 V187 -953.2178342163753
L182_187 V182 V187 -7.684828745735327e-13
C182_187 V182 V187 -3.230801447425624e-19

R182_188 V182 V188 -151.9994008608113
L182_188 V182 V188 -6.919594845920629e-13
C182_188 V182 V188 -2.589497590556222e-19

R182_189 V182 V189 70.82361742734619
L182_189 V182 V189 1.0572500898808664e-11
C182_189 V182 V189 -2.2310299720236664e-19

R182_190 V182 V190 20.058045221632682
L182_190 V182 V190 8.331200506761287e-13
C182_190 V182 V190 3.1996788516181086e-19

R182_191 V182 V191 -305.5799747991368
L182_191 V182 V191 -9.560323536993719e-13
C182_191 V182 V191 -2.0887278910906495e-19

R182_192 V182 V192 -8577.006390665201
L182_192 V182 V192 -4.291863385111471e-12
C182_192 V182 V192 -1.7671904075354608e-19

R182_193 V182 V193 503.6296031434732
L182_193 V182 V193 2.668261940018145e-12
C182_193 V182 V193 1.7916444267920956e-19

R182_194 V182 V194 -45.06233867632417
L182_194 V182 V194 2.0988087184881727e-11
C182_194 V182 V194 1.9494852054072735e-20

R182_195 V182 V195 2067693.283080643
L182_195 V182 V195 5.721725494699588e-13
C182_195 V182 V195 3.662447207577992e-19

R182_196 V182 V196 241.98205512352843
L182_196 V182 V196 4.816221096201346e-13
C182_196 V182 V196 5.497397170696195e-19

R182_197 V182 V197 -114.73857405629782
L182_197 V182 V197 2.3342129592065114e-12
C182_197 V182 V197 1.7492678919178465e-19

R182_198 V182 V198 -22.05581563748955
L182_198 V182 V198 -1.2211408536298592e-12
C182_198 V182 V198 -5.3977199124853376e-20

R182_199 V182 V199 2745.592489427875
L182_199 V182 V199 1.591495509549471e-12
C182_199 V182 V199 2.5231923815970745e-19

R182_200 V182 V200 140.30504171711019
L182_200 V182 V200 -1.6319187902139504e-11
C182_200 V182 V200 2.6785041245365943e-20

R183_183 V183 0 109.62078689267581
L183_183 V183 0 3.8732139253318925e-13
C183_183 V183 0 6.499714353059472e-19

R183_184 V183 V184 129.87273270922088
L183_184 V183 V184 -3.929025513033314e-12
C183_184 V183 V184 2.9530108996221847e-21

R183_185 V183 V185 325.4354451110127
L183_185 V183 V185 1.2865518623882655e-11
C183_185 V183 V185 2.6823765204483877e-20

R183_186 V183 V186 817.1424639423778
L183_186 V183 V186 -5.769590431008071e-12
C183_186 V183 V186 -1.2607290808618902e-20

R183_187 V183 V187 97.24761916156876
L183_187 V183 V187 8.056800397166958e-13
C183_187 V183 V187 6.209955866934886e-20

R183_188 V183 V188 307.04238995240206
L183_188 V183 V188 1.3388315005199221e-12
C183_188 V183 V188 9.463950312060697e-20

R183_189 V183 V189 725.7584841205511
L183_189 V183 V189 1.561121687117049e-11
C183_189 V183 V189 6.596149193173689e-20

R183_190 V183 V190 -198.5027059062477
L183_190 V183 V190 -5.88957507203828e-12
C183_190 V183 V190 -4.605222005439338e-20

R183_191 V183 V191 31.398265745876998
L183_191 V183 V191 1.1471799058260583e-12
C183_191 V183 V191 1.457362139065763e-19

R183_192 V183 V192 3798.2956775417333
L183_192 V183 V192 1.0435311692852594e-11
C183_192 V183 V192 -8.936036909335515e-21

R183_193 V183 V193 -241.91999265198226
L183_193 V183 V193 -4.4532750637152735e-12
C183_193 V183 V193 -4.17654573028713e-20

R183_194 V183 V194 229.95129469972147
L183_194 V183 V194 1.4743828437767308e-11
C183_194 V183 V194 -6.914136248920941e-20

R183_195 V183 V195 -30.155084213911703
L183_195 V183 V195 -8.542292660990724e-13
C183_195 V183 V195 -2.4574745100402746e-19

R183_196 V183 V196 953.1717674576882
L183_196 V183 V196 -1.5969682608928957e-12
C183_196 V183 V196 4.068052711586797e-20

R183_197 V183 V197 -781.6320428867458
L183_197 V183 V197 -4.5378039120241e-12
C183_197 V183 V197 -4.457457266314601e-20

R183_198 V183 V198 422.322607290467
L183_198 V183 V198 7.638239424855035e-12
C183_198 V183 V198 -7.363349034595026e-21

R183_199 V183 V199 -86.46624800606997
L183_199 V183 V199 -2.86856188212868e-12
C183_199 V183 V199 -3.5502950371078144e-20

R183_200 V183 V200 -203.81156776375005
L183_200 V183 V200 -4.530137956398395e-12
C183_200 V183 V200 -5.799091693523372e-20

R184_184 V184 0 26.8231606903837
L184_184 V184 0 2.0557806045048947e-13
C184_184 V184 0 -1.60085979799988e-19

R184_185 V184 V185 -257.96326032136375
L184_185 V184 V185 -9.723208241083733e-12
C184_185 V184 V185 8.537880537230329e-20

R184_186 V184 V186 -160.57165073356552
L184_186 V184 V186 -1.7174589116913415e-12
C184_186 V184 V186 -8.960264933535515e-20

R184_187 V184 V187 -297.42667914588804
L184_187 V184 V187 2.4828778924361205e-11
C184_187 V184 V187 -2.0497899112519803e-20

R184_188 V184 V188 63.111727961515655
L184_188 V184 V188 8.26583956360373e-13
C184_188 V184 V188 2.6342920555680556e-20

R184_189 V184 V189 327.2207646186053
L184_189 V184 V189 8.647628447099617e-12
C184_189 V184 V189 7.912559132205875e-21

R184_190 V184 V190 -598.2991304600426
L184_190 V184 V190 1.575090975444933e-11
C184_190 V184 V190 5.777478605579305e-20

R184_191 V184 V191 440.00554062998197
L184_191 V184 V191 3.045530580046613e-12
C184_191 V184 V191 -2.7714061860718623e-20

R184_192 V184 V192 33.906168191435356
L184_192 V184 V192 6.2266729852838594e-12
C184_192 V184 V192 8.838890516240451e-20

R184_193 V184 V193 295.6741970436475
L184_193 V184 V193 3.083510184158469e-11
C184_193 V184 V193 2.748429391656657e-20

R184_194 V184 V194 155.33152621003177
L184_194 V184 V194 3.798122246422839e-12
C184_194 V184 V194 6.405094718989797e-20

R184_195 V184 V195 1189.1658162837116
L184_195 V184 V195 -2.244329673789768e-12
C184_195 V184 V195 1.4805999663428617e-19

R184_196 V184 V196 -29.96437547975879
L184_196 V184 V196 -4.686976932936924e-12
C184_196 V184 V196 -9.850589468071563e-20

R184_197 V184 V197 -198.1260115892841
L184_197 V184 V197 -8.747758814126853e-12
C184_197 V184 V197 -7.155770677692589e-20

R184_198 V184 V198 336.6913003857473
L184_198 V184 V198 -5.840284532731027e-12
C184_198 V184 V198 1.1494135353145296e-20

R184_199 V184 V199 -1903.2099687378918
L184_199 V184 V199 -5.856604751807077e-12
C184_199 V184 V199 6.4111274206242e-20

R184_200 V184 V200 -62.857075946154026
L184_200 V184 V200 -3.006113236547001e-12
C184_200 V184 V200 -2.9314764830260795e-20

R185_185 V185 0 -77.71271541489344
L185_185 V185 0 -1.482509004221198e-12
C185_185 V185 0 -1.0345198786134139e-18

R185_186 V185 V186 96.81370335447406
L185_186 V185 V186 4.599604151613108e-12
C185_186 V185 V186 2.35706890563554e-19

R185_187 V185 V187 -3423.60242619615
L185_187 V185 V187 -5.2872240237648655e-12
C185_187 V185 V187 3.587425185917528e-20

R185_188 V185 V188 -687.3056694770526
L185_188 V185 V188 -3.065093445048904e-12
C185_188 V185 V188 9.112135777884621e-20

R185_189 V185 V189 59.11146144916768
L185_189 V185 V189 1.4756135293554695e-12
C185_189 V185 V189 -7.414057098387186e-20

R185_190 V185 V190 369.92500450111646
L185_190 V185 V190 1.7040996941211092e-11
C185_190 V185 V190 -5.928249545481034e-20

R185_191 V185 V191 -80.21935568285912
L185_191 V185 V191 -3.2970156554049903e-12
C185_191 V185 V191 3.535013954676138e-20

R185_192 V185 V192 -132.89964688827027
L185_192 V185 V192 5.899335846829236e-12
C185_192 V185 V192 -1.4922896756550957e-19

R185_193 V185 V193 29.055252305743423
L185_193 V185 V193 1.157263174640103e-12
C185_193 V185 V193 -4.999386545849846e-20

R185_194 V185 V194 -59.99933751201708
L185_194 V185 V194 4.3169981492105004e-11
C185_194 V185 V194 -2.1151036119704015e-19

R185_195 V185 V195 930.6124804893439
L185_195 V185 V195 1.0576678066614254e-11
C185_195 V185 V195 -3.081617537852604e-20

R185_196 V185 V196 -654.1743571782779
L185_196 V185 V196 -1.0820294027686795e-11
C185_196 V185 V196 -1.1421845430914754e-19

R185_197 V185 V197 -37.825847232546984
L185_197 V185 V197 -3.362192543764193e-11
C185_197 V185 V197 3.298702185409318e-19

R185_198 V185 V198 107.68261969796616
L185_198 V185 V198 4.32819419367217e-12
C185_198 V185 V198 6.264580151769155e-20

R185_199 V185 V199 49.77505324055291
L185_199 V185 V199 2.3851167301533283e-12
C185_199 V185 V199 -1.3517805631310686e-19

R185_200 V185 V200 63.980222410149175
L185_200 V185 V200 3.661692255320063e-12
C185_200 V185 V200 1.6130789564297644e-19

R186_186 V186 0 33.80489021132693
L186_186 V186 0 2.4765823698851003e-13
C186_186 V186 0 6.331893959335058e-19

R186_187 V186 V187 -429.27387709066795
L186_187 V186 V187 -2.211947289961755e-12
C186_187 V186 V187 5.862876145852969e-20

R186_188 V186 V188 129.51537413293502
L186_188 V186 V188 7.169942502659907e-12
C186_188 V186 V188 5.106725233123344e-22

R186_189 V186 V189 -1247.6712786228147
L186_189 V186 V189 3.5335290918327644e-12
C186_189 V186 V189 5.673439621973896e-20

R186_190 V186 V190 203.87048424966468
L186_190 V186 V190 1.0870971639942675e-12
C186_190 V186 V190 8.742219886962452e-20

R186_191 V186 V191 145.02985093363645
L186_191 V186 V191 2.075262354999241e-12
C186_191 V186 V191 -5.99334461378302e-20

R186_192 V186 V192 135.5242645828233
L186_192 V186 V192 2.4635210822896364e-12
C186_192 V186 V192 1.405079098477807e-19

R186_193 V186 V193 -113.68858222552646
L186_193 V186 V193 7.901468132415677e-12
C186_193 V186 V193 7.342819238022634e-20

R186_194 V186 V194 117.81253844989537
L186_194 V186 V194 2.7649195169389808e-12
C186_194 V186 V194 8.438439800254152e-20

R186_195 V186 V195 346.1003574980374
L186_195 V186 V195 -2.6335022025931536e-11
C186_195 V186 V195 1.1208756734794255e-19

R186_196 V186 V196 -315.6897224085349
L186_196 V186 V196 2.2773974742860544e-12
C186_196 V186 V196 -9.412080839793797e-20

R186_197 V186 V197 -653.4217338104805
L186_197 V186 V197 -1.5483646686168225e-11
C186_197 V186 V197 -2.0194276995548122e-19

R186_198 V186 V198 -298.44122558863694
L186_198 V186 V198 -1.7681247049800744e-12
C186_198 V186 V198 3.1214494916255037e-20

R186_199 V186 V199 -83.86350061471117
L186_199 V186 V199 -7.262187197290926e-12
C186_199 V186 V199 7.48931939766897e-20

R186_200 V186 V200 -73.4548576013108
L186_200 V186 V200 -1.946220802029013e-12
C186_200 V186 V200 -4.867362142730983e-20

R187_187 V187 0 3356.6811375946854
L187_187 V187 0 -1.6268106102265924e-12
C187_187 V187 0 -1.942172799096129e-18

R187_188 V187 V188 477.9971965175492
L187_188 V187 V188 -8.855202735640891e-13
C187_188 V187 V188 -2.8718665355952947e-19

R187_189 V187 V189 -1943.6863623838044
L187_189 V187 V189 -1.2441021051432031e-11
C187_189 V187 V189 -1.7483032267567128e-19

R187_190 V187 V190 1972.7562501203993
L187_190 V187 V190 1.3006312762082867e-12
C187_190 V187 V190 2.6105934850664436e-19

R187_191 V187 V191 -180.48559169586844
L187_191 V187 V191 -2.4135350858370162e-12
C187_191 V187 V191 5.122663283732247e-20

R187_192 V187 V192 -833.6737022526341
L187_192 V187 V192 -2.523675379142644e-12
C187_192 V187 V192 -9.614261199809379e-20

R187_193 V187 V193 619.4762131926306
L187_193 V187 V193 2.143462742515397e-12
C187_193 V187 V193 2.0444903271514426e-19

R187_194 V187 V194 311.76678508740827
L187_194 V187 V194 2.625966728890093e-12
C187_194 V187 V194 2.562457349197364e-19

R187_195 V187 V195 85.54744944799417
L187_195 V187 V195 8.453477032480207e-13
C187_195 V187 V195 1.236056116733227e-19

R187_196 V187 V196 -1925.4011917985902
L187_196 V187 V196 4.777950264509865e-13
C187_196 V187 V196 5.35818709013457e-19

R187_197 V187 V197 -797.8293063856498
L187_197 V187 V197 2.5160919250971646e-12
C187_197 V187 V197 4.708780320685259e-20

R187_198 V187 V198 -532.2654120872907
L187_198 V187 V198 -1.7064302488469793e-12
C187_198 V187 V198 -7.339535335969789e-20

R187_199 V187 V199 684.3278801780282
L187_199 V187 V199 2.9662495217724115e-12
C187_199 V187 V199 2.5175883108631906e-19

R187_200 V187 V200 5404.4556221530365
L187_200 V187 V200 -2.668380343848049e-12
C187_200 V187 V200 -1.3989239693464608e-19

R188_188 V188 0 -46.73604445908895
L188_188 V188 0 -1.5810750300365322e-13
C188_188 V188 0 -1.5996231269479096e-18

R188_189 V188 V189 414.46365419105723
L188_189 V188 V189 2.6517499511866692e-12
C188_189 V188 V189 -9.446750468697804e-20

R188_190 V188 V190 339.4112989688296
L188_190 V188 V190 1.3322510072665572e-12
C188_190 V188 V190 1.7400596705823793e-19

R188_191 V188 V191 -136.59452537992462
L188_191 V188 V191 -5.440693802043326e-13
C188_191 V188 V191 -2.457021345450436e-19

R188_192 V188 V192 -8591.687436301692
L188_192 V188 V192 6.705228014825962e-13
C188_192 V188 V192 2.255362166268882e-19

R188_193 V188 V193 3012.820813270877
L188_193 V188 V193 2.4711279357593408e-12
C188_193 V188 V193 2.152464133962136e-19

R188_194 V188 V194 11077.693132975035
L188_194 V188 V194 1.1280757298934647e-12
C188_194 V188 V194 2.8741588518802675e-19

R188_195 V188 V195 283.01008239986055
L188_195 V188 V195 3.6972034046921823e-13
C188_195 V188 V195 4.937300665416366e-19

R188_196 V188 V196 57.814593503172354
L188_196 V188 V196 2.2187944200459566e-12
C188_196 V188 V196 1.841623122808298e-20

R188_197 V188 V197 -376.1070327437943
L188_197 V188 V197 5.41957568014655e-12
C188_197 V188 V197 -7.667973343128987e-21

R188_198 V188 V198 -159.45918723502663
L188_198 V188 V198 -1.8872302037786494e-12
C188_198 V188 V198 -4.9438952006609056e-20

R188_199 V188 V199 4388.54502386757
L188_199 V188 V199 4.176459658662561e-12
C188_199 V188 V199 8.677513503061557e-20

R188_200 V188 V200 -269.67450151419393
L188_200 V188 V200 -3.914032231008186e-12
C188_200 V188 V200 1.6614616712846728e-20

R189_189 V189 0 -60.87246094461516
L189_189 V189 0 -4.4513721136746334e-13
C189_189 V189 0 -1.1206531574082989e-18

R189_190 V189 V190 -117.3051245693192
L189_190 V189 V190 -3.114150039006492e-12
C189_190 V189 V190 2.5756811633980172e-19

R189_191 V189 V191 525.2865330179982
L189_191 V189 V191 -3.8123478399436914e-12
C189_191 V189 V191 -3.527353151619038e-19

R189_192 V189 V192 -6790.331716829637
L189_192 V189 V192 -1.046380806999927e-12
C189_192 V189 V192 -4.1346368885184067e-19

R189_193 V189 V193 -161.32184302864545
L189_193 V189 V193 9.695762859959597e-13
C189_193 V189 V193 2.1172378887765647e-19

R189_194 V189 V194 194.12947921065327
L189_194 V189 V194 -1.3786958697975847e-12
C189_194 V189 V194 -1.3933105240388023e-19

R189_195 V189 V195 1847.4781005723994
L189_195 V189 V195 3.444301889756241e-12
C189_195 V189 V195 5.639904500268801e-19

R189_196 V189 V196 -515.1422474311438
L189_196 V189 V196 2.731894144677014e-12
C189_196 V189 V196 6.082045577972906e-19

R189_197 V189 V197 48.11325846317951
L189_197 V189 V197 1.0094393853331568e-12
C189_197 V189 V197 3.0466407597987577e-19

R189_198 V189 V198 193.66917168734514
L189_198 V189 V198 2.698390816255673e-12
C189_198 V189 V198 -6.463205466505214e-20

R189_199 V189 V199 -345.5219246562612
L189_199 V189 V199 3.2066985898126533e-12
C189_199 V189 V199 2.1362873824110014e-19

R189_200 V189 V200 -683.3342863332603
L189_200 V189 V200 1.5772436848115917e-12
C189_200 V189 V200 1.2184277735900173e-19

R190_190 V190 0 -490.30853129464765
L190_190 V190 0 -8.307579607779667e-13
C190_190 V190 0 1.6342773753087999e-18

R190_191 V190 V191 -331.3625532959854
L190_191 V190 V191 6.052116088241112e-12
C190_191 V190 V191 2.226904015895547e-19

R190_192 V190 V192 -2055.8780638662006
L190_192 V190 V192 -1.1367615011661364e-11
C190_192 V190 V192 1.672707753788265e-19

R190_193 V190 V193 3431.635238449962
L190_193 V190 V193 -5.119526491733877e-12
C190_193 V190 V193 -1.8432818116507892e-19

R190_194 V190 V194 58.11135093450283
L190_194 V190 V194 6.72024687146934e-12
C190_194 V190 V194 2.948725469757778e-20

R190_195 V190 V195 729.1024772832473
L190_195 V190 V195 -1.723161272701973e-12
C190_195 V190 V195 -4.537818230986902e-19

R190_196 V190 V196 -256.04050118123786
L190_196 V190 V196 -1.0440720908764772e-12
C190_196 V190 V196 -4.3251356118975965e-19

R190_197 V190 V197 115.66377854797025
L190_197 V190 V197 2.335887517204647e-11
C190_197 V190 V197 -1.7208542226177173e-19

R190_198 V190 V198 29.82991515902927
L190_198 V190 V198 1.1546368827425941e-12
C190_198 V190 V198 6.096250232422009e-21

R190_199 V190 V199 283.96298129139365
L190_199 V190 V199 -1.768905346220259e-11
C190_199 V190 V199 -2.7944425118027973e-19

R190_200 V190 V200 509.51235942696684
L190_200 V190 V200 2.940145283668064e-12
C190_200 V190 V200 -2.7088816371365523e-20

R191_191 V191 0 -69.50404952561544
L191_191 V191 0 -2.389235750961092e-13
C191_191 V191 0 -1.0774681631467367e-18

R191_192 V191 V192 -154.93948950577501
L191_192 V191 V192 4.846981737652738e-12
C191_192 V191 V192 -1.5281058589781396e-19

R191_193 V191 V193 88.4892241991763
L191_193 V191 V193 1.8876420277306256e-12
C191_193 V191 V193 1.701865389813719e-19

R191_194 V191 V194 -120.77898603659258
L191_194 V191 V194 9.081599808468583e-12
C191_194 V191 V194 -3.0231874652091553e-20

R191_195 V191 V195 35.12222125165226
L191_195 V191 V195 4.019763645692875e-13
C191_195 V191 V195 1.1115827148688683e-18

R191_196 V191 V196 328.09139847713556
L191_196 V191 V196 3.860685755713312e-12
C191_196 V191 V196 8.274326041125962e-20

R191_197 V191 V197 -586.1109580297862
L191_197 V191 V197 2.581572186238722e-12
C191_197 V191 V197 2.17806283240094e-19

R191_198 V191 V198 196.47069611353848
L191_198 V191 V198 2.5832803696004672e-11
C191_198 V191 V198 -5.312963054146607e-20

R191_199 V191 V199 53.84493242405963
L191_199 V191 V199 1.3791292667936655e-12
C191_199 V191 V199 1.769693659016107e-19

R191_200 V191 V200 75.84044592184406
L191_200 V191 V200 1.935043957832504e-12
C191_200 V191 V200 2.975532275924296e-19

R192_192 V192 0 -28.355144941192716
L192_192 V192 0 -8.419806472336578e-13
C192_192 V192 0 -7.171874839439214e-20

R192_193 V192 V193 146.53063393169222
L192_193 V192 V193 6.4984291863745054e-12
C192_193 V192 V193 -7.131347881426277e-21

R192_194 V192 V194 -112.60996673762273
L192_194 V192 V194 -8.967231175552888e-13
C192_194 V192 V194 -4.3265395090789067e-19

R192_195 V192 V195 245.88849920605776
L192_195 V192 V195 -1.4825583088555072e-12
C192_195 V192 V195 4.5459059915295243e-20

R192_196 V192 V196 58.065279382299764
L192_196 V192 V196 5.314888449847992e-13
C192_196 V192 V196 1.0576041899044336e-18

R192_197 V192 V197 -1038.4022434918468
L192_197 V192 V197 1.9057120992446427e-12
C192_197 V192 V197 4.282335778380299e-19

R192_198 V192 V198 219.81058160033263
L192_198 V192 V198 3.0500725339094796e-12
C192_198 V192 V198 -8.771491931658263e-20

R192_199 V192 V199 93.30015944891736
L192_199 V192 V199 1.7202552730764728e-12
C192_199 V192 V199 2.0091881705732147e-19

R192_200 V192 V200 48.34644354416273
L192_200 V192 V200 1.5026758686585443e-12
C192_200 V192 V200 9.682160344035263e-20

R193_193 V193 0 54.743844654543174
L193_193 V193 0 -1.4344570146248764e-12
C193_193 V193 0 6.1586028449606105e-19

R193_194 V193 V194 72.99993582159982
L193_194 V193 V194 5.9809422040846245e-12
C193_194 V193 V194 -1.1739801182841553e-19

R193_195 V193 V195 -2321.4807121378713
L193_195 V193 V195 -2.153178270354196e-12
C193_195 V193 V195 -3.4534295498162127e-19

R193_196 V193 V196 241.79799579916315
L193_196 V193 V196 -3.0237507910720966e-12
C193_196 V193 V196 -1.868620290182669e-19

R193_197 V193 V197 46.56922457305068
L193_197 V193 V197 4.940050638553876e-12
C193_197 V193 V197 -1.9283442207710634e-20

R193_198 V193 V198 -117.62687628964838
L193_198 V193 V198 -2.8077916147031587e-11
C193_198 V193 V198 3.4404378954734315e-20

R193_199 V193 V199 -58.31645286012606
L193_199 V193 V199 -1.7570658737155775e-12
C193_199 V193 V199 -1.3676812877698313e-19

R193_200 V193 V200 -59.00986578630204
L193_200 V193 V200 -2.346332217862965e-12
C193_200 V193 V200 -1.192408438316485e-20

R194_194 V194 0 -65.25416480434228
L194_194 V194 0 -3.226943537776482e-13
C194_194 V194 0 5.442845331903584e-19

R194_195 V194 V195 -3545.185280129953
L194_195 V194 V195 -2.923146898160784e-12
C194_195 V194 V195 -1.3144180640136585e-19

R194_196 V194 V196 705.3961636874504
L194_196 V194 V196 3.6086191202896102e-12
C194_196 V194 V196 3.401247064548208e-19

R194_197 V194 V197 -265.79443212247946
L194_197 V194 V197 3.861477028256788e-12
C194_197 V194 V197 3.212669629154241e-19

R194_198 V194 V198 -400.0330387664443
L194_198 V194 V198 1.9373004289963237e-12
C194_198 V194 V198 3.4177574327504235e-20

R194_199 V194 V199 72.00231407713756
L194_199 V194 V199 3.4822643097370154e-12
C194_199 V194 V199 -6.689797286930486e-20

R194_200 V194 V200 65.67514342638636
L194_200 V194 V200 1.3789078574347054e-12
C194_200 V194 V200 1.8052054441124404e-19

R195_195 V195 0 370.58891206318134
L195_195 V195 0 2.002662348618664e-13
C195_195 V195 0 3.2046540710320547e-18

R195_196 V195 V196 -421.60772770071117
L195_196 V195 V196 -1.2028553499491023e-12
C195_196 V195 V196 1.1470628417721834e-19

R195_197 V195 V197 1490.505281656796
L195_197 V195 V197 -1.2460529512256529e-12
C195_197 V195 V197 -3.148283759717909e-19

R195_198 V195 V198 -902.057984380959
L195_198 V195 V198 3.0000327794122534e-12
C195_198 V195 V198 1.238832592593469e-20

R195_199 V195 V199 -143.04351621992606
L195_199 V195 V199 -1.767226200829372e-12
C195_199 V195 V199 -3.2490481487811943e-19

R195_200 V195 V200 -316.180470874877
L195_200 V195 V200 -2.173859790229374e-12
C195_200 V195 V200 -4.2110691824022683e-19

R196_196 V196 0 36.15050010214348
L196_196 V196 0 -2.1655683630778223e-12
C196_196 V196 0 1.276914628418997e-19

R196_197 V196 V197 1338.4007764697362
L196_197 V196 V197 -1.1262939031965004e-12
C196_197 V196 V197 -5.072081260068081e-19

R196_198 V196 V198 287.55459793779147
L196_198 V196 V198 1.721378906366985e-12
C196_198 V196 V198 2.446559050260708e-19

R196_199 V196 V199 -1953.3912969374696
L196_199 V196 V199 -9.495452284971155e-13
C196_199 V196 V199 -5.213261126697608e-19

R196_200 V196 V200 -527.7147883143963
L196_200 V196 V200 1.9200076721098264e-12
C196_200 V196 V200 2.3471083037412596e-19

R197_197 V197 0 63.46007724741369
L197_197 V197 0 2.1447024512244507e-13
C197_197 V197 0 1.5426565404035257e-18

R197_198 V197 V198 -333.1007349853041
L197_198 V197 V198 -3.857223141007912e-12
C197_198 V197 V198 1.3751784170093913e-20

R197_199 V197 V199 541.1826122211806
L197_199 V197 V199 -1.738960143680197e-12
C197_199 V197 V199 -1.0362614628578958e-19

R197_200 V197 V200 -1015.3856335863234
L197_200 V197 V200 -1.867478575290406e-12
C197_200 V197 V200 -2.167829448253643e-19

R198_198 V198 0 44.91497735552347
L198_198 V198 0 4.4394872630477206e-13
C198_198 V198 0 4.0857579388022885e-19

R198_199 V198 V199 -65.61836720929374
L198_199 V198 V199 -4.394192117597473e-12
C198_199 V198 V199 2.6418188877297945e-20

R198_200 V198 V200 -302.8875078858766
L198_200 V198 V200 -2.3822581213478022e-12
C198_200 V198 V200 2.5361185540226937e-21

R199_199 V199 0 21.227757455934732
L199_199 V199 0 3.532887238935711e-13
C199_199 V199 0 1.2206939055385753e-18

R199_200 V199 V200 -63.36704148577402
L199_200 V199 V200 -1.9385849649454347e-12
C199_200 V199 V200 9.077069276174104e-20

R200_200 V200 0 36.841390535026065
L200_200 V200 0 2.1862098091294462e-13
C200_200 V200 0 3.9075676392312116e-19

ISRC1_p1 0 V1  ac 1.064553385934121e-01*Ip1
ISRC1_p2 0 V1  ac 9.885765551539263e-03*Ip2
ISRC1_p3 0 V1  ac 1.407097011782252e-02*Ip3
ISRC1_p4 0 V1  ac 1.246401772639715e-02*Ip4

ISRC2_p1 0 V2  ac -3.289874922314183e-02*Ip1
ISRC2_p2 0 V2  ac 1.151348703301520e-01*Ip2
ISRC2_p3 0 V2  ac 1.208308238763943e-02*Ip3
ISRC2_p4 0 V2  ac 1.404957179831909e-02*Ip4

ISRC3_p1 0 V3  ac -2.509892529706435e-02*Ip1
ISRC3_p2 0 V3  ac -3.174423885616620e-02*Ip2
ISRC3_p3 0 V3  ac 1.294002244417553e-01*Ip3
ISRC3_p4 0 V3  ac 3.112103832951167e-03*Ip4

ISRC4_p1 0 V4  ac -1.954126116031075e-02*Ip1
ISRC4_p2 0 V4  ac -2.754089886761033e-02*Ip2
ISRC4_p3 0 V4  ac -2.433399909658278e-02*Ip3
ISRC4_p4 0 V4  ac 1.418953874747593e-01*Ip4

ISRC5_p1 0 V5  ac 3.977279028018596e-02*Ip1
ISRC5_p2 0 V5  ac 8.998875849843853e-03*Ip2
ISRC5_p3 0 V5  ac 1.012527959263409e-02*Ip3
ISRC5_p4 0 V5  ac 1.268646725409618e-02*Ip4

ISRC6_p1 0 V6  ac -7.637529762056741e-03*Ip1
ISRC6_p2 0 V6  ac 1.782299303554434e-02*Ip2
ISRC6_p3 0 V6  ac 1.903545198954385e-02*Ip3
ISRC6_p4 0 V6  ac 2.186315488804201e-02*Ip4

ISRC7_p1 0 V7  ac -6.034088753907411e-03*Ip1
ISRC7_p2 0 V7  ac -6.605244120468883e-03*Ip2
ISRC7_p3 0 V7  ac -1.220788946719124e-02*Ip3
ISRC7_p4 0 V7  ac 3.761607789154967e-02*Ip4

ISRC8_p1 0 V8  ac 9.677876337867933e-04*Ip1
ISRC8_p2 0 V8  ac -1.947809160723713e-04*Ip2
ISRC8_p3 0 V8  ac -1.748820315209653e-03*Ip3
ISRC8_p4 0 V8  ac -5.103676500195518e-02*Ip4

ISRC9_p1 0 V9  ac -8.469330962994324e-02*Ip1
ISRC9_p2 0 V9  ac 4.188545909805909e-03*Ip2
ISRC9_p3 0 V9  ac 2.124005020098187e-03*Ip3
ISRC9_p4 0 V9  ac 3.749404573261545e-03*Ip4

ISRC10_p1 0 V10  ac 9.534056792040479e-03*Ip1
ISRC10_p2 0 V10  ac -5.333099815344879e-02*Ip2
ISRC10_p3 0 V10  ac -3.158046509419913e-04*Ip3
ISRC10_p4 0 V10  ac -1.417055112745353e-03*Ip4

ISRC11_p1 0 V11  ac 1.156198658093865e-02*Ip1
ISRC11_p2 0 V11  ac 1.219653006860806e-02*Ip2
ISRC11_p3 0 V11  ac -3.959434098941371e-02*Ip3
ISRC11_p4 0 V11  ac -6.853675605346481e-03*Ip4

ISRC12_p1 0 V12  ac 7.861785738433491e-03*Ip1
ISRC12_p2 0 V12  ac 1.186607359060020e-02*Ip2
ISRC12_p3 0 V12  ac 1.037637620836932e-02*Ip3
ISRC12_p4 0 V12  ac -2.708870824692164e-02*Ip4

ISRC13_p1 0 V13  ac 3.094509028002145e-02*Ip1
ISRC13_p2 0 V13  ac 3.454371605918731e-03*Ip2
ISRC13_p3 0 V13  ac 4.166447826200361e-03*Ip3
ISRC13_p4 0 V13  ac 6.039882183935082e-03*Ip4

ISRC14_p1 0 V14  ac -1.071170649510741e-02*Ip1
ISRC14_p2 0 V14  ac 1.752779916338945e-02*Ip2
ISRC14_p3 0 V14  ac 8.689764838044787e-03*Ip3
ISRC14_p4 0 V14  ac 1.194936203782196e-02*Ip4

ISRC15_p1 0 V15  ac -9.534946905422947e-03*Ip1
ISRC15_p2 0 V15  ac -5.437714900034983e-03*Ip2
ISRC15_p3 0 V15  ac 1.712003741361888e-03*Ip3
ISRC15_p4 0 V15  ac 1.715937693256592e-02*Ip4

ISRC16_p1 0 V16  ac -6.327890355247883e-03*Ip1
ISRC16_p2 0 V16  ac -3.073074028508607e-03*Ip2
ISRC16_p3 0 V16  ac -3.169228959279274e-03*Ip3
ISRC16_p4 0 V16  ac -1.421349775304866e-02*Ip4

ISRC17_p1 0 V17  ac -5.101879789818612e-03*Ip1
ISRC17_p2 0 V17  ac -3.078579601669633e-03*Ip2
ISRC17_p3 0 V17  ac -4.024171576769096e-03*Ip3
ISRC17_p4 0 V17  ac -6.436577683489982e-03*Ip4

ISRC18_p1 0 V18  ac 3.797747910509557e-04*Ip1
ISRC18_p2 0 V18  ac 6.714406212632103e-04*Ip2
ISRC18_p3 0 V18  ac -9.739888162112763e-03*Ip3
ISRC18_p4 0 V18  ac -1.446927970010249e-02*Ip4

ISRC19_p1 0 V19  ac -1.251044410573520e-03*Ip1
ISRC19_p2 0 V19  ac -7.642152608904459e-04*Ip2
ISRC19_p3 0 V19  ac -3.086164138027966e-03*Ip3
ISRC19_p4 0 V19  ac -9.488481560116495e-03*Ip4

ISRC20_p1 0 V20  ac -2.108799359782761e-03*Ip1
ISRC20_p2 0 V20  ac -1.153852719636614e-03*Ip2
ISRC20_p3 0 V20  ac -4.891932747269603e-03*Ip3
ISRC20_p4 0 V20  ac -1.126664199800508e-02*Ip4

ISRC21_p1 0 V21  ac 6.276094647060905e-02*Ip1
ISRC21_p2 0 V21  ac -3.442237073245447e-03*Ip2
ISRC21_p3 0 V21  ac -2.499409603884970e-03*Ip3
ISRC21_p4 0 V21  ac -4.725819952106287e-03*Ip4

ISRC22_p1 0 V22  ac -7.355013721468268e-03*Ip1
ISRC22_p2 0 V22  ac 3.048918559166735e-02*Ip2
ISRC22_p3 0 V22  ac 3.831684767846498e-03*Ip3
ISRC22_p4 0 V22  ac 3.952797235236571e-03*Ip4

ISRC23_p1 0 V23  ac -7.047139662162913e-03*Ip1
ISRC23_p2 0 V23  ac -6.303118658173635e-03*Ip2
ISRC23_p3 0 V23  ac 2.501044696035065e-02*Ip3
ISRC23_p4 0 V23  ac 1.737379112855615e-03*Ip4

ISRC24_p1 0 V24  ac -5.015532505739845e-03*Ip1
ISRC24_p2 0 V24  ac -6.565142836976160e-03*Ip2
ISRC24_p3 0 V24  ac -3.566842491611761e-03*Ip3
ISRC24_p4 0 V24  ac 1.634603251732231e-02*Ip4

ISRC25_p1 0 V25  ac -6.299452169639454e-02*Ip1
ISRC25_p2 0 V25  ac -4.191224307968065e-03*Ip2
ISRC25_p3 0 V25  ac -3.909031479721647e-03*Ip3
ISRC25_p4 0 V25  ac -6.016313326859806e-03*Ip4

ISRC26_p1 0 V26  ac 7.993155239201497e-03*Ip1
ISRC26_p2 0 V26  ac -2.497564636120427e-02*Ip2
ISRC26_p3 0 V26  ac -1.229186519171024e-02*Ip3
ISRC26_p4 0 V26  ac -1.795361653890191e-02*Ip4

ISRC27_p1 0 V27  ac 8.624353694309113e-03*Ip1
ISRC27_p2 0 V27  ac 5.451316583042930e-03*Ip2
ISRC27_p3 0 V27  ac -1.755023596477593e-02*Ip3
ISRC27_p4 0 V27  ac -1.642426920182681e-02*Ip4

ISRC28_p1 0 V28  ac 5.835139927730089e-03*Ip1
ISRC28_p2 0 V28  ac 4.983160941345400e-03*Ip2
ISRC28_p3 0 V28  ac 2.048161515035386e-03*Ip3
ISRC28_p4 0 V28  ac -1.357512204334800e-02*Ip4

ISRC29_p1 0 V29  ac -4.934243596917237e-02*Ip1
ISRC29_p2 0 V29  ac 3.911679640121136e-03*Ip2
ISRC29_p3 0 V29  ac 3.078602819360878e-03*Ip3
ISRC29_p4 0 V29  ac 3.713740665566660e-03*Ip4

ISRC30_p1 0 V30  ac 6.720116614696111e-03*Ip1
ISRC30_p2 0 V30  ac -2.906308340434324e-02*Ip2
ISRC30_p3 0 V30  ac 2.054760169267779e-03*Ip3
ISRC30_p4 0 V30  ac 3.297032137136703e-03*Ip4

ISRC31_p1 0 V31  ac 7.553407390817403e-03*Ip1
ISRC31_p2 0 V31  ac 3.348565045215622e-03*Ip2
ISRC31_p3 0 V31  ac -6.339784081834158e-03*Ip3
ISRC31_p4 0 V31  ac -4.269130439006110e-03*Ip4

ISRC32_p1 0 V32  ac 3.857358101066122e-03*Ip1
ISRC32_p2 0 V32  ac 1.866499616267574e-03*Ip2
ISRC32_p3 0 V32  ac 5.696979201072420e-03*Ip3
ISRC32_p4 0 V32  ac 1.864196714842760e-02*Ip4

ISRC33_p1 0 V33  ac -4.410104431199773e-02*Ip1
ISRC33_p2 0 V33  ac -7.918700505729201e-03*Ip2
ISRC33_p3 0 V33  ac -8.617302425782675e-03*Ip3
ISRC33_p4 0 V33  ac -1.010767595652246e-02*Ip4

ISRC34_p1 0 V34  ac 8.764988302185524e-03*Ip1
ISRC34_p2 0 V34  ac -1.288071382302024e-02*Ip2
ISRC34_p3 0 V34  ac -1.156362392435279e-02*Ip3
ISRC34_p4 0 V34  ac -1.363441475596117e-02*Ip4

ISRC35_p1 0 V35  ac 8.644795439710883e-03*Ip1
ISRC35_p2 0 V35  ac 4.629609822747795e-03*Ip2
ISRC35_p3 0 V35  ac -4.698205686700862e-04*Ip3
ISRC35_p4 0 V35  ac -1.712431116640557e-02*Ip4

ISRC36_p1 0 V36  ac 4.411167806607764e-03*Ip1
ISRC36_p2 0 V36  ac 2.643570340983159e-03*Ip2
ISRC36_p3 0 V36  ac 2.045267609037755e-03*Ip3
ISRC36_p4 0 V36  ac 2.726178511453871e-02*Ip4

ISRC37_p1 0 V37  ac 2.763030193182794e-02*Ip1
ISRC37_p2 0 V37  ac -5.689804748402769e-03*Ip2
ISRC37_p3 0 V37  ac -3.810418838006437e-03*Ip3
ISRC37_p4 0 V37  ac -3.618520701049493e-03*Ip4

ISRC38_p1 0 V38  ac -4.432488259461918e-04*Ip1
ISRC38_p2 0 V38  ac 1.368188604733325e-02*Ip2
ISRC38_p3 0 V38  ac -4.433735449132514e-03*Ip3
ISRC38_p4 0 V38  ac -2.162522463299118e-03*Ip4

ISRC39_p1 0 V39  ac -3.066799762576146e-03*Ip1
ISRC39_p2 0 V39  ac -2.960093333005583e-03*Ip2
ISRC39_p3 0 V39  ac 1.599366814737212e-02*Ip3
ISRC39_p4 0 V39  ac -6.913012326041273e-03*Ip4

ISRC40_p1 0 V40  ac -4.249149407101513e-03*Ip1
ISRC40_p2 0 V40  ac -4.669118231644642e-03*Ip2
ISRC40_p3 0 V40  ac -3.494684231099457e-03*Ip3
ISRC40_p4 0 V40  ac 2.316110041720301e-02*Ip4

ISRC41_p1 0 V41  ac -2.532952498923222e-02*Ip1
ISRC41_p2 0 V41  ac -2.965087322408071e-03*Ip2
ISRC41_p3 0 V41  ac -2.192274783298315e-03*Ip3
ISRC41_p4 0 V41  ac -3.395848178839711e-03*Ip4

ISRC42_p1 0 V42  ac 3.164874988926015e-03*Ip1
ISRC42_p2 0 V42  ac -1.769864281596540e-04*Ip2
ISRC42_p3 0 V42  ac -7.908004713214923e-03*Ip3
ISRC42_p4 0 V42  ac -1.212091149067668e-02*Ip4

ISRC43_p1 0 V43  ac 3.844432778475996e-03*Ip1
ISRC43_p2 0 V43  ac 3.932030887783973e-03*Ip2
ISRC43_p3 0 V43  ac 2.665916258915953e-03*Ip3
ISRC43_p4 0 V43  ac -1.017995605068883e-02*Ip4

ISRC44_p1 0 V44  ac 2.279457104326765e-03*Ip1
ISRC44_p2 0 V44  ac 3.685737082374333e-03*Ip2
ISRC44_p3 0 V44  ac 3.943672707701714e-03*Ip3
ISRC44_p4 0 V44  ac 8.778674512055509e-03*Ip4

ISRC45_p1 0 V45  ac -2.341612629248979e-02*Ip1
ISRC45_p2 0 V45  ac 1.207137358718455e-03*Ip2
ISRC45_p3 0 V45  ac 1.369904547784649e-03*Ip3
ISRC45_p4 0 V45  ac 6.982087370800037e-04*Ip4

ISRC46_p1 0 V46  ac 1.745634132138401e-03*Ip1
ISRC46_p2 0 V46  ac -3.608130902226872e-03*Ip2
ISRC46_p3 0 V46  ac 2.066957513204919e-03*Ip3
ISRC46_p4 0 V46  ac 4.962106998202304e-04*Ip4

ISRC47_p1 0 V47  ac 4.709696545089532e-03*Ip1
ISRC47_p2 0 V47  ac 3.909060741851198e-03*Ip2
ISRC47_p3 0 V47  ac -5.080183349852568e-03*Ip3
ISRC47_p4 0 V47  ac -2.776750388030336e-04*Ip4

ISRC48_p1 0 V48  ac 3.772187001815300e-03*Ip1
ISRC48_p2 0 V48  ac 4.350499893641255e-03*Ip2
ISRC48_p3 0 V48  ac 4.087425824627722e-03*Ip3
ISRC48_p4 0 V48  ac -8.647719456494282e-03*Ip4

ISRC49_p1 0 V49  ac -5.090487530944270e-02*Ip1
ISRC49_p2 0 V49  ac -3.270407887088175e-03*Ip2
ISRC49_p3 0 V49  ac -6.257032032392691e-03*Ip3
ISRC49_p4 0 V49  ac -9.033939941003585e-03*Ip4

ISRC50_p1 0 V50  ac 8.627511470398072e-03*Ip1
ISRC50_p2 0 V50  ac -1.612587733462518e-02*Ip2
ISRC50_p3 0 V50  ac -9.763761931455292e-03*Ip3
ISRC50_p4 0 V50  ac -1.277903317812252e-02*Ip4

ISRC51_p1 0 V51  ac 9.349647151883201e-03*Ip1
ISRC51_p2 0 V51  ac 4.490765252069876e-03*Ip2
ISRC51_p3 0 V51  ac -4.919317748534397e-03*Ip3
ISRC51_p4 0 V51  ac -1.821800312198825e-02*Ip4

ISRC52_p1 0 V52  ac 7.493704074601864e-03*Ip1
ISRC52_p2 0 V52  ac 3.597163735013071e-03*Ip2
ISRC52_p3 0 V52  ac 1.169660116085664e-03*Ip3
ISRC52_p4 0 V52  ac 1.649956679022428e-02*Ip4

ISRC53_p1 0 V53  ac 1.087702420716670e-03*Ip1
ISRC53_p2 0 V53  ac -4.095994661093978e-03*Ip2
ISRC53_p3 0 V53  ac -5.745609139713166e-03*Ip3
ISRC53_p4 0 V53  ac -5.615030704099642e-03*Ip4

ISRC54_p1 0 V54  ac 2.969940940361963e-03*Ip1
ISRC54_p2 0 V54  ac 7.543388004127026e-03*Ip2
ISRC54_p3 0 V54  ac -7.567761966826809e-03*Ip3
ISRC54_p4 0 V54  ac -4.853639690926584e-03*Ip4

ISRC55_p1 0 V55  ac 7.945660773770325e-04*Ip1
ISRC55_p2 0 V55  ac 2.145836287990734e-03*Ip2
ISRC55_p3 0 V55  ac 4.465499651673252e-03*Ip3
ISRC55_p4 0 V55  ac -8.019814516018174e-03*Ip4

ISRC56_p1 0 V56  ac -1.256834826740014e-03*Ip1
ISRC56_p2 0 V56  ac 1.191711587028407e-03*Ip2
ISRC56_p3 0 V56  ac -3.373783586799434e-03*Ip3
ISRC56_p4 0 V56  ac 2.733016846393329e-02*Ip4

ISRC57_p1 0 V57  ac -2.232602797754398e-02*Ip1
ISRC57_p2 0 V57  ac -4.551574462164671e-03*Ip2
ISRC57_p3 0 V57  ac -6.084014788918131e-03*Ip3
ISRC57_p4 0 V57  ac -8.822816978112016e-03*Ip4

ISRC58_p1 0 V58  ac 1.018722953110818e-02*Ip1
ISRC58_p2 0 V58  ac -1.612426742028542e-02*Ip2
ISRC58_p3 0 V58  ac -3.625469270237909e-03*Ip3
ISRC58_p4 0 V58  ac -7.261709982161198e-03*Ip4

ISRC59_p1 0 V59  ac 7.339729996322285e-03*Ip1
ISRC59_p2 0 V59  ac 2.185078097454532e-03*Ip2
ISRC59_p3 0 V59  ac -7.368489681682210e-03*Ip3
ISRC59_p4 0 V59  ac -9.807266624957929e-03*Ip4

ISRC60_p1 0 V60  ac 7.174496982814181e-03*Ip1
ISRC60_p2 0 V60  ac 1.774953324906171e-03*Ip2
ISRC60_p3 0 V60  ac -2.075582947728587e-04*Ip3
ISRC60_p4 0 V60  ac -2.526978702432712e-04*Ip4

ISRC61_p1 0 V61  ac 4.527382996279265e-03*Ip1
ISRC61_p2 0 V61  ac 2.830217699361713e-03*Ip2
ISRC61_p3 0 V61  ac 3.699623516277351e-03*Ip3
ISRC61_p4 0 V61  ac 5.880181677497633e-03*Ip4

ISRC62_p1 0 V62  ac -2.950552315040490e-03*Ip1
ISRC62_p2 0 V62  ac 6.128203343700713e-03*Ip2
ISRC62_p3 0 V62  ac -6.105861912131524e-04*Ip3
ISRC62_p4 0 V62  ac -8.809327608619626e-04*Ip4

ISRC63_p1 0 V63  ac -9.115321685990989e-04*Ip1
ISRC63_p2 0 V63  ac -4.896094466020496e-04*Ip2
ISRC63_p3 0 V63  ac 6.696011265926864e-03*Ip3
ISRC63_p4 0 V63  ac -1.057510598737472e-03*Ip4

ISRC64_p1 0 V64  ac -2.139917258604182e-03*Ip1
ISRC64_p2 0 V64  ac -1.242332739091441e-03*Ip2
ISRC64_p3 0 V64  ac 2.393143712728887e-03*Ip3
ISRC64_p4 0 V64  ac 1.693594248285024e-02*Ip4

ISRC65_p1 0 V65  ac -4.349005836961142e-02*Ip1
ISRC65_p2 0 V65  ac -3.044158925196999e-03*Ip2
ISRC65_p3 0 V65  ac -4.582039871029183e-03*Ip3
ISRC65_p4 0 V65  ac -7.485707683256867e-03*Ip4

ISRC66_p1 0 V66  ac 5.403565938467778e-03*Ip1
ISRC66_p2 0 V66  ac -1.285607568322445e-02*Ip2
ISRC66_p3 0 V66  ac -9.481278639243291e-03*Ip3
ISRC66_p4 0 V66  ac -1.234212406817545e-02*Ip4

ISRC67_p1 0 V67  ac 3.701893249635747e-03*Ip1
ISRC67_p2 0 V67  ac 2.340491262082087e-03*Ip2
ISRC67_p3 0 V67  ac -6.162577723510735e-03*Ip3
ISRC67_p4 0 V67  ac -7.807788087699882e-03*Ip4

ISRC68_p1 0 V68  ac 2.357991777170757e-03*Ip1
ISRC68_p2 0 V68  ac 2.258228695382048e-03*Ip2
ISRC68_p3 0 V68  ac -1.605513136109961e-03*Ip3
ISRC68_p4 0 V68  ac 1.838259553753410e-03*Ip4

ISRC69_p1 0 V69  ac -6.983974595464238e-03*Ip1
ISRC69_p2 0 V69  ac 6.441898783751959e-04*Ip2
ISRC69_p3 0 V69  ac -3.862235518706718e-03*Ip3
ISRC69_p4 0 V69  ac 1.551376865508921e-03*Ip4

ISRC70_p1 0 V70  ac 4.741984598391168e-03*Ip1
ISRC70_p2 0 V70  ac -7.488137883177536e-03*Ip2
ISRC70_p3 0 V70  ac 4.647965850133573e-03*Ip3
ISRC70_p4 0 V70  ac 9.797084506301037e-03*Ip4

ISRC71_p1 0 V71  ac 6.511751127016892e-03*Ip1
ISRC71_p2 0 V71  ac 1.447640194077371e-03*Ip2
ISRC71_p3 0 V71  ac -1.417592299222011e-02*Ip3
ISRC71_p4 0 V71  ac 1.348212592908153e-02*Ip4

ISRC72_p1 0 V72  ac 1.107634813001143e-02*Ip1
ISRC72_p2 0 V72  ac 2.988637334016987e-03*Ip2
ISRC72_p3 0 V72  ac -2.065689446984980e-04*Ip3
ISRC72_p4 0 V72  ac -1.525650606191884e-02*Ip4

ISRC73_p1 0 V73  ac 4.236996807445851e-03*Ip1
ISRC73_p2 0 V73  ac -1.023722947635832e-02*Ip2
ISRC73_p3 0 V73  ac -8.801811968805725e-03*Ip3
ISRC73_p4 0 V73  ac -1.156799565781176e-02*Ip4

ISRC74_p1 0 V74  ac 1.582925025942338e-03*Ip1
ISRC74_p2 0 V74  ac -2.070634729703284e-03*Ip2
ISRC74_p3 0 V74  ac -2.456618069464487e-03*Ip3
ISRC74_p4 0 V74  ac -3.597653853537358e-03*Ip4

ISRC75_p1 0 V75  ac -1.879063220677189e-03*Ip1
ISRC75_p2 0 V75  ac -4.035913552856572e-03*Ip2
ISRC75_p3 0 V75  ac 1.122928072525312e-02*Ip3
ISRC75_p4 0 V75  ac -1.685112556736483e-02*Ip4

ISRC76_p1 0 V76  ac -3.997288541227213e-03*Ip1
ISRC76_p2 0 V76  ac -5.656459867536486e-03*Ip2
ISRC76_p3 0 V76  ac 7.432246403578978e-04*Ip3
ISRC76_p4 0 V76  ac 1.859863103304499e-02*Ip4

ISRC77_p1 0 V77  ac -9.316616218590109e-03*Ip1
ISRC77_p2 0 V77  ac -1.569016860919551e-03*Ip2
ISRC77_p3 0 V77  ac 4.761199461208163e-03*Ip3
ISRC77_p4 0 V77  ac 5.093403555299010e-04*Ip4

ISRC78_p1 0 V78  ac -4.460196224767124e-03*Ip1
ISRC78_p2 0 V78  ac -3.478450943499225e-03*Ip2
ISRC78_p3 0 V78  ac 8.235212902705576e-03*Ip3
ISRC78_p4 0 V78  ac 4.967656317267365e-03*Ip4

ISRC79_p1 0 V79  ac -2.776365881509120e-03*Ip1
ISRC79_p2 0 V79  ac 1.463187581714342e-03*Ip2
ISRC79_p3 0 V79  ac 1.437636521216112e-02*Ip3
ISRC79_p4 0 V79  ac -3.715456106099636e-04*Ip4

ISRC80_p1 0 V80  ac -3.596268823511706e-03*Ip1
ISRC80_p2 0 V80  ac 1.824859274423669e-03*Ip2
ISRC80_p3 0 V80  ac 1.083341969952222e-02*Ip3
ISRC80_p4 0 V80  ac 1.392832780020418e-02*Ip4

ISRC81_p1 0 V81  ac -7.022847241727172e-02*Ip1
ISRC81_p2 0 V81  ac -6.297291286270419e-03*Ip2
ISRC81_p3 0 V81  ac 4.719198422020762e-05*Ip3
ISRC81_p4 0 V81  ac -9.875603132643098e-03*Ip4

ISRC82_p1 0 V82  ac 1.098447027041419e-02*Ip1
ISRC82_p2 0 V82  ac -6.478680570717284e-03*Ip2
ISRC82_p3 0 V82  ac -3.408974315909798e-03*Ip3
ISRC82_p4 0 V82  ac -7.390580731378229e-03*Ip4

ISRC83_p1 0 V83  ac 2.068452916086180e-02*Ip1
ISRC83_p2 0 V83  ac 5.831370912791993e-03*Ip2
ISRC83_p3 0 V83  ac 4.055208806637234e-03*Ip3
ISRC83_p4 0 V83  ac -1.821917570683409e-02*Ip4

ISRC84_p1 0 V84  ac 1.427210330187201e-02*Ip1
ISRC84_p2 0 V84  ac 4.977124945309690e-03*Ip2
ISRC84_p3 0 V84  ac 4.795109554287330e-03*Ip3
ISRC84_p4 0 V84  ac 1.320181019086249e-02*Ip4

ISRC85_p1 0 V85  ac -8.442092113149604e-03*Ip1
ISRC85_p2 0 V85  ac 8.792116183070775e-03*Ip2
ISRC85_p3 0 V85  ac 4.111416460587654e-03*Ip3
ISRC85_p4 0 V85  ac 6.510384312423102e-03*Ip4

ISRC86_p1 0 V86  ac 2.794675000082851e-02*Ip1
ISRC86_p2 0 V86  ac -8.905437434395569e-03*Ip2
ISRC86_p3 0 V86  ac -4.770473718398365e-03*Ip3
ISRC86_p4 0 V86  ac -6.391538764491039e-03*Ip4

ISRC87_p1 0 V87  ac 5.185778705875230e-03*Ip1
ISRC87_p2 0 V87  ac 3.245476677559363e-03*Ip2
ISRC87_p3 0 V87  ac -1.286848925570786e-02*Ip3
ISRC87_p4 0 V87  ac 5.686932429862197e-03*Ip4

ISRC88_p1 0 V88  ac 8.914219336067590e-03*Ip1
ISRC88_p2 0 V88  ac 4.028686797344659e-03*Ip2
ISRC88_p3 0 V88  ac 1.883376421241431e-03*Ip3
ISRC88_p4 0 V88  ac -2.149874753567729e-02*Ip4

ISRC89_p1 0 V89  ac -3.192662058064219e-03*Ip1
ISRC89_p2 0 V89  ac -3.280181739791781e-03*Ip2
ISRC89_p3 0 V89  ac -7.432375723756647e-03*Ip3
ISRC89_p4 0 V89  ac -9.476358408880472e-03*Ip4

ISRC90_p1 0 V90  ac -1.756005579429375e-02*Ip1
ISRC90_p2 0 V90  ac 1.101657262851554e-02*Ip2
ISRC90_p3 0 V90  ac -8.207373415918429e-03*Ip3
ISRC90_p4 0 V90  ac -1.530986161796139e-02*Ip4

ISRC91_p1 0 V91  ac -4.613197032756059e-03*Ip1
ISRC91_p2 0 V91  ac 5.663191973650803e-03*Ip2
ISRC91_p3 0 V91  ac 4.064797286071130e-03*Ip3
ISRC91_p4 0 V91  ac -1.104299744267396e-02*Ip4

ISRC92_p1 0 V92  ac 1.831807600581663e-03*Ip1
ISRC92_p2 0 V92  ac 4.868058951730602e-03*Ip2
ISRC92_p3 0 V92  ac 2.322968246695981e-03*Ip3
ISRC92_p4 0 V92  ac 3.689614040490742e-02*Ip4

ISRC93_p1 0 V93  ac -2.265962377968248e-02*Ip1
ISRC93_p2 0 V93  ac -8.715313767176682e-03*Ip2
ISRC93_p3 0 V93  ac -4.141801336405042e-03*Ip3
ISRC93_p4 0 V93  ac -1.212551638221688e-02*Ip4

ISRC94_p1 0 V94  ac -1.139471722023971e-02*Ip1
ISRC94_p2 0 V94  ac 1.441837969141160e-02*Ip2
ISRC94_p3 0 V94  ac -1.550808076741854e-03*Ip3
ISRC94_p4 0 V94  ac -7.629957586578746e-03*Ip4

ISRC95_p1 0 V95  ac -4.943656181522936e-03*Ip1
ISRC95_p2 0 V95  ac -4.519609227269510e-03*Ip2
ISRC95_p3 0 V95  ac 8.275129018377304e-03*Ip3
ISRC95_p4 0 V95  ac 2.479422814734026e-04*Ip4

ISRC96_p1 0 V96  ac -1.221898667419119e-02*Ip1
ISRC96_p2 0 V96  ac -5.561638818003388e-03*Ip2
ISRC96_p3 0 V96  ac -1.846275855110432e-03*Ip3
ISRC96_p4 0 V96  ac -6.295618963235728e-03*Ip4

ISRC97_p1 0 V97  ac -3.852719646230263e-02*Ip1
ISRC97_p2 0 V97  ac 2.859112454327756e-03*Ip2
ISRC97_p3 0 V97  ac -2.752116419127173e-03*Ip3
ISRC97_p4 0 V97  ac -7.346953850715947e-03*Ip4

ISRC98_p1 0 V98  ac 4.600000495711222e-02*Ip1
ISRC98_p2 0 V98  ac -3.299259542288193e-02*Ip2
ISRC98_p3 0 V98  ac 6.705881251327870e-04*Ip3
ISRC98_p4 0 V98  ac 2.881508623358328e-03*Ip4

ISRC99_p1 0 V99  ac 3.770513776080353e-02*Ip1
ISRC99_p2 0 V99  ac 1.652265319663298e-02*Ip2
ISRC99_p3 0 V99  ac -1.333504681650178e-02*Ip3
ISRC99_p4 0 V99  ac -1.964851519648511e-02*Ip4

ISRC100_p1 0 V100  ac 3.670005359095647e-02*Ip1
ISRC100_p2 0 V100  ac 1.687783931522490e-02*Ip2
ISRC100_p3 0 V100  ac 1.145039269267273e-02*Ip3
ISRC100_p4 0 V100  ac 4.028320969819161e-03*Ip4

ISRC101_p1 0 V101  ac -2.185513748227067e-04*Ip1
ISRC101_p2 0 V101  ac -4.555741391468536e-03*Ip2
ISRC101_p3 0 V101  ac -5.302194998663588e-03*Ip3
ISRC101_p4 0 V101  ac -1.352061982850475e-02*Ip4

ISRC102_p1 0 V102  ac 1.094316251880759e-03*Ip1
ISRC102_p2 0 V102  ac 5.897876691271365e-03*Ip2
ISRC102_p3 0 V102  ac -3.222088255297933e-04*Ip3
ISRC102_p4 0 V102  ac -1.310169687764743e-03*Ip4

ISRC103_p1 0 V103  ac 3.345390593829145e-03*Ip1
ISRC103_p2 0 V103  ac -3.388663613326631e-03*Ip2
ISRC103_p3 0 V103  ac 8.610083960219743e-03*Ip3
ISRC103_p4 0 V103  ac -9.049043080685220e-03*Ip4

ISRC104_p1 0 V104  ac 4.579089142799786e-03*Ip1
ISRC104_p2 0 V104  ac -4.309155107563545e-03*Ip2
ISRC104_p3 0 V104  ac -2.307124205762066e-03*Ip3
ISRC104_p4 0 V104  ac 1.015900885356369e-02*Ip4

ISRC105_p1 0 V105  ac -6.714045947806549e-02*Ip1
ISRC105_p2 0 V105  ac -5.248416729482176e-03*Ip2
ISRC105_p3 0 V105  ac -7.563743191631118e-03*Ip3
ISRC105_p4 0 V105  ac -8.053516609652027e-03*Ip4

ISRC106_p1 0 V106  ac 5.803492302237197e-03*Ip1
ISRC106_p2 0 V106  ac -1.024808771095798e-02*Ip2
ISRC106_p3 0 V106  ac -2.142613818914409e-03*Ip3
ISRC106_p4 0 V106  ac -1.239275833141363e-03*Ip4

ISRC107_p1 0 V107  ac -8.080147037114857e-03*Ip1
ISRC107_p2 0 V107  ac -3.524533096303123e-03*Ip2
ISRC107_p3 0 V107  ac -6.296397990490722e-03*Ip3
ISRC107_p4 0 V107  ac 1.443669961398773e-03*Ip4

ISRC108_p1 0 V108  ac -8.401322833657946e-03*Ip1
ISRC108_p2 0 V108  ac -3.474044111865911e-03*Ip2
ISRC108_p3 0 V108  ac -7.760423361325197e-03*Ip3
ISRC108_p4 0 V108  ac -2.139263749567766e-02*Ip4

ISRC109_p1 0 V109  ac 1.470597047515707e-02*Ip1
ISRC109_p2 0 V109  ac 3.680075898045226e-03*Ip2
ISRC109_p3 0 V109  ac -6.083924748872178e-03*Ip3
ISRC109_p4 0 V109  ac -5.644657330200380e-03*Ip4

ISRC110_p1 0 V110  ac -6.106375711274602e-03*Ip1
ISRC110_p2 0 V110  ac 1.951896243721862e-03*Ip2
ISRC110_p3 0 V110  ac 4.062247751301749e-03*Ip3
ISRC110_p4 0 V110  ac 1.050901155074040e-02*Ip4

ISRC111_p1 0 V111  ac 1.048998485368235e-02*Ip1
ISRC111_p2 0 V111  ac 7.249631197415612e-03*Ip2
ISRC111_p3 0 V111  ac -2.824838430175881e-02*Ip3
ISRC111_p4 0 V111  ac 1.196955253397806e-02*Ip4

ISRC112_p1 0 V112  ac 1.555387711015356e-02*Ip1
ISRC112_p2 0 V112  ac 8.717600471887908e-03*Ip2
ISRC112_p3 0 V112  ac -6.995061827642067e-05*Ip3
ISRC112_p4 0 V112  ac -1.719959237852735e-02*Ip4

ISRC113_p1 0 V113  ac -1.622541318800517e-02*Ip1
ISRC113_p2 0 V113  ac -8.198592072597159e-03*Ip2
ISRC113_p3 0 V113  ac 2.207846971428019e-03*Ip3
ISRC113_p4 0 V113  ac 5.113648493720657e-03*Ip4

ISRC114_p1 0 V114  ac 4.909802248907243e-03*Ip1
ISRC114_p2 0 V114  ac 2.872182897348084e-03*Ip2
ISRC114_p3 0 V114  ac 3.611809020140942e-03*Ip3
ISRC114_p4 0 V114  ac 9.379230965223508e-03*Ip4

ISRC115_p1 0 V115  ac 8.754918597668002e-03*Ip1
ISRC115_p2 0 V115  ac -4.966965341061574e-03*Ip2
ISRC115_p3 0 V115  ac -3.846986014471723e-03*Ip3
ISRC115_p4 0 V115  ac 1.341168533370973e-02*Ip4

ISRC116_p1 0 V116  ac 5.932674047511899e-03*Ip1
ISRC116_p2 0 V116  ac -4.787917284804065e-03*Ip2
ISRC116_p3 0 V116  ac 3.024425175735793e-03*Ip3
ISRC116_p4 0 V116  ac 1.289703448141753e-03*Ip4

ISRC117_p1 0 V117  ac -3.878998164284536e-02*Ip1
ISRC117_p2 0 V117  ac -1.814052169573436e-03*Ip2
ISRC117_p3 0 V117  ac -4.641111772407185e-03*Ip3
ISRC117_p4 0 V117  ac -1.505256799862051e-03*Ip4

ISRC118_p1 0 V118  ac 9.164705990736032e-03*Ip1
ISRC118_p2 0 V118  ac -1.274711274220891e-02*Ip2
ISRC118_p3 0 V118  ac -3.393060157595444e-03*Ip3
ISRC118_p4 0 V118  ac -1.675215639105227e-03*Ip4

ISRC119_p1 0 V119  ac 2.230601630632587e-03*Ip1
ISRC119_p2 0 V119  ac 1.933052420227220e-04*Ip2
ISRC119_p3 0 V119  ac -1.004150014919197e-02*Ip3
ISRC119_p4 0 V119  ac 5.839363426097100e-03*Ip4

ISRC120_p1 0 V120  ac 8.525816943504495e-03*Ip1
ISRC120_p2 0 V120  ac 2.026456354856588e-03*Ip2
ISRC120_p3 0 V120  ac -3.128680806845299e-03*Ip3
ISRC120_p4 0 V120  ac -1.928805013066257e-03*Ip4

ISRC121_p1 0 V121  ac -1.327719260607884e-02*Ip1
ISRC121_p2 0 V121  ac -5.993487168116922e-03*Ip2
ISRC121_p3 0 V121  ac -1.109993577555694e-02*Ip3
ISRC121_p4 0 V121  ac -1.214448099560918e-02*Ip4

ISRC122_p1 0 V122  ac 5.094912859981850e-03*Ip1
ISRC122_p2 0 V122  ac -8.554035166477091e-03*Ip2
ISRC122_p3 0 V122  ac -1.635787688971508e-03*Ip3
ISRC122_p4 0 V122  ac 5.627924379089261e-03*Ip4

ISRC123_p1 0 V123  ac 2.687223271800871e-03*Ip1
ISRC123_p2 0 V123  ac -8.245727028496800e-04*Ip2
ISRC123_p3 0 V123  ac -9.100231166051862e-04*Ip3
ISRC123_p4 0 V123  ac -4.600047829870858e-03*Ip4

ISRC124_p1 0 V124  ac -6.273939053177414e-03*Ip1
ISRC124_p2 0 V124  ac -3.770668217384737e-03*Ip2
ISRC124_p3 0 V124  ac -3.413960371187892e-03*Ip3
ISRC124_p4 0 V124  ac 7.727428884169710e-03*Ip4

ISRC125_p1 0 V125  ac -2.572235509103546e-02*Ip1
ISRC125_p2 0 V125  ac 1.905641148807220e-03*Ip2
ISRC125_p3 0 V125  ac -2.079579844713993e-03*Ip3
ISRC125_p4 0 V125  ac 1.039234442371656e-03*Ip4

ISRC126_p1 0 V126  ac -5.505557442320114e-03*Ip1
ISRC126_p2 0 V126  ac 1.035689003141785e-02*Ip2
ISRC126_p3 0 V126  ac 1.294480885164417e-02*Ip3
ISRC126_p4 0 V126  ac 2.333218985087444e-02*Ip4

ISRC127_p1 0 V127  ac -6.713064655025361e-03*Ip1
ISRC127_p2 0 V127  ac -3.245007935507910e-03*Ip2
ISRC127_p3 0 V127  ac 6.050303314071669e-03*Ip3
ISRC127_p4 0 V127  ac 1.787732565675711e-02*Ip4

ISRC128_p1 0 V128  ac -7.996003232790417e-03*Ip1
ISRC128_p2 0 V128  ac -2.021139148010768e-03*Ip2
ISRC128_p3 0 V128  ac 1.246492275567762e-03*Ip3
ISRC128_p4 0 V128  ac -1.225534609709604e-02*Ip4

ISRC129_p1 0 V129  ac -4.766392815144431e-03*Ip1
ISRC129_p2 0 V129  ac 5.860137166510808e-04*Ip2
ISRC129_p3 0 V129  ac 6.618924844710068e-03*Ip3
ISRC129_p4 0 V129  ac 4.612618237510146e-03*Ip4

ISRC130_p1 0 V130  ac -6.056524882365515e-04*Ip1
ISRC130_p2 0 V130  ac -7.887843577311898e-03*Ip2
ISRC130_p3 0 V130  ac 6.825801943115826e-03*Ip3
ISRC130_p4 0 V130  ac 4.948571901724662e-03*Ip4

ISRC131_p1 0 V131  ac 1.261406625415807e-02*Ip1
ISRC131_p2 0 V131  ac 3.792224004291014e-03*Ip2
ISRC131_p3 0 V131  ac -6.556717893936332e-04*Ip3
ISRC131_p4 0 V131  ac -1.428376836981988e-02*Ip4

ISRC132_p1 0 V132  ac 2.764520085054679e-02*Ip1
ISRC132_p2 0 V132  ac 4.187390399527384e-03*Ip2
ISRC132_p3 0 V132  ac 4.693476383943962e-03*Ip3
ISRC132_p4 0 V132  ac -1.562294170076672e-03*Ip4

ISRC133_p1 0 V133  ac 2.480156460481891e-02*Ip1
ISRC133_p2 0 V133  ac -6.177835531011336e-03*Ip2
ISRC133_p3 0 V133  ac 3.882174059461310e-03*Ip3
ISRC133_p4 0 V133  ac 9.497913913734337e-03*Ip4

ISRC134_p1 0 V134  ac 1.144794077648058e-02*Ip1
ISRC134_p2 0 V134  ac -1.940487035420162e-02*Ip2
ISRC134_p3 0 V134  ac 3.734803763693945e-03*Ip3
ISRC134_p4 0 V134  ac 1.274902709353365e-02*Ip4

ISRC135_p1 0 V135  ac -7.915591217097884e-03*Ip1
ISRC135_p2 0 V135  ac -1.045033501616771e-02*Ip2
ISRC135_p3 0 V135  ac -1.346634052265049e-02*Ip3
ISRC135_p4 0 V135  ac 1.544020000103929e-02*Ip4

ISRC136_p1 0 V136  ac -1.148693946544295e-02*Ip1
ISRC136_p2 0 V136  ac -1.260126670736977e-02*Ip2
ISRC136_p3 0 V136  ac -7.502502615857376e-03*Ip3
ISRC136_p4 0 V136  ac -7.309603295467193e-03*Ip4

ISRC137_p1 0 V137  ac -4.427486835070243e-02*Ip1
ISRC137_p2 0 V137  ac -1.261024529014118e-02*Ip2
ISRC137_p3 0 V137  ac -1.105568619255578e-02*Ip3
ISRC137_p4 0 V137  ac -2.068166422768994e-03*Ip4

ISRC138_p1 0 V138  ac -2.448010248026448e-02*Ip1
ISRC138_p2 0 V138  ac 1.262305162351754e-02*Ip2
ISRC138_p3 0 V138  ac 8.708606574147638e-03*Ip3
ISRC138_p4 0 V138  ac 1.279277418294510e-02*Ip4

ISRC139_p1 0 V139  ac 5.212478990784465e-03*Ip1
ISRC139_p2 0 V139  ac 3.194856281248549e-03*Ip2
ISRC139_p3 0 V139  ac 1.099572104511356e-03*Ip3
ISRC139_p4 0 V139  ac 1.947867811800501e-02*Ip4

ISRC140_p1 0 V140  ac 7.055065919251113e-03*Ip1
ISRC140_p2 0 V140  ac 3.418137041952891e-03*Ip2
ISRC140_p3 0 V140  ac 1.307111000418973e-02*Ip3
ISRC140_p4 0 V140  ac 6.589412666971300e-03*Ip4

ISRC141_p1 0 V141  ac 2.362196010933740e-02*Ip1
ISRC141_p2 0 V141  ac 1.164407094131003e-03*Ip2
ISRC141_p3 0 V141  ac -7.881875559396619e-03*Ip3
ISRC141_p4 0 V141  ac -1.044912389919838e-03*Ip4

ISRC142_p1 0 V142  ac 2.372623821345798e-02*Ip1
ISRC142_p2 0 V142  ac -1.741431350883275e-02*Ip2
ISRC142_p3 0 V142  ac -1.299373804111490e-02*Ip3
ISRC142_p4 0 V142  ac -6.493289871902621e-03*Ip4

ISRC143_p1 0 V143  ac 1.387163273253914e-02*Ip1
ISRC143_p2 0 V143  ac 1.644476355537701e-04*Ip2
ISRC143_p3 0 V143  ac -2.746411852639585e-02*Ip3
ISRC143_p4 0 V143  ac -4.264974932036757e-03*Ip4

ISRC144_p1 0 V144  ac 1.060076840625014e-02*Ip1
ISRC144_p2 0 V144  ac 2.043514071926547e-03*Ip2
ISRC144_p3 0 V144  ac -1.307578729835372e-02*Ip3
ISRC144_p4 0 V144  ac 3.892086589426044e-02*Ip4

ISRC145_p1 0 V145  ac -4.787821429284701e-02*Ip1
ISRC145_p2 0 V145  ac 3.350333520627571e-03*Ip2
ISRC145_p3 0 V145  ac 1.200174989441409e-02*Ip3
ISRC145_p4 0 V145  ac 5.697427221591206e-03*Ip4

ISRC146_p1 0 V146  ac 2.064301657773689e-02*Ip1
ISRC146_p2 0 V146  ac 2.250760136584003e-02*Ip2
ISRC146_p3 0 V146  ac 9.862468350515796e-03*Ip3
ISRC146_p4 0 V146  ac 1.313338153197388e-03*Ip4

ISRC147_p1 0 V147  ac -1.443291473427060e-02*Ip1
ISRC147_p2 0 V147  ac 5.894269894845359e-03*Ip2
ISRC147_p3 0 V147  ac 8.330551785054904e-02*Ip3
ISRC147_p4 0 V147  ac 1.005503052923308e-02*Ip4

ISRC148_p1 0 V148  ac -1.457162173496649e-02*Ip1
ISRC148_p2 0 V148  ac -7.812179107000578e-03*Ip2
ISRC148_p3 0 V148  ac 1.872718918512845e-02*Ip3
ISRC148_p4 0 V148  ac -4.505821382284891e-02*Ip4

ISRC149_p1 0 V149  ac 7.803965338572787e-02*Ip1
ISRC149_p2 0 V149  ac -1.128895202231376e-02*Ip2
ISRC149_p3 0 V149  ac -1.520916154967457e-02*Ip3
ISRC149_p4 0 V149  ac -2.595827502037034e-02*Ip4

ISRC150_p1 0 V150  ac -1.838145257209180e-02*Ip1
ISRC150_p2 0 V150  ac -6.456058233474332e-02*Ip2
ISRC150_p3 0 V150  ac -2.628387307415905e-02*Ip3
ISRC150_p4 0 V150  ac -3.280759713796646e-02*Ip4

ISRC151_p1 0 V151  ac -3.418919982455481e-03*Ip1
ISRC151_p2 0 V151  ac 3.793270273764938e-03*Ip2
ISRC151_p3 0 V151  ac -1.010211326719188e-01*Ip3
ISRC151_p4 0 V151  ac -1.814370111925634e-02*Ip4

ISRC152_p1 0 V152  ac 1.302535928216251e-02*Ip1
ISRC152_p2 0 V152  ac 2.330060701532994e-02*Ip2
ISRC152_p3 0 V152  ac -1.870887069950088e-02*Ip3
ISRC152_p4 0 V152  ac 8.090632881334712e-03*Ip4

ISRC153_p1 0 V153  ac -5.404120356653935e-02*Ip1
ISRC153_p2 0 V153  ac -8.482434591828404e-03*Ip2
ISRC153_p3 0 V153  ac -4.500935230526409e-03*Ip3
ISRC153_p4 0 V153  ac 4.563846498229053e-04*Ip4

ISRC154_p1 0 V154  ac -3.617778688371115e-03*Ip1
ISRC154_p2 0 V154  ac 4.901447169333658e-02*Ip2
ISRC154_p3 0 V154  ac -7.408123744690831e-03*Ip3
ISRC154_p4 0 V154  ac 4.867800750030657e-03*Ip4

ISRC155_p1 0 V155  ac 8.676004720543189e-03*Ip1
ISRC155_p2 0 V155  ac 5.760576820892756e-03*Ip2
ISRC155_p3 0 V155  ac 1.779623589151156e-01*Ip3
ISRC155_p4 0 V155  ac -2.783693915067740e-03*Ip4

ISRC156_p1 0 V156  ac 4.449523209069742e-03*Ip1
ISRC156_p2 0 V156  ac -3.377521551058466e-02*Ip2
ISRC156_p3 0 V156  ac -4.444345483182234e-03*Ip3
ISRC156_p4 0 V156  ac -1.944214525530798e-02*Ip4

ISRC157_p1 0 V157  ac -6.166516700186617e-02*Ip1
ISRC157_p2 0 V157  ac 1.451259161489638e-03*Ip2
ISRC157_p3 0 V157  ac 8.151747890732744e-03*Ip3
ISRC157_p4 0 V157  ac -1.196191211392234e-02*Ip4

ISRC158_p1 0 V158  ac 1.693731307477685e-02*Ip1
ISRC158_p2 0 V158  ac -3.447498311778689e-02*Ip2
ISRC158_p3 0 V158  ac 2.016882970319882e-03*Ip3
ISRC158_p4 0 V158  ac -1.709421208676824e-02*Ip4

ISRC159_p1 0 V159  ac 8.562008797333594e-03*Ip1
ISRC159_p2 0 V159  ac -1.127159295936232e-02*Ip2
ISRC159_p3 0 V159  ac -7.840364905489458e-02*Ip3
ISRC159_p4 0 V159  ac -3.047124123512891e-02*Ip4

ISRC160_p1 0 V160  ac 1.271892476086758e-03*Ip1
ISRC160_p2 0 V160  ac 3.174568699169161e-03*Ip2
ISRC160_p3 0 V160  ac 1.056889730379459e-02*Ip3
ISRC160_p4 0 V160  ac 3.819249820225047e-02*Ip4

ISRC161_p1 0 V161  ac -3.228070393673621e-02*Ip1
ISRC161_p2 0 V161  ac 8.530217303083631e-03*Ip2
ISRC161_p3 0 V161  ac -6.552676983492012e-04*Ip3
ISRC161_p4 0 V161  ac -1.017021084071755e-02*Ip4

ISRC162_p1 0 V162  ac 2.341028831769454e-02*Ip1
ISRC162_p2 0 V162  ac -7.346445832212813e-03*Ip2
ISRC162_p3 0 V162  ac -8.449979911116791e-03*Ip3
ISRC162_p4 0 V162  ac -1.826259267429926e-02*Ip4

ISRC163_p1 0 V163  ac 3.022137851023103e-02*Ip1
ISRC163_p2 0 V163  ac 1.223681193345087e-02*Ip2
ISRC163_p3 0 V163  ac 3.349896622374243e-02*Ip3
ISRC163_p4 0 V163  ac -1.159561158543618e-02*Ip4

ISRC164_p1 0 V164  ac 2.136134296487368e-02*Ip1
ISRC164_p2 0 V164  ac 1.376525516633009e-02*Ip2
ISRC164_p3 0 V164  ac -2.902733509396533e-03*Ip3
ISRC164_p4 0 V164  ac -2.942815525117056e-02*Ip4

ISRC165_p1 0 V165  ac -1.950211017956653e-02*Ip1
ISRC165_p2 0 V165  ac -1.803509508288141e-02*Ip2
ISRC165_p3 0 V165  ac -3.541536538193785e-03*Ip3
ISRC165_p4 0 V165  ac -1.675914121943873e-02*Ip4

ISRC166_p1 0 V166  ac 2.947705358270832e-02*Ip1
ISRC166_p2 0 V166  ac -1.439654182783156e-02*Ip2
ISRC166_p3 0 V166  ac 2.751075944413870e-03*Ip3
ISRC166_p4 0 V166  ac -1.404023249025646e-02*Ip4

ISRC167_p1 0 V167  ac 6.875677690116823e-03*Ip1
ISRC167_p2 0 V167  ac -9.892089817770207e-04*Ip2
ISRC167_p3 0 V167  ac -5.313363481338271e-02*Ip3
ISRC167_p4 0 V167  ac -1.810456209994458e-02*Ip4

ISRC168_p1 0 V168  ac 1.673301124156163e-02*Ip1
ISRC168_p2 0 V168  ac 5.391726411068827e-03*Ip2
ISRC168_p3 0 V168  ac 2.147567119673164e-02*Ip3
ISRC168_p4 0 V168  ac 1.994763663332341e-02*Ip4

ISRC169_p1 0 V169  ac 2.453979740547674e-03*Ip1
ISRC169_p2 0 V169  ac -1.366970966241734e-02*Ip2
ISRC169_p3 0 V169  ac -1.715431561174883e-02*Ip3
ISRC169_p4 0 V169  ac -2.099994104613713e-02*Ip4

ISRC170_p1 0 V170  ac -5.418538062632982e-02*Ip1
ISRC170_p2 0 V170  ac 3.833825178252607e-02*Ip2
ISRC170_p3 0 V170  ac -5.022411274056412e-03*Ip3
ISRC170_p4 0 V170  ac -8.895043136002449e-03*Ip4

ISRC171_p1 0 V171  ac -4.476118273911465e-02*Ip1
ISRC171_p2 0 V171  ac -1.221689196874923e-02*Ip2
ISRC171_p3 0 V171  ac 6.581013408062222e-02*Ip3
ISRC171_p4 0 V171  ac -1.481380494429165e-02*Ip4

ISRC172_p1 0 V172  ac -2.999932703651284e-02*Ip1
ISRC172_p2 0 V172  ac -1.917950945115731e-02*Ip2
ISRC172_p3 0 V172  ac -3.082162694671326e-03*Ip3
ISRC172_p4 0 V172  ac 4.422152314720591e-02*Ip4

ISRC173_p1 0 V173  ac -3.949898789305574e-02*Ip1
ISRC173_p2 0 V173  ac 1.852214385526292e-02*Ip2
ISRC173_p3 0 V173  ac 2.114928195067277e-04*Ip3
ISRC173_p4 0 V173  ac 2.148954193432623e-03*Ip4

ISRC174_p1 0 V174  ac 1.171454404938804e-02*Ip1
ISRC174_p2 0 V174  ac -2.632869038937073e-02*Ip2
ISRC174_p3 0 V174  ac -6.278302017946043e-03*Ip3
ISRC174_p4 0 V174  ac 3.777180103607067e-03*Ip4

ISRC175_p1 0 V175  ac 2.910611997290782e-02*Ip1
ISRC175_p2 0 V175  ac -3.758932400358629e-03*Ip2
ISRC175_p3 0 V175  ac -2.792597166999780e-02*Ip3
ISRC175_p4 0 V175  ac 1.520176667938286e-02*Ip4

ISRC176_p1 0 V176  ac 1.944749995903122e-02*Ip1
ISRC176_p2 0 V176  ac -3.949856198861897e-03*Ip2
ISRC176_p3 0 V176  ac 3.459211555914911e-03*Ip3
ISRC176_p4 0 V176  ac -1.134099038612104e-02*Ip4

ISRC177_p1 0 V177  ac -5.385955744358731e-03*Ip1
ISRC177_p2 0 V177  ac -1.161594158928995e-03*Ip2
ISRC177_p3 0 V177  ac -3.366962212314372e-03*Ip3
ISRC177_p4 0 V177  ac -1.025462788412333e-02*Ip4

ISRC178_p1 0 V178  ac 1.280103583443455e-02*Ip1
ISRC178_p2 0 V178  ac -1.158475304106715e-02*Ip2
ISRC178_p3 0 V178  ac 6.416807653214267e-03*Ip3
ISRC178_p4 0 V178  ac 1.164495138025793e-02*Ip4

ISRC179_p1 0 V179  ac 9.955019151620460e-03*Ip1
ISRC179_p2 0 V179  ac 9.101606500778554e-03*Ip2
ISRC179_p3 0 V179  ac 4.239337429737586e-02*Ip3
ISRC179_p4 0 V179  ac 9.253970623143251e-03*Ip4

ISRC180_p1 0 V180  ac 5.453894533977014e-03*Ip1
ISRC180_p2 0 V180  ac 2.054358303946953e-02*Ip2
ISRC180_p3 0 V180  ac -3.274959186339564e-03*Ip3
ISRC180_p4 0 V180  ac -3.485568863846736e-03*Ip4

ISRC181_p1 0 V181  ac 1.286618679067355e-02*Ip1
ISRC181_p2 0 V181  ac -1.391176597013612e-02*Ip2
ISRC181_p3 0 V181  ac -4.789271708817364e-03*Ip3
ISRC181_p4 0 V181  ac 1.667326163335450e-03*Ip4

ISRC182_p1 0 V182  ac -7.694916553845941e-03*Ip1
ISRC182_p2 0 V182  ac -2.717922223389572e-02*Ip2
ISRC182_p3 0 V182  ac 3.976277638822431e-03*Ip3
ISRC182_p4 0 V182  ac 1.511066908091950e-03*Ip4

ISRC183_p1 0 V183  ac -1.261133834552144e-02*Ip1
ISRC183_p2 0 V183  ac 2.700190662464953e-03*Ip2
ISRC183_p3 0 V183  ac -2.022418731398606e-02*Ip3
ISRC183_p4 0 V183  ac 5.276706666305136e-03*Ip4

ISRC184_p1 0 V184  ac -1.122099602366624e-02*Ip1
ISRC184_p2 0 V184  ac 7.100326361685911e-04*Ip2
ISRC184_p3 0 V184  ac 6.874111294410131e-03*Ip3
ISRC184_p4 0 V184  ac 2.788761252548204e-02*Ip4

ISRC185_p1 0 V185  ac -1.712185006096005e-02*Ip1
ISRC185_p2 0 V185  ac 1.289963575847937e-02*Ip2
ISRC185_p3 0 V185  ac 1.890289366070598e-03*Ip3
ISRC185_p4 0 V185  ac 2.198345677967066e-03*Ip4

ISRC186_p1 0 V186  ac 2.102978333730294e-02*Ip1
ISRC186_p2 0 V186  ac -9.521261215054769e-03*Ip2
ISRC186_p3 0 V186  ac -6.490121466933202e-03*Ip3
ISRC186_p4 0 V186  ac 8.472522165518307e-03*Ip4

ISRC187_p1 0 V187  ac 6.162246952581637e-03*Ip1
ISRC187_p2 0 V187  ac -8.481824789532279e-03*Ip2
ISRC187_p3 0 V187  ac -2.189701306483527e-02*Ip3
ISRC187_p4 0 V187  ac 1.894950775530693e-02*Ip4

ISRC188_p1 0 V188  ac -2.174021683779193e-05*Ip1
ISRC188_p2 0 V188  ac -6.215641777665142e-03*Ip2
ISRC188_p3 0 V188  ac 1.145652626325245e-02*Ip3
ISRC188_p4 0 V188  ac -4.099048979391923e-02*Ip4

ISRC189_p1 0 V189  ac 5.411403537001305e-02*Ip1
ISRC189_p2 0 V189  ac 2.304682299766027e-03*Ip2
ISRC189_p3 0 V189  ac -3.371348043229985e-03*Ip3
ISRC189_p4 0 V189  ac 4.685481581649037e-03*Ip4

ISRC190_p1 0 V190  ac -6.408115830514835e-03*Ip1
ISRC190_p2 0 V190  ac -1.901271560435754e-02*Ip2
ISRC190_p3 0 V190  ac -1.174176948020015e-02*Ip3
ISRC190_p4 0 V190  ac -2.627895111441924e-02*Ip4

ISRC191_p1 0 V191  ac -1.887532784624662e-02*Ip1
ISRC191_p2 0 V191  ac 1.256703477676590e-03*Ip2
ISRC191_p3 0 V191  ac -1.249051039108148e-02*Ip3
ISRC191_p4 0 V191  ac -3.697327012155605e-02*Ip4

ISRC192_p1 0 V192  ac -1.015931556660456e-02*Ip1
ISRC192_p2 0 V192  ac 3.787886274584768e-03*Ip2
ISRC192_p3 0 V192  ac -2.360867430702373e-02*Ip3
ISRC192_p4 0 V192  ac 2.897608702587812e-02*Ip4

ISRC193_p1 0 V193  ac -6.760869951021223e-03*Ip1
ISRC193_p2 0 V193  ac 1.848238542232917e-03*Ip2
ISRC193_p3 0 V193  ac -1.082222382895082e-03*Ip3
ISRC193_p4 0 V193  ac 8.527753624809462e-03*Ip4

ISRC194_p1 0 V194  ac -2.657409766995441e-02*Ip1
ISRC194_p2 0 V194  ac -7.041915008944384e-03*Ip2
ISRC194_p3 0 V194  ac 5.224462437293228e-03*Ip3
ISRC194_p4 0 V194  ac -6.584796757252977e-03*Ip4

ISRC195_p1 0 V195  ac -6.142809965468050e-04*Ip1
ISRC195_p2 0 V195  ac 2.337326180408065e-04*Ip2
ISRC195_p3 0 V195  ac 3.176176909773838e-02*Ip3
ISRC195_p4 0 V195  ac 7.317217953623584e-03*Ip4

ISRC196_p1 0 V196  ac -6.550315757960008e-03*Ip1
ISRC196_p2 0 V196  ac 9.140427113656712e-03*Ip2
ISRC196_p3 0 V196  ac -1.728634687174757e-02*Ip3
ISRC196_p4 0 V196  ac -1.899767138801580e-02*Ip4

ISRC197_p1 0 V197  ac -5.853769819391637e-02*Ip1
ISRC197_p2 0 V197  ac 1.092409247643439e-02*Ip2
ISRC197_p3 0 V197  ac -1.023873145954302e-02*Ip3
ISRC197_p4 0 V197  ac 1.017196134626943e-02*Ip4

ISRC198_p1 0 V198  ac 2.741250580113968e-02*Ip1
ISRC198_p2 0 V198  ac 1.301835119676763e-03*Ip2
ISRC198_p3 0 V198  ac -1.661009789440840e-02*Ip3
ISRC198_p4 0 V198  ac -3.328833456810678e-02*Ip4

ISRC199_p1 0 V199  ac 4.581784172651988e-02*Ip1
ISRC199_p2 0 V199  ac 6.877799370912243e-04*Ip2
ISRC199_p3 0 V199  ac 7.564181653188793e-03*Ip3
ISRC199_p4 0 V199  ac -6.364316449912448e-02*Ip4

ISRC200_p1 0 V200  ac 2.235188496521608e-02*Ip1
ISRC200_p2 0 V200  ac 3.708839248587317e-03*Ip2
ISRC200_p3 0 V200  ac 1.031252917511086e-02*Ip3
ISRC200_p4 0 V200  ac 4.955674117142042e-02*Ip4


.ends subckt equivalent_circuit

.end

