* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 
X_11 node_1 0 yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 0 yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 0 yp33
X_34 node_3 node_4 yp34
X_44 node_4 0 yp44
.ends


* Y'11
.subckt yp11 node_1 0
* Branch 0
Rabr0 node_1 netRa0 326.61057146937475
Lbr0 netRa0 netL0 -5.117381476432755e-13
Rbbr0 netL0 0 -2200.7948202195016
Cbr0 netL0 0 -4.80803259443911e-19

* Branch 1
Rabr1 node_1 netRa1 222.5438694403912
Lbr1 netRa1 netL1 -4.3751691175770625e-13
Rbbr1 netL1 0 -2098.2632006837534
Cbr1 netL1 0 -5.869597624192263e-19

* Branch 2
Rabr2 node_1 netRa2 142.47643687284696
Lbr2 netRa2 netL2 -3.4035622605774203e-13
Rbbr2 netL2 0 -1809.8816661859219
Cbr2 netL2 0 -7.700609982977301e-19

* Branch 3
Rabr3 node_1 netRa3 139.02936140865506
Lbr3 netRa3 netL3 -4.901189529746543e-13
Rbbr3 netL3 0 -3075.9955135807954
Cbr3 netL3 0 -5.628061455421911e-19

* Branch 4
Rabr4 node_1 netRa4 -333.6325910193248
Lbr4 netRa4 netL4 -6.452279938227414e-13
Rbbr4 netL4 0 9253.363871967975
Cbr4 netL4 0 -4.347845159698791e-19

* Branch 5
Rabr5 node_1 netRa5 -10369272.719332574
Lbr5 netRa5 netL5 7.245707165438178e-11
Rbbr5 netL5 0 10370990.502703767
Cbr5 netL5 0 6.726862004870602e-25

* Branch 6
Rabr6 node_1 netRa6 193.04356122351857
Lbr6 netRa6 netL6 3.1980595716464953e-13
Rbbr6 netL6 0 -2687.5383501761826
Cbr6 netL6 0 8.6979661357187e-19

* Branch 7
Rabr7 node_1 netRa7 59280.70426488376
Lbr7 netRa7 netL7 2.050982390663445e-12
Rbbr7 netL7 0 -59511.583691876716
Cbr7 netL7 0 5.833565020857678e-22

* Branch 8
Rabr8 node_1 netRa8 -1823.319412902136
Lbr8 netRa8 netL8 -2.154908265435155e-12
Rbbr8 netL8 0 11168.34584993483
Cbr8 netL8 0 -1.1413185330448228e-19

* Branch 9
Rabr9 node_1 netRa9 -5049979.818094138
Lbr9 netRa9 netL9 -4.375765037755529e-11
Rbbr9 netL9 0 5051220.249074346
Cbr9 netL9 0 -1.7161651642923957e-24

* Branch 10
Rabr10 node_1 netRa10 -1144398.2386926573
Lbr10 netRa10 netL10 -4.9088653209177065e-11
Rbbr10 netL10 0 1145805.7453336774
Cbr10 netL10 0 -3.7507957114850805e-23

* Branch 11
Rabr11 node_1 netRa11 20603.887876752688
Lbr11 netRa11 netL11 -4.564807896757151e-12
Rbbr11 netL11 0 -23264.007296597272
Cbr11 netL11 0 -9.441268976294865e-21

* Branch 12
Rabr12 node_1 netRa12 -46736.78260657894
Lbr12 netRa12 netL12 -1.4260555523559178e-11
Rbbr12 netL12 0 49688.63935857222
Cbr12 netL12 0 -6.211598197261353e-21

* Branch 13
Rabr13 node_1 netRa13 -27602.921503384157
Lbr13 netRa13 netL13 1.2919029998912039e-11
Rbbr13 netL13 0 31608.410593550707
Cbr13 netL13 0 1.455668465068999e-20

* Branch 14
Rabr14 node_1 netRa14 -1777.6683249726939
Lbr14 netRa14 netL14 1.4867687118991373e-12
Rbbr14 netL14 0 5515.356095693521
Cbr14 netL14 0 1.472828411570406e-19

* Branch 15
Rabr15 node_1 netRa15 -341.58694345764366
Lbr15 netRa15 netL15 -4.003741529026911e-13
Rbbr15 netL15 0 1650.3563542423067
Cbr15 netL15 0 -7.405338810746267e-19

* Branch 16
Rabr16 node_1 netRa16 124100.31787191561
Lbr16 netRa16 netL16 -1.0956067466657093e-11
Rbbr16 netL16 0 -126650.89549764723
Cbr16 netL16 0 -6.950601382966993e-22

* Branch 17
Rabr17 node_1 netRa17 58.424673291437344
Lbr17 netRa17 netL17 7.594594201968031e-12
Rbbr17 netL17 0 208118.91488447445
Cbr17 netL17 0 1.952157727377674e-19

* Branch 18
Rabr18 node_1 netRa18 52422.7456705161
Lbr18 netRa18 netL18 -1.3528658028606826e-11
Rbbr18 netL18 0 -62078.190715320525
Cbr18 netL18 0 -4.123842069669665e-21

* Branch 19
Rabr19 node_1 netRa19 185083.38969726217
Lbr19 netRa19 netL19 -1.2251434122690868e-11
Rbbr19 netL19 0 -187225.85252011352
Cbr19 netL19 0 -3.5282736784601276e-22

* Branch 20
Rabr20 node_1 netRa20 3787.448115736157
Lbr20 netRa20 netL20 1.8736448074001828e-12
Rbbr20 netL20 0 -6286.08933929191
Cbr20 netL20 0 7.989568336804851e-20

* Branch 21
Rabr21 node_1 netRa21 -1814.4320964489339
Lbr21 netRa21 netL21 3.8052156196048495e-12
Rbbr21 netL21 0 24496.215352854837
Cbr21 netL21 0 8.053778925672055e-20

* Branch 22
Rabr22 node_1 netRa22 -350.3376052935576
Lbr22 netRa22 netL22 4.136531853416352e-12
Rbbr22 netL22 0 107341.26305336072
Cbr22 netL22 0 8.142573760492006e-20

* Branch 23
Rabr23 node_1 netRa23 -276.73200264299714
Lbr23 netRa23 netL23 -8.984847766876161e-13
Rbbr23 netL23 0 2405.497093098574
Cbr23 netL23 0 -1.48704375532406e-18

* Branch 24
Rabr24 node_1 netRa24 17273.91172599369
Lbr24 netRa24 netL24 1.0588943296080566e-11
Rbbr24 netL24 0 -36238.36734656803
Cbr24 netL24 0 1.7195681343448043e-20

* Branch 25
Rabr25 node_1 netRa25 -112.74018590543525
Lbr25 netRa25 netL25 2.040304706451264e-12
Rbbr25 netL25 0 78913.27882042492
Cbr25 netL25 0 1.553991209051218e-19

* Branch 26
Rabr26 node_1 netRa26 461.4730849100955
Lbr26 netRa26 netL26 5.612857163850537e-13
Rbbr26 netL26 0 -2306.750070354589
Cbr26 netL26 0 5.441595157630696e-19

* Branch 27
Rabr27 node_1 netRa27 -25357872.322337534
Lbr27 netRa27 netL27 -1.4252430511442698e-10
Rbbr27 netL27 0 25359981.75436609
Cbr27 netL27 0 -2.216606863487908e-25

* Branch 28
Rabr28 node_1 netRa28 2200.7989479536436
Lbr28 netRa28 netL28 1.5330269510144953e-12
Rbbr28 netL28 0 -4975.040272513325
Cbr28 netL28 0 1.423715958862726e-19

* Branch 29
Rabr29 node_1 netRa29 17262.635173079467
Lbr29 netRa29 netL29 5.4273271111523705e-12
Rbbr29 netL29 0 -19993.918390318202
Cbr29 netL29 0 1.5829936686277327e-20

* Branch 30
Rabr30 node_1 netRa30 520.5020402560228
Lbr30 netRa30 netL30 7.352860081171223e-13
Rbbr30 netL30 0 -2337.9042233404425
Cbr30 netL30 0 6.2247228851436495e-19

* Branch 31
Rabr31 node_1 netRa31 -5918.902399224241
Lbr31 netRa31 netL31 3.2579457027520616e-12
Rbbr31 netL31 0 7137.3293389943765
Cbr31 netL31 0 7.625914175992438e-20

* Branch 32
Rabr32 node_1 netRa32 44853.56595508354
Lbr32 netRa32 netL32 -8.62110198404899e-12
Rbbr32 netL32 0 -48182.467784042165
Cbr32 netL32 0 -3.973646533697732e-21

* Branch 33
Rabr33 node_1 netRa33 14130.481723862635
Lbr33 netRa33 netL33 2.8036112979619105e-12
Rbbr33 netL33 0 -15431.810975632883
Cbr33 netL33 0 1.2907683605629048e-20

* Branch 34
Rabr34 node_1 netRa34 -161.01256982311358
Lbr34 netRa34 netL34 7.826308362812545e-13
Rbbr34 netL34 0 5917.735542519768
Cbr34 netL34 0 7.508164121500441e-19

* Branch 35
Rabr35 node_1 netRa35 31017.49654827111
Lbr35 netRa35 netL35 4.723430356299044e-12
Rbbr35 netL35 0 -32740.463315814537
Cbr35 netL35 0 4.66480860233561e-21

* Branch 36
Rabr36 node_1 netRa36 -2273.5704724688712
Lbr36 netRa36 netL36 -2.803348864585759e-12
Rbbr36 netL36 0 4478.0301923137595
Cbr36 netL36 0 -2.8194038261707407e-19

* Branch 37
Rabr37 node_1 netRa37 51448.13306862744
Lbr37 netRa37 netL37 6.15634444797698e-12
Rbbr37 netL37 0 -52899.589340679224
Cbr37 netL37 0 2.2671406726640717e-21

* Branch 38
Rabr38 node_1 netRa38 700.3628370330492
Lbr38 netRa38 netL38 9.100956924364867e-13
Rbbr38 netL38 0 -2580.3616137400554
Cbr38 netL38 0 5.161446231093987e-19

* Branch 39
Rabr39 node_1 netRa39 -27890.66605062626
Lbr39 netRa39 netL39 7.1908794233927366e-12
Rbbr39 netL39 0 30403.7017298787
Cbr39 netL39 0 8.441243248499901e-21

* Branch 40
Rabr40 node_1 netRa40 -1081.5901546583084
Lbr40 netRa40 netL40 1.068276180864409e-12
Rbbr40 netL40 0 2396.826720344499
Cbr40 netL40 0 4.0516894578742746e-19

* Branch 41
Rabr41 node_1 netRa41 177865.4572332121
Lbr41 netRa41 netL41 -1.594616468664118e-10
Rbbr41 netL41 0 -654752.9508268264
Cbr41 netL41 0 -1.3484694708046026e-21

* Branch 42
Rabr42 node_1 netRa42 3943.5914502195938
Lbr42 netRa42 netL42 3.5514578803468695e-12
Rbbr42 netL42 0 -8265.361280645271
Cbr42 netL42 0 1.10645702705794e-19

* Branch 43
Rabr43 node_1 netRa43 35662.20017553108
Lbr43 netRa43 netL43 6.480447620630142e-12
Rbbr43 netL43 0 -38604.2202882075
Cbr43 netL43 0 4.721624751407409e-21

* Branch 44
Rabr44 node_1 netRa44 224.2770737519292
Lbr44 netRa44 netL44 8.698323702567144e-13
Rbbr44 netL44 0 -5367.716455632127
Cbr44 netL44 0 7.727511832800663e-19

* Branch 45
Rabr45 node_1 netRa45 -446.54374225664026
Lbr45 netRa45 netL45 8.591095508189552e-13
Rbbr45 netL45 0 2880.811467789878
Cbr45 netL45 0 6.471012361299801e-19

* Branch 46
Rabr46 node_1 netRa46 208.69141063802607
Lbr46 netRa46 netL46 9.296485377009404e-13
Rbbr46 netL46 0 -6002.348540280618
Cbr46 netL46 0 8.005268316411923e-19

* Branch 47
Rabr47 node_1 netRa47 2080.578033111982
Lbr47 netRa47 netL47 1.1033096538579315e-12
Rbbr47 netL47 0 -3395.238266815175
Cbr47 netL47 0 1.5751802847288386e-19

* Branch 48
Rabr48 node_1 netRa48 101.40059339867325
Lbr48 netRa48 netL48 7.875093511254381e-13
Rbbr48 netL48 0 -8273.936325682202
Cbr48 netL48 0 1.0701843774940229e-18

* Branch 49
Rabr49 node_1 netRa49 182802.47652732432
Lbr49 netRa49 netL49 2.1483978663561614e-11
Rbbr49 netL49 0 -186479.76279242104
Cbr49 netL49 0 6.314064488193606e-22

* Branch 50
Rabr50 node_1 netRa50 10237.89104255574
Lbr50 netRa50 netL50 1.2109734378165194e-11
Rbbr50 netL50 0 -16510.67837595354
Cbr50 netL50 0 7.297816748530808e-20

* Branch 51
Rabr51 node_1 netRa51 -106610326.97515523
Lbr51 netRa51 netL51 4.900958605546951e-10
Rbbr51 netL51 0 106614983.99205525
Cbr51 netL51 0 4.3115438406904124e-26

* Branch 52
Rabr52 node_1 netRa52 -781.7371189632361
Lbr52 netRa52 netL52 1.2347670226061218e-12
Rbbr52 netL52 0 3437.2189256176594
Cbr52 netL52 0 4.490685894396322e-19

* Branch 53
Rabr53 node_1 netRa53 -254.50325956569117
Lbr53 netRa53 netL53 6.261594846643179e-13
Rbbr53 netL53 0 3397.2347821377243
Cbr53 netL53 0 6.991525960473434e-19

* Branch 54
Rabr54 node_1 netRa54 -751157.6034091921
Lbr54 netRa54 netL54 3.838334509194316e-11
Rbbr54 netL54 0 754343.682771699
Cbr54 netL54 0 6.768944637103557e-23

* Branch 55
Rabr55 node_1 netRa55 12371.213557069053
Lbr55 netRa55 netL55 8.32304830062498e-12
Rbbr55 netL55 0 -19178.99516816798
Cbr55 netL55 0 3.5420660802418403e-20

* Branch 56
Rabr56 node_1 netRa56 -1071894.1614082514
Lbr56 netRa56 netL56 -4.58086909450481e-11
Rbbr56 netL56 0 1074317.5576580246
Cbr56 netL56 0 -3.9803957824100895e-23

* Branch 57
Rabr57 node_1 netRa57 -37133560.51184464
Lbr57 netRa57 netL57 -3.5090762566176124e-10
Rbbr57 netL57 0 37139432.90770302
Cbr57 netL57 0 -2.5447728645126814e-25

* Branch 58
Rabr58 node_1 netRa58 791880.6371782444
Lbr58 netRa58 netL58 -3.267906546732189e-11
Rbbr58 netL58 0 -794213.3367142725
Cbr58 netL58 0 -5.193012445957823e-23

* Branch 59
Rabr59 node_1 netRa59 -15431.678529042287
Lbr59 netRa59 netL59 5.373965898318151e-12
Rbbr59 netL59 0 18199.718750608623
Cbr59 netL59 0 1.9041493085078785e-20

* Branch 60
Rabr60 node_1 netRa60 -87921.69660529992
Lbr60 netRa60 netL60 2.8517469738082418e-11
Rbbr60 netL60 0 117574.69702014008
Cbr60 netL60 0 2.746254234178302e-21

* Branch 61
Rabr61 node_1 netRa61 -2758.6047807833684
Lbr61 netRa61 netL61 5.0768454724818796e-12
Rbbr61 netL61 0 11661.254537811003
Cbr61 netL61 0 1.5389958480575577e-19

* Branch 62
Rabr62 node_1 netRa62 3608.199795103456
Lbr62 netRa62 netL62 1.8275903073134565e-12
Rbbr62 netL62 0 -5734.463257883422
Cbr62 netL62 0 8.894540892214946e-20

* Branch 63
Rabr63 node_1 netRa63 4121.630245053233
Lbr63 netRa63 netL63 1.729159796507296e-12
Rbbr63 netL63 0 -5521.571763599154
Cbr63 netL63 0 7.641741068267683e-20

* Branch 64
Rabr64 node_1 netRa64 -646788.3706456515
Lbr64 netRa64 netL64 -3.439887645277958e-11
Rbbr64 netL64 0 648114.8554668574
Cbr64 netL64 0 -8.211717673884694e-23

* Branch 65
Rabr65 node_1 netRa65 299.30324748757573
Lbr65 netRa65 netL65 5.582858263359128e-13
Rbbr65 netL65 0 -2625.586990924519
Cbr65 netL65 0 7.280445183031181e-19

* Branch 66
Rabr66 node_1 netRa66 -1654.4923263232033
Lbr66 netRa66 netL66 1.1026065535940383e-12
Rbbr66 netL66 0 2975.900939229699
Cbr66 netL66 0 2.220622504806648e-19

* Branch 67
Rabr67 node_1 netRa67 -68613.84445567628
Lbr67 netRa67 netL67 -1.3565745075553794e-11
Rbbr67 netL67 0 70178.7104136802
Cbr67 netL67 0 -2.8242274960729374e-21

* Branch 68
Rabr68 node_1 netRa68 -306.2740252444531
Lbr68 netRa68 netL68 9.822211625529298e-13
Rbbr68 netL68 0 3524.837809453759
Cbr68 netL68 0 8.751824573200287e-19

* Branch 69
Rabr69 node_1 netRa69 27992.472773769015
Lbr69 netRa69 netL69 7.0787139435636524e-12
Rbbr69 netL69 0 -32376.482815303636
Cbr69 netL69 0 7.833553532313383e-21

* Branch 70
Rabr70 node_1 netRa70 -3147.5192021681337
Lbr70 netRa70 netL70 1.7543473916268218e-12
Rbbr70 netL70 0 4264.056312722721
Cbr70 netL70 0 1.2989226420599677e-19

* Branch 71
Rabr71 node_1 netRa71 -288.44971497413894
Lbr71 netRa71 netL71 8.470251659990217e-13
Rbbr71 netL71 0 4740.779220139339
Cbr71 netL71 0 5.994240796988328e-19

* Branch 72
Rabr72 node_1 netRa72 -6843.948324285896
Lbr72 netRa72 netL72 -5.2651218423799e-12
Rbbr72 netL72 0 9261.981052881341
Cbr72 netL72 0 -8.37041562149798e-20

* Branch 73
Rabr73 node_1 netRa73 -91358.42310207002
Lbr73 netRa73 netL73 8.7315590367256e-12
Rbbr73 netL73 0 93157.9989621604
Cbr73 netL73 0 1.0250296646418747e-21

* Branch 74
Rabr74 node_1 netRa74 1009.0203293234782
Lbr74 netRa74 netL74 8.751740485655757e-13
Rbbr74 netL74 0 -2445.340109674062
Cbr74 netL74 0 3.5756484811041946e-19

* Branch 75
Rabr75 node_1 netRa75 73792.98903068753
Lbr75 netRa75 netL75 -3.41089380585003e-11
Rbbr75 netL75 0 -90788.94974292065
Cbr75 netL75 0 -5.0697846830520264e-21

* Branch 76
Rabr76 node_1 netRa76 9053.064921250978
Lbr76 netRa76 netL76 2.8925432643462623e-12
Rbbr76 netL76 0 -10749.399032972593
Cbr76 netL76 0 2.9808919400144065e-20

* Branch 77
Rabr77 node_1 netRa77 -106835.2072796009
Lbr77 netRa77 netL77 1.5267868673151566e-11
Rbbr77 netL77 0 109270.23902604092
Cbr77 netL77 0 1.3061936162179833e-21

* Branch 78
Rabr78 node_1 netRa78 18287.40960103391
Lbr78 netRa78 netL78 -4.298746309609517e-12
Rbbr78 netL78 0 -20431.063398093807
Cbr78 netL78 0 -1.1489690912780342e-20

* Branch 79
Rabr79 node_1 netRa79 -237.03633715170267
Lbr79 netRa79 netL79 7.075827103931839e-13
Rbbr79 netL79 0 1841.6131843369715
Cbr79 netL79 0 1.5946468707612137e-18

* Branch 80
Rabr80 node_1 netRa80 -111542.99288386511
Lbr80 netRa80 netL80 -3.31570626780147e-11
Rbbr80 netL80 0 120285.60306327025
Cbr80 netL80 0 -2.4746091615804093e-21

* Branch 81
Rabr81 node_1 netRa81 504.2350908736966
Lbr81 netRa81 netL81 1.3741467242731394e-12
Rbbr81 netL81 0 -3532.9290118091612
Cbr81 netL81 0 7.805309270774924e-19

* Branch 82
Rabr82 node_1 netRa82 -4798.047606674113
Lbr82 netRa82 netL82 5.150872996261945e-12
Rbbr82 netL82 0 10340.728051307735
Cbr82 netL82 0 1.0334909085792359e-19

* Branch 83
Rabr83 node_1 netRa83 -396.0156383466338
Lbr83 netRa83 netL83 -5.837659281084559e-13
Rbbr83 netL83 0 1056.9463548959234
Cbr83 netL83 0 -1.4029413951994692e-18

* Branch 84
Rabr84 node_1 netRa84 -965.4915139931123
Lbr84 netRa84 netL84 1.992881487019154e-12
Rbbr84 netL84 0 4883.657801284634
Cbr84 netL84 0 4.192427997091575e-19

* Branch 85
Rabr85 node_1 netRa85 3290.800845604087
Lbr85 netRa85 netL85 -2.9265528575280903e-12
Rbbr85 netL85 0 -4785.737917684861
Cbr85 netL85 0 -1.8522882725218438e-19

* Branch 86
Rabr86 node_1 netRa86 605.306536640312
Lbr86 netRa86 netL86 3.1796857930429164e-12
Rbbr86 netL86 0 -14743.321736710837
Cbr86 netL86 0 3.6144468347092254e-19

* Branch 87
Rabr87 node_1 netRa87 -2368.6234665813354
Lbr87 netRa87 netL87 2.701338793533445e-12
Rbbr87 netL87 0 5564.232336150656
Cbr87 netL87 0 2.0445725547614257e-19

* Branch 88
Rabr88 node_1 netRa88 -123.60764123262216
Lbr88 netRa88 netL88 2.0643784155084733e-12
Rbbr88 netL88 0 32223.783434402005
Cbr88 netL88 0 5.177433499631307e-19

* Branch 89
Rabr89 node_1 netRa89 2517.8333510573516
Lbr89 netRa89 netL89 5.53212059185336e-12
Rbbr89 netL89 0 -13076.827986546066
Cbr89 netL89 0 1.6802228317522746e-19

* Branch 90
Rabr90 node_1 netRa90 649.5798299926325
Lbr90 netRa90 netL90 2.077814197826197e-12
Rbbr90 netL90 0 -6622.291026756326
Cbr90 netL90 0 4.832278279627673e-19

* Branch 91
Rabr91 node_1 netRa91 25134.060744343362
Lbr91 netRa91 netL91 5.1894018418779663e-11
Rbbr91 netL91 0 -72554.4943349116
Cbr91 netL91 0 2.848231375565605e-20

* Branch 92
Rabr92 node_1 netRa92 684.5834664431213
Lbr92 netRa92 netL92 -2.257577494057299e-12
Rbbr92 netL92 0 -4614.456481010133
Cbr92 netL92 0 -7.129723208911178e-19

* Branch 93
Rabr93 node_1 netRa93 1085.0906909213165
Lbr93 netRa93 netL93 -2.5099113693286366e-12
Rbbr93 netL93 0 -4265.982360849354
Cbr93 netL93 0 -5.405153445130858e-19

* Branch 94
Rabr94 node_1 netRa94 513.5716353140076
Lbr94 netRa94 netL94 -3.2609705988202728e-12
Rbbr94 netL94 0 -10846.661169576775
Cbr94 netL94 0 -5.791392936183597e-19

* Branch 95
Rabr95 node_1 netRa95 242.5879497903749
Lbr95 netRa95 netL95 -3.650435865172915e-12
Rbbr95 netL95 0 -25704.5808776694
Cbr95 netL95 0 -5.667624749194518e-19

* Branch 96
Rabr96 node_1 netRa96 254.19377071019727
Lbr96 netRa96 netL96 -3.6715152831432734e-12
Rbbr96 netL96 0 -23567.207800566244
Cbr96 netL96 0 -5.896912635294459e-19

* Branch 97
Rabr97 node_1 netRa97 7990.031200947222
Lbr97 netRa97 netL97 -1.7856971234302524e-12
Rbbr97 netL97 0 -9040.740601949528
Cbr97 netL97 0 -2.457689397823807e-20

* Branch 98
Rabr98 node_1 netRa98 -11539.073688878661
Lbr98 netRa98 netL98 1.0917132717723217e-11
Rbbr98 netL98 0 18280.933088231912
Cbr98 netL98 0 5.0103322436264375e-20

* Branch 99
Rabr99 node_1 netRa99 226.37305748538049
Lbr99 netRa99 netL99 -3.9366613323596333e-13
Rbbr99 netL99 0 -1789.79745392947
Cbr99 netL99 0 -6.341640074570584e-19

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 169808951.3172598
Lbr0 netRa0 netL0 4.479281388528496e-09
Rbbr0 netL0 node_2 -170001222.2893393
Cbr0 netL0 node_2 1.5785156359682692e-25

* Branch 1
Rabr1 node_1 netRa1 166567623.82609943
Lbr1 netRa1 netL1 4.143678367817688e-09
Rbbr1 netL1 node_2 -166738222.78163382
Cbr1 netL1 node_2 1.5153107916040185e-25

* Branch 2
Rabr2 node_1 netRa2 915730642.8564659
Lbr2 netRa2 netL2 -8.82286344127248e-09
Rbbr2 netL2 node_2 -915871159.0443059
Cbr2 netL2 node_2 -1.046296076086981e-26

* Branch 3
Rabr3 node_1 netRa3 26281771.411704186
Lbr3 netRa3 netL3 -1.3347204745095725e-09
Rbbr3 netL3 node_2 -26394251.011932455
Cbr3 netL3 node_2 -1.8774857987817946e-24

* Branch 4
Rabr4 node_1 netRa4 2044122.4010606175
Lbr4 netRa4 netL4 -3.2398116683481204e-10
Rbbr4 netL4 node_2 -2127915.285887631
Cbr4 netL4 node_2 -7.052441502798898e-23

* Branch 5
Rabr5 node_1 netRa5 301064.8942012801
Lbr5 netRa5 netL5 -9.342122306335802e-11
Rbbr5 netL5 node_2 -353435.41712570866
Cbr5 netL5 node_2 -8.647204443363676e-22

* Branch 6
Rabr6 node_1 netRa6 10210.58776740934
Lbr6 netRa6 netL6 7.035751259769162e-12
Rbbr6 netL6 node_2 -25908.340265988092
Cbr6 netL6 node_2 2.6950308530394606e-20

* Branch 7
Rabr7 node_1 netRa7 -1263.1804462822445
Lbr7 netRa7 netL7 3.994888457253101e-12
Rbbr7 netL7 node_2 39761.88426214638
Cbr7 netL7 node_2 7.510353279260003e-20

* Branch 8
Rabr8 node_1 netRa8 122643.86239589774
Lbr8 netRa8 netL8 -6.805075055557287e-11
Rbbr8 netL8 node_2 -183730.59225280964
Cbr8 netL8 node_2 -2.990715772655852e-21

* Branch 9
Rabr9 node_1 netRa9 8999.744476563445
Lbr9 netRa9 netL9 8.629773519041832e-12
Rbbr9 netL9 node_2 -34699.02241881427
Cbr9 netL9 node_2 2.8063579356263115e-20

* Branch 10
Rabr10 node_1 netRa10 112982.94352813651
Lbr10 netRa10 netL10 -4.771068353870332e-11
Rbbr10 netL10 node_2 -124237.3924518753
Cbr10 netL10 node_2 -3.37921506156419e-21

* Branch 11
Rabr11 node_1 netRa11 3269.6187604203474
Lbr11 netRa11 netL11 -1.3260043096387568e-11
Rbbr11 netL11 node_2 -28792.64717622359
Cbr11 netL11 node_2 -1.3335899670717273e-19

* Branch 12
Rabr12 node_1 netRa12 31645.927936333115
Lbr12 netRa12 netL12 2.246594390080263e-11
Rbbr12 netL12 node_2 -39421.03699795083
Cbr12 netL12 node_2 1.818387394023412e-20

* Branch 13
Rabr13 node_1 netRa13 -927.7944103522165
Lbr13 netRa13 netL13 1.279649273006556e-11
Rbbr13 netL13 node_2 81425.81509118291
Cbr13 netL13 node_2 1.4266398954093212e-19

* Branch 14
Rabr14 node_1 netRa14 655.2386663446703
Lbr14 netRa14 netL14 3.8236637571354825e-12
Rbbr14 netL14 node_2 -80332.14200894648
Cbr14 netL14 node_2 7.879979583814671e-20

* Branch 15
Rabr15 node_1 netRa15 -195949921.59082758
Lbr15 netRa15 netL15 1.9089064934523897e-09
Rbbr15 netL15 node_2 195959603.86798024
Cbr15 netL15 node_2 4.9706879918585425e-26

* Branch 16
Rabr16 node_1 netRa16 1676.3765517208458
Lbr16 netRa16 netL16 1.0803458841467192e-11
Rbbr16 netL16 node_2 -36888.99787875653
Cbr16 netL16 node_2 1.9067745790386845e-19

* Branch 17
Rabr17 node_1 netRa17 -16219.595809083636
Lbr17 netRa17 netL17 1.990277753660919e-11
Rbbr17 netL17 node_2 26913.200035857422
Cbr17 netL17 node_2 4.4880698644796613e-20

* Branch 18
Rabr18 node_1 netRa18 -3881.272721354793
Lbr18 netRa18 netL18 1.8605635982814637e-11
Rbbr18 netL18 node_2 54796.41084102967
Cbr18 netL18 node_2 8.247614342758465e-20

* Branch 19
Rabr19 node_1 netRa19 -49854.89670140304
Lbr19 netRa19 netL19 -4.626871109637935e-11
Rbbr19 netL19 node_2 68397.04503312052
Cbr19 netL19 node_2 -1.3725264738069545e-20

* Branch 20
Rabr20 node_1 netRa20 -6304.067354620804
Lbr20 netRa20 netL20 -1.1228370931002218e-11
Rbbr20 netL20 node_2 18227.252789362472
Cbr20 netL20 node_2 -9.980430074770153e-20

* Branch 21
Rabr21 node_1 netRa21 820.4538358075656
Lbr21 netRa21 netL21 3.825101781539649e-12
Rbbr21 netL21 node_2 -64139.70434237396
Cbr21 netL21 node_2 7.683424745744214e-20

* Branch 22
Rabr22 node_1 netRa22 329272.28737271944
Lbr22 netRa22 netL22 -9.023785045666763e-11
Rbbr22 netL22 node_2 -376756.54171136324
Cbr22 netL22 node_2 -7.251142026678774e-22

* Branch 23
Rabr23 node_1 netRa23 40243.91076986043
Lbr23 netRa23 netL23 -3.808469228290112e-11
Rbbr23 netL23 node_2 -70768.13492415102
Cbr23 netL23 node_2 -1.3229497748314076e-20

* Branch 24
Rabr24 node_1 netRa24 27719.503749673357
Lbr24 netRa24 netL24 1.1559004557021956e-11
Rbbr24 netL24 node_2 -41745.533788597895
Cbr24 netL24 node_2 1.003368419420715e-20

* Branch 25
Rabr25 node_1 netRa25 -17228.712771515755
Lbr25 netRa25 netL25 -4.735444978717804e-11
Rbbr25 netL25 node_2 145395.28270625524
Cbr25 netL25 node_2 -1.9467849331751542e-20

* Branch 26
Rabr26 node_1 netRa26 -18657.646716775143
Lbr26 netRa26 netL26 -3.6253820793073687e-11
Rbbr26 netL26 node_2 69684.96690168076
Cbr26 netL26 node_2 -2.8417158937973924e-20

* Branch 27
Rabr27 node_1 netRa27 -11752.727985018813
Lbr27 netRa27 netL27 -2.9073677540468922e-11
Rbbr27 netL27 node_2 61536.61027587581
Cbr27 netL27 node_2 -4.1150107387507435e-20

* Branch 28
Rabr28 node_1 netRa28 413.43777761521534
Lbr28 netRa28 netL28 4.007937728751795e-12
Rbbr28 netL28 node_2 -146278.30865559753
Cbr28 netL28 node_2 7.260594561198036e-20

* Branch 29
Rabr29 node_1 netRa29 -27569.34198560533
Lbr29 netRa29 netL29 -3.2454309317462925e-11
Rbbr29 netL29 node_2 52530.40106046663
Cbr29 netL29 node_2 -2.2640698508745934e-20

* Branch 30
Rabr30 node_1 netRa30 75923.5481053151
Lbr30 netRa30 netL30 -5.886382074139075e-11
Rbbr30 netL30 node_2 -144505.08231729036
Cbr30 netL30 node_2 -5.3322206823999756e-21

* Branch 31
Rabr31 node_1 netRa31 1248320.263938297
Lbr31 netRa31 netL31 9.761587607365594e-11
Rbbr31 netL31 node_2 -1268507.3351136844
Cbr31 netL31 node_2 6.168308816069327e-23

* Branch 32
Rabr32 node_1 netRa32 4879.29797383358
Lbr32 netRa32 netL32 4.403436442814524e-12
Rbbr32 netL32 node_2 -17452.66975096981
Cbr32 netL32 node_2 5.20617181215237e-20

* Branch 33
Rabr33 node_1 netRa33 -1260.7097765759163
Lbr33 netRa33 netL33 3.46278011655018e-12
Rbbr33 netL33 node_2 33909.73540521138
Cbr33 netL33 node_2 7.94966092591838e-20

* Branch 34
Rabr34 node_1 netRa34 3803.3215568091873
Lbr34 netRa34 netL34 3.9118638062161145e-12
Rbbr34 netL34 node_2 -16289.485670563245
Cbr34 netL34 node_2 6.355780405488456e-20

* Branch 35
Rabr35 node_1 netRa35 -29975.40003144745
Lbr35 netRa35 netL35 -4.6663012547127104e-11
Rbbr35 netL35 node_2 107994.51811109913
Cbr35 netL35 node_2 -1.4558832625976287e-20

* Branch 36
Rabr36 node_1 netRa36 47723.806692038655
Lbr36 netRa36 netL36 -5.324874531301988e-11
Rbbr36 netL36 node_2 -130576.54544776872
Cbr36 netL36 node_2 -8.485046590092343e-21

* Branch 37
Rabr37 node_1 netRa37 -2193983.6095282575
Lbr37 netRa37 netL37 -1.74127348395648e-10
Rbbr37 netL37 node_2 2204733.70513981
Cbr37 netL37 node_2 -3.6015196065789706e-23

* Branch 38
Rabr38 node_1 netRa38 23418.35527261634
Lbr38 netRa38 netL38 -4.610330880186845e-11
Rbbr38 netL38 node_2 -139029.3071975478
Cbr38 netL38 node_2 -1.4015834147168468e-20

* Branch 39
Rabr39 node_1 netRa39 1454952.410589981
Lbr39 netRa39 netL39 -1.509607694069948e-10
Rbbr39 netL39 node_2 -1490215.0975636337
Cbr39 netL39 node_2 -6.958762999211678e-23

* Branch 40
Rabr40 node_1 netRa40 733497.515103407
Lbr40 netRa40 netL40 -1.161555416444788e-10
Rbbr40 netL40 node_2 -772761.4234045654
Cbr40 netL40 node_2 -2.047603418118933e-22

* Branch 41
Rabr41 node_1 netRa41 24682002.13966927
Lbr41 netRa41 netL41 4.924545871774469e-10
Rbbr41 netL41 node_2 -24706972.072812617
Cbr41 netL41 node_2 8.076248404590255e-25

* Branch 42
Rabr42 node_1 netRa42 28987.111632984546
Lbr42 netRa42 netL42 1.322231604298157e-11
Rbbr42 netL42 node_2 -45438.890078541524
Cbr42 netL42 node_2 1.0061103363983317e-20

* Branch 43
Rabr43 node_1 netRa43 -18821.780189149827
Lbr43 netRa43 netL43 1.3652128125011883e-11
Rbbr43 netL43 node_2 27460.529124832246
Cbr43 netL43 node_2 2.6335264562996668e-20

* Branch 44
Rabr44 node_1 netRa44 3672.0796058433566
Lbr44 netRa44 netL44 8.499265097784467e-12
Rbbr44 netL44 node_2 -22308.64080854959
Cbr44 netL44 node_2 1.0473450549645599e-19

* Branch 45
Rabr45 node_1 netRa45 171998.16285050262
Lbr45 netRa45 netL45 -7.33960457959008e-11
Rbbr45 netL45 node_2 -226448.19214846747
Cbr45 netL45 node_2 -1.8812888584332258e-21

* Branch 46
Rabr46 node_1 netRa46 9524.609426221443
Lbr46 netRa46 netL46 1.1107110734616982e-11
Rbbr46 netL46 node_2 -20376.047584795782
Cbr46 netL46 node_2 5.744747352658171e-20

* Branch 47
Rabr47 node_1 netRa47 197921.08977372074
Lbr47 netRa47 netL47 -4.038347914013548e-11
Rbbr47 netL47 node_2 -204181.6456184265
Cbr47 netL47 node_2 -9.98739808213303e-22

* Branch 48
Rabr48 node_1 netRa48 3339926.1212129835
Lbr48 netRa48 netL48 -2.1006869118479978e-10
Rbbr48 netL48 node_2 -3371117.2021075683
Cbr48 netL48 node_2 -1.865424598400655e-23

* Branch 49
Rabr49 node_1 netRa49 -5554.423747770516
Lbr49 netRa49 netL49 1.4439355630470783e-11
Rbbr49 netL49 node_2 39364.084233649315
Cbr49 netL49 node_2 6.563587969435999e-20

* Branch 50
Rabr50 node_1 netRa50 -1215.3765694825559
Lbr50 netRa50 netL50 9.991875431828072e-12
Rbbr50 netL50 node_2 85685.59390981618
Cbr50 netL50 node_2 9.415325047117502e-20

* Branch 51
Rabr51 node_1 netRa51 -494.37419759804607
Lbr51 netRa51 netL51 1.7819116577261115e-11
Rbbr51 netL51 node_2 478763.16502422397
Cbr51 netL51 node_2 6.962059979107642e-20

* Branch 52
Rabr52 node_1 netRa52 -43588.526296664386
Lbr52 netRa52 netL52 1.9023315306397393e-11
Rbbr52 netL52 node_2 51710.295420965
Cbr52 netL52 node_2 8.43421368384126e-21

* Branch 53
Rabr53 node_1 netRa53 3655.4338964957974
Lbr53 netRa53 netL53 -4.080133881661546e-11
Rbbr53 netL53 node_2 -532967.7572676779
Cbr53 netL53 node_2 -2.0664633716613762e-20

* Branch 54
Rabr54 node_1 netRa54 156291.08506668426
Lbr54 netRa54 netL54 -7.874120346110147e-11
Rbbr54 netL54 node_2 -181050.41480188604
Cbr54 netL54 node_2 -2.781183192551519e-21

* Branch 55
Rabr55 node_1 netRa55 -55044.80947021395
Lbr55 netRa55 netL55 2.959572672936781e-11
Rbbr55 netL55 node_2 71149.96909287352
Cbr55 netL55 node_2 7.55347430538843e-21

* Branch 56
Rabr56 node_1 netRa56 67045.39755428776
Lbr56 netRa56 netL56 -5.380647789634709e-11
Rbbr56 netL56 node_2 -97811.53652859855
Cbr56 netL56 node_2 -8.204274286122315e-21

* Branch 57
Rabr57 node_1 netRa57 -21533.838556288636
Lbr57 netRa57 netL57 -4.42640981081652e-11
Rbbr57 netL57 node_2 80926.43644671506
Cbr57 netL57 node_2 -2.5403637782670502e-20

* Branch 58
Rabr58 node_1 netRa58 -1925.4216977869382
Lbr58 netRa58 netL58 -4.507316940334605e-11
Rbbr58 netL58 node_2 722442.127296396
Cbr58 netL58 node_2 -3.243970899831925e-20

* Branch 59
Rabr59 node_1 netRa59 -2094563.8374034017
Lbr59 netRa59 netL59 1.4608317217593601e-10
Rbbr59 netL59 node_2 2105633.4265085654
Cbr59 netL59 node_2 3.3122474823535196e-23

* Branch 60
Rabr60 node_1 netRa60 70308.94308526626
Lbr60 netRa60 netL60 1.5162206753120544e-11
Rbbr60 netL60 node_2 -79209.73792622656
Cbr60 netL60 node_2 2.7225504680284423e-21

* Branch 61
Rabr61 node_1 netRa61 1817172.6660893685
Lbr61 netRa61 netL61 1.7807701351593705e-10
Rbbr61 netL61 node_2 -1858767.4721108952
Cbr61 netL61 node_2 5.272142762374596e-23

* Branch 62
Rabr62 node_1 netRa62 142263.23170495036
Lbr62 netRa62 netL62 2.71802237714685e-11
Rbbr62 netL62 node_2 -157039.90807843968
Cbr62 netL62 node_2 1.2166103575125199e-21

* Branch 63
Rabr63 node_1 netRa63 696650.5193133559
Lbr63 netRa63 netL63 1.3568708850122396e-10
Rbbr63 netL63 node_2 -758194.2219739226
Cbr63 netL63 node_2 2.5689068976485382e-22

* Branch 64
Rabr64 node_1 netRa64 569783.9610679746
Lbr64 netRa64 netL64 1.4263373832247316e-10
Rbbr64 netL64 node_2 -645294.924186664
Cbr64 netL64 node_2 3.879370978796793e-22

* Branch 65
Rabr65 node_1 netRa65 505140.79082142893
Lbr65 netRa65 netL65 1.0237292915125013e-10
Rbbr65 netL65 node_2 -556923.1649724812
Cbr65 netL65 node_2 3.639015099124991e-22

* Branch 66
Rabr66 node_1 netRa66 497898.9054102991
Lbr66 netRa66 netL66 1.3372621539114195e-10
Rbbr66 netL66 node_2 -571992.0168950477
Cbr66 netL66 node_2 4.695632178880182e-22

* Branch 67
Rabr67 node_1 netRa67 469608.03644676716
Lbr67 netRa67 netL67 1.3135463016286327e-10
Rbbr67 netL67 node_2 -541660.669590043
Cbr67 netL67 node_2 5.164064197953828e-22

* Branch 68
Rabr68 node_1 netRa68 345388.4666085766
Lbr68 netRa68 netL68 1.1631594462691056e-10
Rbbr68 netL68 node_2 -420252.28372208046
Cbr68 netL68 node_2 8.013688035493409e-22

* Branch 69
Rabr69 node_1 netRa69 444976.7878646631
Lbr69 netRa69 netL69 1.2630159757738905e-10
Rbbr69 netL69 node_2 -517094.82816912804
Cbr69 netL69 node_2 5.489221080600681e-22

* Branch 70
Rabr70 node_1 netRa70 367325.95956712397
Lbr70 netRa70 netL70 1.2827398726024627e-10
Rbbr70 netL70 node_2 -450727.4010907072
Cbr70 netL70 node_2 7.747915193201315e-22

* Branch 71
Rabr71 node_1 netRa71 470405.49477590085
Lbr71 netRa71 netL71 1.2657434178912043e-10
Rbbr71 netL71 node_2 -546032.6733609517
Cbr71 netL71 node_2 4.9279226981038345e-22

* Branch 72
Rabr72 node_1 netRa72 278368.35495924397
Lbr72 netRa72 netL72 1.2146198532922674e-10
Rbbr72 netL72 node_2 -369410.0523224699
Cbr72 netL72 node_2 1.181209518558202e-21

* Branch 73
Rabr73 node_1 netRa73 249430.3288380024
Lbr73 netRa73 netL73 1.1611479897492592e-10
Rbbr73 netL73 node_2 -339759.1695799241
Cbr73 netL73 node_2 1.3701987677885856e-21

* Branch 74
Rabr74 node_1 netRa74 299076.1145213708
Lbr74 netRa74 netL74 1.1545747139373964e-10
Rbbr74 netL74 node_2 -377752.9834601814
Cbr74 netL74 node_2 1.0219898973018323e-21

* Branch 75
Rabr75 node_1 netRa75 281664.5814184761
Lbr75 netRa75 netL75 1.1247316048472426e-10
Rbbr75 netL75 node_2 -363100.19393305876
Cbr75 netL75 node_2 1.0997776272007693e-21

* Branch 76
Rabr76 node_1 netRa76 461503.7212830943
Lbr76 netRa76 netL76 1.0529089262417924e-10
Rbbr76 netL76 node_2 -516134.4463764065
Cbr76 netL76 node_2 4.420395912225574e-22

* Branch 77
Rabr77 node_1 netRa77 182269.86610622387
Lbr77 netRa77 netL77 1.0427112687184858e-10
Rbbr77 netL77 node_2 -279203.9370061047
Cbr77 netL77 node_2 2.0490348110424063e-21

* Branch 78
Rabr78 node_1 netRa78 172750.41673129305
Lbr78 netRa78 netL78 1.0822883242139893e-10
Rbbr78 netL78 node_2 -276817.84449023067
Cbr78 netL78 node_2 2.26336162023969e-21

* Branch 79
Rabr79 node_1 netRa79 170468.94112029494
Lbr79 netRa79 netL79 1.0471184960973877e-10
Rbbr79 netL79 node_2 -272068.62439975806
Cbr79 netL79 node_2 2.257855090165868e-21

* Branch 80
Rabr80 node_1 netRa80 391004.5748247919
Lbr80 netRa80 netL80 1.0996868485982959e-10
Rbbr80 netL80 node_2 -458036.0857910417
Cbr80 netL80 node_2 6.140430403145721e-22

* Branch 81
Rabr81 node_1 netRa81 120773.64516987675
Lbr81 netRa81 netL81 1.0181043120552204e-10
Rbbr81 netL81 node_2 -248711.82078644857
Cbr81 netL81 node_2 3.389690663128025e-21

* Branch 82
Rabr82 node_1 netRa82 34637.11198874462
Lbr82 netRa82 netL82 1.1838424156258652e-10
Rbbr82 netL82 node_2 -552525.8602847754
Cbr82 netL82 node_2 6.18798861665738e-21

* Branch 83
Rabr83 node_1 netRa83 103741.02135650282
Lbr83 netRa83 netL83 1.029006863821528e-10
Rbbr83 netL83 node_2 -247076.12014950125
Cbr83 netL83 node_2 4.014953396869999e-21

* Branch 84
Rabr84 node_1 netRa84 120635.42303489674
Lbr84 netRa84 netL84 1.0518290745508983e-10
Rbbr84 netL84 node_2 -253355.34892135483
Cbr84 netL84 node_2 3.4417452584885105e-21

* Branch 85
Rabr85 node_1 netRa85 358566.02209344285
Lbr85 netRa85 netL85 8.657087537898374e-11
Rbbr85 netL85 node_2 -409554.46454844833
Cbr85 netL85 node_2 5.895245374779144e-22

* Branch 86
Rabr86 node_1 netRa86 230900.9050487869
Lbr86 netRa86 netL86 6.258620674185588e-11
Rbbr86 netL86 node_2 -275185.9311273105
Cbr86 netL86 node_2 9.850083835177842e-22

* Branch 87
Rabr87 node_1 netRa87 66403.91973981033
Lbr87 netRa87 netL87 9.940916156868916e-11
Rbbr87 netL87 node_2 -269127.4804362036
Cbr87 netL87 node_2 5.563510153238901e-21

* Branch 88
Rabr88 node_1 netRa88 49624.24527637453
Lbr88 netRa88 netL88 1.0463544461967691e-10
Rbbr88 netL88 node_2 -341018.1769220511
Cbr88 netL88 node_2 6.184637743125271e-21

* Branch 89
Rabr89 node_1 netRa89 185864.93597849153
Lbr89 netRa89 netL89 4.884676492549557e-11
Rbbr89 netL89 node_2 -218631.55100096483
Cbr89 netL89 node_2 1.2021017380585217e-21

* Branch 90
Rabr90 node_1 netRa90 -582662.3365884358
Lbr90 netRa90 netL90 1.144262794505781e-10
Rbbr90 netL90 node_2 607897.4695361658
Cbr90 netL90 node_2 3.2304765294548474e-22

* Branch 91
Rabr91 node_1 netRa91 -22903.987931986325
Lbr91 netRa91 netL91 8.964578091899908e-11
Rbbr91 netL91 node_2 457472.68081011437
Cbr91 netL91 node_2 8.55062417106208e-21

* Branch 92
Rabr92 node_1 netRa92 -76758.80866932744
Lbr92 netRa92 netL92 9.075532406452258e-11
Rbbr92 netL92 node_2 205468.5502649473
Cbr92 netL92 node_2 5.753329639119494e-21

* Branch 93
Rabr93 node_1 netRa93 -107832.33828373947
Lbr93 netRa93 netL93 6.728016879799907e-11
Rbbr93 netL93 node_2 156559.87129847123
Cbr93 netL93 node_2 3.984730942527187e-21

* Branch 94
Rabr94 node_1 netRa94 101998.85200976716
Lbr94 netRa94 netL94 2.6787731417197277e-11
Rbbr94 netL94 node_2 -121599.11376889351
Cbr94 netL94 node_2 2.1599623755962097e-21

* Branch 95
Rabr95 node_1 netRa95 50602.1679832866
Lbr95 netRa95 netL95 2.2825560953973994e-11
Rbbr95 netL95 node_2 -78078.85706919357
Cbr95 netL95 node_2 5.778244000067135e-21

* Branch 96
Rabr96 node_1 netRa96 21033.581053614515
Lbr96 netRa96 netL96 7.467389058905235e-12
Rbbr96 netL96 node_2 -28727.13090132454
Cbr96 netL96 node_2 1.2360945572251246e-20

* Branch 97
Rabr97 node_1 netRa97 15438.898116978904
Lbr97 netRa97 netL97 6.698646121863135e-12
Rbbr97 netL97 node_2 -24055.4976234382
Cbr97 netL97 node_2 1.8045886838914422e-20

* Branch 98
Rabr98 node_1 netRa98 7551.630821584635
Lbr98 netRa98 netL98 3.967114292637416e-12
Rbbr98 netL98 node_2 -13848.85396597243
Cbr98 netL98 node_2 3.7969804382014474e-20

* Branch 99
Rabr99 node_1 netRa99 -6723.847335513704
Lbr99 netRa99 netL99 3.672197636346571e-12
Rbbr99 netL99 node_2 13875.869753924002
Cbr99 netL99 node_2 3.931993418722382e-20

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 -71466284.67849602
Lbr0 netRa0 netL0 1.408029580426109e-09
Rbbr0 netL0 node_3 71554155.40209906
Cbr0 netL0 node_3 2.7507132404231944e-25

* Branch 1
Rabr1 node_1 netRa1 -4465735.171256416
Lbr1 netRa1 netL1 5.431159317019115e-10
Rbbr1 netL1 node_3 4640098.675646492
Cbr1 netL1 node_3 2.6072821106784893e-23

* Branch 2
Rabr2 node_1 netRa2 -12165066.259611245
Lbr2 netRa2 netL2 6.090991974469992e-10
Rbbr2 netL2 node_3 12260112.658437086
Cbr2 netL2 node_3 4.075311064111188e-24

* Branch 3
Rabr3 node_1 netRa3 -48057510.06493399
Lbr3 netRa3 netL3 1.0819460764999927e-09
Rbbr3 netL3 node_3 48135978.6770833
Cbr3 netL3 node_3 4.672870093347104e-25

* Branch 4
Rabr4 node_1 netRa4 -4256180.434532034
Lbr4 netRa4 netL4 5.114491953046574e-10
Rbbr4 netL4 node_3 4421651.188006404
Cbr4 netL4 node_3 2.705320470378721e-23

* Branch 5
Rabr5 node_1 netRa5 -3340862.112605553
Lbr5 netRa5 netL5 3.678171028337995e-10
Rbbr5 netL5 node_3 3461505.2488635876
Cbr5 netL5 node_3 3.171436406310371e-23

* Branch 6
Rabr6 node_1 netRa6 -2568100.901726931
Lbr6 netRa6 netL6 5.703309080003867e-10
Rbbr6 netL6 node_3 2836933.078490669
Cbr6 netL6 node_3 7.784604443148855e-23

* Branch 7
Rabr7 node_1 netRa7 -3274722.8154639457
Lbr7 netRa7 netL7 4.4899079512835935e-10
Rbbr7 netL7 node_3 3440574.623742548
Cbr7 netL7 node_3 3.9714783719156414e-23

* Branch 8
Rabr8 node_1 netRa8 -2446533.782405937
Lbr8 netRa8 netL8 5.668958098834992e-10
Rbbr8 netL8 node_3 2722250.917312104
Cbr8 netL8 node_3 8.476451654919826e-23

* Branch 9
Rabr9 node_1 netRa9 -2676232.556039192
Lbr9 netRa9 netL9 4.782018313492777e-10
Rbbr9 netL9 node_3 2885197.008050948
Cbr9 netL9 node_3 6.173460592074374e-23

* Branch 10
Rabr10 node_1 netRa10 -1745806.9912464689
Lbr10 netRa10 netL10 9.250978057804966e-10
Rbbr10 netL10 node_3 2218379.5197115717
Cbr10 netL10 node_3 2.3666212732985365e-22

* Branch 11
Rabr11 node_1 netRa11 -1856030.7625974868
Lbr11 netRa11 netL11 9.024703602742539e-10
Rbbr11 netL11 node_3 2314625.5289234784
Cbr11 netL11 node_3 2.0830767866945542e-22

* Branch 12
Rabr12 node_1 netRa12 -1632845.7700964648
Lbr12 netRa12 netL12 9.465193258650081e-10
Rbbr12 netL12 node_3 2118973.7953784396
Cbr12 netL12 node_3 2.708354912528185e-22

* Branch 13
Rabr13 node_1 netRa13 -1518469.2015472413
Lbr13 netRa13 netL13 9.667919195871672e-10
Rbbr13 netL13 node_3 2017718.1680714998
Cbr13 netL13 node_3 3.1215050913117353e-22

* Branch 14
Rabr14 node_1 netRa14 -7264.0115889568715
Lbr14 netRa14 netL14 -6.019344868450137e-11
Rbbr14 netL14 node_3 1993921.8225462853
Cbr14 netL14 node_3 -4.82666806065027e-21

* Branch 15
Rabr15 node_1 netRa15 -1963384.0645567526
Lbr15 netRa15 netL15 8.776125613233533e-10
Rbbr15 netL15 node_3 2407325.136341325
Cbr15 netL15 node_3 1.8434389802322813e-22

* Branch 16
Rabr16 node_1 netRa16 -2155930.219028675
Lbr16 netRa16 netL16 8.243902598594174e-10
Rbbr16 netL16 node_3 2569621.8213103125
Cbr16 netL16 node_3 1.4791169121651026e-22

* Branch 17
Rabr17 node_1 netRa17 -2278762.774697587
Lbr17 netRa17 netL17 8.013641602867822e-10
Rbbr17 netL17 node_3 2675808.0435234685
Cbr17 netL17 node_3 1.3071667031638864e-22

* Branch 18
Rabr18 node_1 netRa18 -1293313.215466186
Lbr18 netRa18 netL18 1.0056514069175816e-09
Rbbr18 netL18 node_3 1817290.7726447724
Cbr18 netL18 node_3 4.22865281941623e-22

* Branch 19
Rabr19 node_1 netRa19 -2061911.7796260316
Lbr19 netRa19 netL19 8.524681749761172e-10
Rbbr19 netL19 node_3 2491613.7277693534
Cbr19 netL19 node_3 1.649093617973969e-22

* Branch 20
Rabr20 node_1 netRa20 -1404878.4720714544
Lbr20 netRa20 netL20 9.87096360504648e-10
Rbbr20 netL20 node_3 1917686.3744044886
Cbr20 netL20 node_3 3.6259273416953666e-22

* Branch 21
Rabr21 node_1 netRa21 -1181026.1801839187
Lbr21 netRa21 netL21 1.0234661631933664e-09
Rbbr21 netL21 node_3 1717218.9387113666
Cbr21 netL21 node_3 4.986937339731535e-22

* Branch 22
Rabr22 node_1 netRa22 -2301415.8892554883
Lbr22 netRa22 netL22 7.661633998766882e-10
Rbbr22 netL22 node_3 2685448.751867965
Cbr22 netL22 node_3 1.2341880948215986e-22

* Branch 23
Rabr23 node_1 netRa23 -957908.4206788708
Lbr23 netRa23 netL23 1.0573654418731873e-09
Rbbr23 netL23 node_3 1514858.170638505
Cbr23 netL23 node_3 7.186551230773757e-22

* Branch 24
Rabr24 node_1 netRa24 -2363502.333802859
Lbr24 netRa24 netL24 4.945550517477085e-10
Rbbr24 netL24 node_3 2600991.604948785
Cbr24 netL24 node_3 8.02423611736223e-23

* Branch 25
Rabr25 node_1 netRa25 -1068334.4379471
Lbr25 netRa25 netL25 1.0412058983497837e-09
Rbbr25 netL25 node_3 1615231.5729292356
Cbr25 netL25 node_3 5.964316590769096e-22

* Branch 26
Rabr26 node_1 netRa26 -2056597.1660649462
Lbr26 netRa26 netL26 5.971832062527471e-10
Rbbr26 netL26 node_3 2378332.476848623
Cbr26 netL26 node_3 1.2173971300797966e-22

* Branch 27
Rabr27 node_1 netRa27 -2364165.861071747
Lbr27 netRa27 netL27 7.39959378716372e-10
Rbbr27 netL27 node_3 2738231.2653172533
Cbr27 netL27 node_3 1.1396448309387132e-22

* Branch 28
Rabr28 node_1 netRa28 -1990004.854293761
Lbr28 netRa28 netL28 6.248956174360634e-10
Rbbr28 netL28 node_3 2336360.250241641
Cbr28 netL28 node_3 1.34007264583168e-22

* Branch 29
Rabr29 node_1 netRa29 -2334853.2002616706
Lbr29 netRa29 netL29 5.730458311970185e-10
Rbbr29 netL29 node_3 2620040.5726024336
Cbr29 netL29 node_3 9.349383857542475e-23

* Branch 30
Rabr30 node_1 netRa30 236241.67562071388
Lbr30 netRa30 netL30 -1.7714039734093275e-09
Rbbr30 netL30 node_3 -37602769.91704199
Cbr30 netL30 node_3 -1.9699049597531308e-22

* Branch 31
Rabr31 node_1 netRa31 -2921407.531233787
Lbr31 netRa31 netL31 -3.4963071165121693e-09
Rbbr31 netL31 node_3 14590633.103059718
Cbr31 netL31 node_3 -8.208257952324189e-23

* Branch 32
Rabr32 node_1 netRa32 -3752406.411437343
Lbr32 netRa32 netL32 -5.485222809750532e-09
Rbbr32 netL32 node_3 16787017.413364395
Cbr32 netL32 node_3 -8.711976488266776e-23

* Branch 33
Rabr33 node_1 netRa33 -6332599.346354952
Lbr33 netRa33 netL33 -4.2902802225701274e-09
Rbbr33 netL33 node_3 11464133.806197466
Cbr33 netL33 node_3 -5.910924584965652e-23

* Branch 34
Rabr34 node_1 netRa34 -14140495.790780198
Lbr34 netRa34 netL34 -7.155889858375208e-09
Rbbr34 netL34 node_3 20361835.788884547
Cbr34 netL34 node_3 -2.48569039279429e-23

* Branch 35
Rabr35 node_1 netRa35 -46364351.59102785
Lbr35 netRa35 netL35 -1.2028376962020736e-08
Rbbr35 netL35 node_3 51293423.456701435
Cbr35 netL35 node_3 -5.058114230030876e-24

* Branch 36
Rabr36 node_1 netRa36 -7834027689.796539
Lbr36 netRa36 netL36 -1.0671773181279063e-07
Rbbr36 netL36 node_3 7837255674.280837
Cbr36 netL36 node_3 -1.7381548650599366e-27

* Branch 37
Rabr37 node_1 netRa37 -25992607.989125066
Lbr37 netRa37 netL37 -5.01847964797734e-09
Rbbr37 netL37 node_3 28635490.432040382
Cbr37 netL37 node_3 -6.74249170305328e-24

* Branch 38
Rabr38 node_1 netRa38 -604665436.4471807
Lbr38 netRa38 netL38 3.0704428364603544e-08
Rbbr38 netL38 node_3 608044489.613893
Cbr38 netL38 node_3 8.351223301024807e-26

* Branch 39
Rabr39 node_1 netRa39 -46096844.40704829
Lbr39 netRa39 netL39 1.8372129391526834e-08
Rbbr39 netL39 node_3 51535616.83560853
Cbr39 netL39 node_3 7.733538007837745e-24

* Branch 40
Rabr40 node_1 netRa40 -46365694.538370006
Lbr40 netRa40 netL40 2.0904644301205823e-08
Rbbr40 netL40 node_3 51983912.3766401
Cbr40 netL40 node_3 8.673100122023806e-24

* Branch 41
Rabr41 node_1 netRa41 -215629712.96117097
Lbr41 netRa41 netL41 2.1830941884635522e-08
Rbbr41 netL41 node_3 219853517.6991263
Cbr41 netL41 node_3 4.605004610854945e-25

* Branch 42
Rabr42 node_1 netRa42 -34208803.02207873
Lbr42 netRa42 netL42 2.0809759344289477e-08
Rbbr42 netL42 node_3 40101796.386163905
Cbr42 netL42 node_3 1.5169251183720032e-23

* Branch 43
Rabr43 node_1 netRa43 -30464250.563579954
Lbr43 netRa43 netL43 1.88765977907434e-08
Rbbr43 netL43 node_3 36199612.64872377
Cbr43 netL43 node_3 1.711701849734196e-23

* Branch 44
Rabr44 node_1 netRa44 -38453910.45936399
Lbr44 netRa44 netL44 1.8447660371783816e-08
Rbbr44 netL44 node_3 43977443.49791635
Cbr44 netL44 node_3 1.0908622194032997e-23

* Branch 45
Rabr45 node_1 netRa45 -32819545.884784307
Lbr45 netRa45 netL45 2.0918585284444646e-08
Rbbr45 netL45 node_3 38704013.06482025
Cbr45 netL45 node_3 1.646807012112771e-23

* Branch 46
Rabr46 node_1 netRa46 -30861516.5888555
Lbr46 netRa46 netL46 2.0901776199498592e-08
Rbbr46 netL46 node_3 36776116.564192794
Cbr46 netL46 node_3 1.8416167090738802e-23

* Branch 47
Rabr47 node_1 netRa47 -34172036.151603095
Lbr47 netRa47 netL47 1.9434401393617603e-08
Rbbr47 netL47 node_3 39873275.501319066
Cbr47 netL47 node_3 1.4263225333323717e-23

* Branch 48
Rabr48 node_1 netRa48 -29349405.621929
Lbr48 netRa48 netL48 2.1028157459852412e-08
Rbbr48 netL48 node_3 35299308.44086747
Cbr48 netL48 node_3 2.0297144281919957e-23

* Branch 49
Rabr49 node_1 netRa49 -34036824.838352785
Lbr49 netRa49 netL49 1.8123592023444677e-08
Rbbr49 netL49 node_3 39524928.28336677
Cbr49 netL49 node_3 1.3471737340936835e-23

* Branch 50
Rabr50 node_1 netRa50 -39978074.119629495
Lbr50 netRa50 netL50 1.847364398465269e-08
Rbbr50 netL50 node_3 45550927.64853931
Cbr50 netL50 node_3 1.0144561597787118e-23

* Branch 51
Rabr51 node_1 netRa51 -35841837.819213174
Lbr51 netRa51 netL51 1.6975696777659657e-08
Rbbr51 netL51 node_3 41326498.940993726
Cbr51 netL51 node_3 1.1460632858405486e-23

* Branch 52
Rabr52 node_1 netRa52 -41160725.71996506
Lbr52 netRa52 netL52 1.770999430942463e-08
Rbbr52 netL52 node_3 46587226.70003083
Cbr52 netL52 node_3 9.235672438446934e-24

* Branch 53
Rabr53 node_1 netRa53 -14313184.56727283
Lbr53 netRa53 netL53 1.2942529680585616e-08
Rbbr53 netL53 node_3 20655529.846570726
Cbr53 netL53 node_3 4.3776999228817586e-23

* Branch 54
Rabr54 node_1 netRa54 -251926669.91963083
Lbr54 netRa54 netL54 -3.8670436157662155e-08
Rbbr54 netL54 node_3 256903917.03882512
Cbr54 netL54 node_3 -5.974951051693424e-25

* Branch 55
Rabr55 node_1 netRa55 -79176664.08226584
Lbr55 netRa55 netL55 -2.0496562849389536e-08
Rbbr55 netL55 node_3 84164555.06777816
Cbr55 netL55 node_3 -3.0757779227037412e-24

* Branch 56
Rabr56 node_1 netRa56 -47523461.98469654
Lbr56 netRa56 netL56 -1.6294583120037242e-08
Rbbr56 netL56 node_3 52582817.22272752
Cbr56 netL56 node_3 -6.520664506094129e-24

* Branch 57
Rabr57 node_1 netRa57 -36799665.414526366
Lbr57 netRa57 netL57 -1.5741445374477023e-08
Rbbr57 netL57 node_3 42226548.681217544
Cbr57 netL57 node_3 -1.013014910427639e-23

* Branch 58
Rabr58 node_1 netRa58 -21123207.625088487
Lbr58 netRa58 netL58 -1.1613422068549293e-08
Rbbr58 netL58 node_3 26689079.39413298
Cbr58 netL58 node_3 -2.060002134068124e-23

* Branch 59
Rabr59 node_1 netRa59 -38566997.39830398
Lbr59 netRa59 netL59 -1.4103657823146674e-08
Rbbr59 netL59 node_3 43596645.03941362
Cbr59 netL59 node_3 -8.388099334524442e-24

* Branch 60
Rabr60 node_1 netRa60 -47756270.67916401
Lbr60 netRa60 netL60 -1.5292918106545883e-08
Rbbr60 netL60 node_3 52707238.667862915
Cbr60 netL60 node_3 -6.075616198397572e-24

* Branch 61
Rabr61 node_1 netRa61 -28170888.095805317
Lbr61 netRa61 netL61 -1.4220165013070038e-08
Rbbr61 netL61 node_3 33726910.58758687
Cbr61 netL61 node_3 -1.496679710422514e-23

* Branch 62
Rabr62 node_1 netRa62 -32428480.88830544
Lbr62 netRa62 netL62 -1.247685294242122e-08
Rbbr62 netL62 node_3 37456494.772631906
Cbr62 netL62 node_3 -1.0271936779897895e-23

* Branch 63
Rabr63 node_1 netRa63 -48825028.72545902
Lbr63 netRa63 netL63 -1.4719217964416938e-08
Rbbr63 netL63 node_3 53637240.31061014
Cbr63 netL63 node_3 -5.620521678979537e-24

* Branch 64
Rabr64 node_1 netRa64 -60735098.34322831
Lbr64 netRa64 netL64 -1.610437490160227e-08
Rbbr64 netL64 node_3 65527047.2051161
Cbr64 netL64 node_3 -4.04654509734453e-24

* Branch 65
Rabr65 node_1 netRa65 -44030537.76524635
Lbr65 netRa65 netL65 -1.334387321398929e-08
Rbbr65 netL65 node_3 48723767.20917831
Cbr65 netL65 node_3 -6.2199687418398344e-24

* Branch 66
Rabr66 node_1 netRa66 -49759299.05231397
Lbr66 netRa66 netL66 -1.398276763716396e-08
Rbbr66 netL66 node_3 54472638.88580914
Cbr66 netL66 node_3 -5.1587178056208255e-24

* Branch 67
Rabr67 node_1 netRa67 -96607243.57214159
Lbr67 netRa67 netL67 -1.874497728333693e-08
Rbbr67 netL67 node_3 101114312.75074494
Cbr67 netL67 node_3 -1.9189501646221828e-24

* Branch 68
Rabr68 node_1 netRa68 -60432620.97367551
Lbr68 netRa68 netL68 -1.4390811616447339e-08
Rbbr68 netL68 node_3 64957436.9089837
Cbr68 netL68 node_3 -3.665956496787425e-24

* Branch 69
Rabr69 node_1 netRa69 -23898308.661669366
Lbr69 netRa69 netL69 -9.536308809176706e-09
Rbbr69 netL69 node_3 28767141.46794307
Cbr69 netL69 node_3 -1.387140387360034e-23

* Branch 70
Rabr70 node_1 netRa70 -14935070438.121784
Lbr70 netRa70 netL70 1.3096889082839265e-07
Rbbr70 netL70 node_3 14937808237.23394
Cbr70 netL70 node_3 5.870483936029953e-28

* Branch 71
Rabr71 node_1 netRa71 -65258609.83593523
Lbr71 netRa71 netL71 -1.4766333987068472e-08
Rbbr71 netL71 node_3 69809267.22556327
Cbr71 netL71 node_3 -3.2413367046094084e-24

* Branch 72
Rabr72 node_1 netRa72 -82910473.06603399
Lbr72 netRa72 netL72 -2.075032683839803e-08
Rbbr72 netL72 node_3 90880012.41955045
Cbr72 netL72 node_3 -2.7539264549714224e-24

* Branch 73
Rabr73 node_1 netRa73 -129648260.782479
Lbr73 netRa73 netL73 -2.1309828195050732e-08
Rbbr73 netL73 node_3 135998726.1502744
Cbr73 netL73 node_3 -1.2085988611497834e-24

* Branch 74
Rabr74 node_1 netRa74 -5689387.498269622
Lbr74 netRa74 netL74 -4.951549680561666e-09
Rbbr74 netL74 node_3 11740893.4243924
Cbr74 netL74 node_3 -7.413040942922704e-23

* Branch 75
Rabr75 node_1 netRa75 -11661612.872781783
Lbr75 netRa75 netL75 -5.211705306666747e-09
Rbbr75 netL75 node_3 15998017.50028048
Cbr75 netL75 node_3 -2.7936385297332575e-23

* Branch 76
Rabr76 node_1 netRa76 -4101503.397476933
Lbr76 netRa76 netL76 -4.51531000745857e-09
Rbbr76 netL76 node_3 11295166.679588819
Cbr76 netL76 node_3 -9.747447841611815e-23

* Branch 77
Rabr77 node_1 netRa77 -17170030.049334202
Lbr77 netRa77 netL77 -4.92509133089364e-09
Rbbr77 netL77 node_3 20459859.357097857
Cbr77 netL77 node_3 -1.4020142678537178e-23

* Branch 78
Rabr78 node_1 netRa78 -15353792.03644039
Lbr78 netRa78 netL78 -4.589072764264325e-09
Rbbr78 netL78 node_3 18473298.527810175
Cbr78 netL78 node_3 -1.618000677700262e-23

* Branch 79
Rabr79 node_1 netRa79 -3513224.8182573216
Lbr79 netRa79 netL79 -2.607167516478133e-09
Rbbr79 netL79 node_3 7605322.308713122
Cbr79 netL79 node_3 -9.758575835362106e-23

* Branch 80
Rabr80 node_1 netRa80 -1495753.2894245412
Lbr80 netRa80 netL80 -2.3287155215037317e-09
Rbbr80 netL80 node_3 8791217.68411539
Cbr80 netL80 node_3 -1.7713530531371393e-22

* Branch 81
Rabr81 node_1 netRa81 822356.2488255586
Lbr81 netRa81 netL81 -3.356976113261903e-09
Rbbr81 netL81 node_3 -21236465.326483816
Cbr81 netL81 node_3 -1.9210398976815375e-22

* Branch 82
Rabr82 node_1 netRa82 -3427765.0334689966
Lbr82 netRa82 netL82 -2.091024819628199e-09
Rbbr82 netL82 node_3 6540052.952139069
Cbr82 netL82 node_3 -9.328428309176263e-23

* Branch 83
Rabr83 node_1 netRa83 1460374.4546107957
Lbr83 netRa83 netL83 -2.11298885011282e-09
Rbbr83 netL83 node_3 -7766465.741568255
Cbr83 netL83 node_3 -1.8625490890646478e-22

* Branch 84
Rabr84 node_1 netRa84 -4213288.744609897
Lbr84 netRa84 netL84 -6.2797017332579635e-09
Rbbr84 netL84 node_3 19857469.65099775
Cbr84 netL84 node_3 -7.507777517152941e-23

* Branch 85
Rabr85 node_1 netRa85 -580671023.1047786
Lbr85 netRa85 netL85 -1.6995374199050504e-08
Rbbr85 netL85 node_3 582373794.5369569
Cbr85 netL85 node_3 -5.0257534544401404e-26

* Branch 86
Rabr86 node_1 netRa86 -1591432.0623940781
Lbr86 netRa86 netL86 -2.7408609390654427e-09
Rbbr86 netL86 node_3 10852018.924725648
Cbr86 netL86 node_3 -1.5875895834804229e-22

* Branch 87
Rabr87 node_1 netRa87 -2592497.997056714
Lbr87 netRa87 netL87 -1.9480153557219415e-09
Rbbr87 netL87 node_3 6246565.632822372
Cbr87 netL87 node_3 -1.203094063667365e-22

* Branch 88
Rabr88 node_1 netRa88 -1999777.0786529782
Lbr88 netRa88 netL88 -1.4320182227870255e-09
Rbbr88 netL88 node_3 4737159.670676781
Cbr88 netL88 node_3 -1.5118765417817346e-22

* Branch 89
Rabr89 node_1 netRa89 -1861735.9186118233
Lbr89 netRa89 netL89 -1.6366536680577263e-09
Rbbr89 netL89 node_3 5535816.5484995255
Cbr89 netL89 node_3 -1.5883304868458466e-22

* Branch 90
Rabr90 node_1 netRa90 -1104845.3124504315
Lbr90 netRa90 netL90 -1.3174177465487238e-09
Rbbr90 netL90 node_3 5207347.761150681
Cbr90 netL90 node_3 -2.290456337029294e-22

* Branch 91
Rabr91 node_1 netRa91 -65327.18909421534
Lbr91 netRa91 netL91 -4.891765960384366e-10
Rbbr91 netL91 node_3 11451997.22664188
Cbr91 netL91 node_3 -6.566422279874339e-22

* Branch 92
Rabr92 node_1 netRa92 -113497.88183159671
Lbr92 netRa92 netL92 -4.3562200912383463e-10
Rbbr92 netL92 node_3 5407520.128745571
Cbr92 netL92 node_3 -7.114830201364196e-22

* Branch 93
Rabr93 node_1 netRa93 -80566.63176479202
Lbr93 netRa93 netL93 -5.690238078832868e-10
Rbbr93 netL93 node_3 12321935.100088246
Cbr93 netL93 node_3 -5.7574825294046945e-22

* Branch 94
Rabr94 node_1 netRa94 -352971.4408756905
Lbr94 netRa94 netL94 -4.601362674782577e-10
Rbbr94 netL94 node_3 2287598.519445864
Cbr94 netL94 node_3 -5.703860463067452e-22

* Branch 95
Rabr95 node_1 netRa95 -23520509913.565907
Lbr95 netRa95 netL95 1.1980784977437485e-07
Rbbr95 netL95 node_3 23522554895.719658
Cbr95 netL95 node_3 2.1654714665731033e-28

* Branch 96
Rabr96 node_1 netRa96 -1151442.8280979756
Lbr96 netRa96 netL96 -7.952164663196181e-10
Rbbr96 netL96 node_3 2957116.8787769917
Cbr96 netL96 node_3 -2.3368082435600953e-22

* Branch 97
Rabr97 node_1 netRa97 591127.1192291913
Lbr97 netRa97 netL97 -6.022367516201421e-10
Rbbr97 netL97 node_3 -2412288.605119564
Cbr97 netL97 node_3 -4.2197580775815993e-22

* Branch 98
Rabr98 node_1 netRa98 9797926.37666514
Lbr98 netRa98 netL98 -1.9141211917410416e-09
Rbbr98 netL98 node_3 -10885910.908759203
Cbr98 netL98 node_3 -1.7942448473971258e-23

* Branch 99
Rabr99 node_1 netRa99 360604.0469816219
Lbr99 netRa99 netL99 1.244264993516603e-10
Rbbr99 netL99 node_3 -509608.90319206665
Cbr99 netL99 node_3 6.821730707931636e-22

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 542689.1513992626
Lbr0 netRa0 netL0 -1.2267421465734285e-10
Rbbr0 netL0 node_4 -628399.0415099346
Cbr0 netL0 node_4 -3.534065437676932e-22

* Branch 1
Rabr1 node_1 netRa1 447206.85416959616
Lbr1 netRa1 netL1 -1.0732557605363012e-10
Rbbr1 netL1 node_4 -527536.6621936715
Cbr1 netL1 node_4 -4.476193366551902e-22

* Branch 2
Rabr2 node_1 netRa2 380122.5877658833
Lbr2 netRa2 netL2 -9.2272151505239e-11
Rbbr2 netL2 node_4 -451216.1641861466
Cbr2 netL2 node_4 -5.311361053109372e-22

* Branch 3
Rabr3 node_1 netRa3 560907537.1725335
Lbr3 netRa3 netL3 -5.174266822948842e-09
Rbbr3 netL3 node_4 -561035492.4153266
Cbr3 netL3 node_4 -1.6435529335340026e-26

* Branch 4
Rabr4 node_1 netRa4 97778119.38477397
Lbr4 netRa4 netL4 2.1771652361123505e-09
Rbbr4 netL4 node_4 -97908645.83929859
Cbr4 netL4 node_4 2.275723446995548e-25

* Branch 5
Rabr5 node_1 netRa5 364730.8381495859
Lbr5 netRa5 netL5 -7.980251265808303e-11
Rbbr5 netL5 node_4 -422193.383585675
Cbr5 netL5 node_4 -5.150122526448769e-22

* Branch 6
Rabr6 node_1 netRa6 100667.65955059578
Lbr6 netRa6 netL6 -7.654728093084315e-11
Rbbr6 netL6 node_4 -272749.04783180926
Cbr6 netL6 node_4 -2.7390546196792237e-21

* Branch 7
Rabr7 node_1 netRa7 610633.6714629335
Lbr7 netRa7 netL7 -2.18979792138355e-10
Rbbr7 netL7 node_4 -779782.4769747141
Cbr7 netL7 node_4 -4.561540611272696e-22

* Branch 8
Rabr8 node_1 netRa8 604807.967681163
Lbr8 netRa8 netL8 -2.2671699856584267e-10
Rbbr8 netL8 node_4 -782812.9093945642
Cbr8 netL8 node_4 -4.751812406776017e-22

* Branch 9
Rabr9 node_1 netRa9 798400.3228721467
Lbr9 netRa9 netL9 -2.1821667495494331e-10
Rbbr9 netL9 node_4 -938056.9287507643
Cbr9 netL9 node_4 -2.899962783375214e-22

* Branch 10
Rabr10 node_1 netRa10 310299.3372515673
Lbr10 netRa10 netL10 -3.1887062697250817e-10
Rbbr10 netL10 node_4 -625206.1780833984
Cbr10 netL10 node_4 -1.6172581681546202e-21

* Branch 11
Rabr11 node_1 netRa11 3026634.467024937
Lbr11 netRa11 netL11 -3.710714986975806e-10
Rbbr11 netL11 node_4 -3141850.975184557
Cbr11 netL11 node_4 -3.8946417559700293e-23

* Branch 12
Rabr12 node_1 netRa12 288443.907257376
Lbr12 netRa12 netL12 -3.25686091884457e-10
Rbbr12 netL12 node_4 -613093.282639334
Cbr12 netL12 node_4 -1.8095024371067116e-21

* Branch 13
Rabr13 node_1 netRa13 181052.81947096097
Lbr13 netRa13 netL13 -7.373760512150967e-10
Rbbr13 netL13 node_4 -8050433.181386143
Cbr13 netL13 node_4 -4.760291857272652e-22

* Branch 14
Rabr14 node_1 netRa14 332771.79010588204
Lbr14 netRa14 netL14 -3.117158724884379e-10
Rbbr14 netL14 node_4 -637452.954290281
Cbr14 netL14 node_4 -1.4487277444869423e-21

* Branch 15
Rabr15 node_1 netRa15 266782.5552360517
Lbr15 netRa15 netL15 -3.321195788625964e-10
Rbbr15 netL15 node_4 -600883.0608837282
Cbr15 netL15 node_4 -2.0331068413572197e-21

* Branch 16
Rabr16 node_1 netRa16 17761803.320297956
Lbr16 netRa16 netL16 8.954938862268284e-10
Rbbr16 netL16 node_4 -17882132.355406746
Cbr16 netL16 node_4 2.821506900957534e-24

* Branch 17
Rabr17 node_1 netRa17 245426.41386833906
Lbr17 netRa17 netL17 -3.3844001959118264e-10
Rbbr17 netL17 node_4 -588873.2604443784
Cbr17 netL17 node_4 -2.295453650823669e-21

* Branch 18
Rabr18 node_1 netRa18 405366.46629150095
Lbr18 netRa18 netL18 -2.9033609120102335e-10
Rbbr18 netL18 node_4 -678471.5322364895
Cbr18 netL18 node_4 -1.0447889427442817e-21

* Branch 19
Rabr19 node_1 netRa19 441060.09830102546
Lbr19 netRa19 netL19 -2.853634849578652e-10
Rbbr19 netL19 node_4 -701691.8940509865
Cbr19 netL19 node_4 -9.13754418293771e-22

* Branch 20
Rabr20 node_1 netRa20 224543.8557587763
Lbr20 netRa20 netL20 -3.44674936570988e-10
Rbbr20 netL20 node_4 -577026.4252926718
Cbr20 netL20 node_4 -2.604784993926788e-21

* Branch 21
Rabr21 node_1 netRa21 356872.9972737932
Lbr21 netRa21 netL21 -3.0460669028192175e-10
Rbbr21 netL21 node_4 -650907.4965507705
Cbr21 netL21 node_4 -1.2960948269802043e-21

* Branch 22
Rabr22 node_1 netRa22 204056.3930925654
Lbr22 netRa22 netL22 -3.507537670393374e-10
Rbbr22 netL22 node_4 -565279.7521305572
Cbr22 netL22 node_4 -2.9724011634231445e-21

* Branch 23
Rabr23 node_1 netRa23 382843.94903294934
Lbr23 netRa23 netL23 -2.98682790732954e-10
Rbbr23 netL23 node_4 -666924.7635008798
Cbr23 netL23 node_4 -1.1579757937750426e-21

* Branch 24
Rabr24 node_1 netRa24 184209.4176679176
Lbr24 netRa24 netL24 -3.5673079434461714e-10
Rbbr24 netL24 node_4 -553974.9055500918
Cbr24 netL24 node_4 -3.410389714126335e-21

* Branch 25
Rabr25 node_1 netRa25 165191.92892422588
Lbr25 netRa25 netL25 -3.6310255270970943e-10
Rbbr25 netL25 node_4 -542962.3488308816
Cbr25 netL25 node_4 -3.9420649865350185e-21

* Branch 26
Rabr26 node_1 netRa26 447976.590380895
Lbr26 netRa26 netL26 -2.7733741034413695e-10
Rbbr26 netL26 node_4 -707159.4142151418
Cbr26 netL26 node_4 -8.689719422340481e-22

* Branch 27
Rabr27 node_1 netRa27 272887.8340014151
Lbr27 netRa27 netL27 -1.8643278120434933e-10
Rbbr27 netL27 node_4 -617457.8098015024
Cbr27 netL27 node_4 -1.0974553917946942e-21

* Branch 28
Rabr28 node_1 netRa28 547927.9456490262
Lbr28 netRa28 netL28 -2.7267142961848684e-10
Rbbr28 netL28 node_4 -771629.5415777316
Cbr28 netL28 node_4 -6.425276870739961e-22

* Branch 29
Rabr29 node_1 netRa29 424579.386174464
Lbr29 netRa29 netL29 -2.2956869471104288e-10
Rbbr29 netL29 node_4 -643784.5679918395
Cbr29 netL29 node_4 -8.366437227712949e-22

* Branch 30
Rabr30 node_1 netRa30 488721.77281750226
Lbr30 netRa30 netL30 -2.2930370100429297e-10
Rbbr30 netL30 node_4 -690898.2529552222
Cbr30 netL30 node_4 -6.773396749454134e-22

* Branch 31
Rabr31 node_1 netRa31 736310.6618638322
Lbr31 netRa31 netL31 -2.512217173384756e-10
Rbbr31 netL31 node_4 -912059.6667053038
Cbr31 netL31 node_4 -3.7351330673719953e-22

* Branch 32
Rabr32 node_1 netRa32 -632841.0259563685
Lbr32 netRa32 netL32 4.505070243920217e-10
Rbbr32 netL32 node_4 1563331.77512591
Cbr32 netL32 node_4 4.542254535722797e-22

* Branch 33
Rabr33 node_1 netRa33 8028100.236855678
Lbr33 netRa33 netL33 -1.2309212135583314e-09
Rbbr33 netL33 node_4 -8675021.977770152
Cbr33 netL33 node_4 -1.767410227758547e-23

* Branch 34
Rabr34 node_1 netRa34 -17593710.629390817
Lbr34 netRa34 netL34 -2.592014008985538e-09
Rbbr34 netL34 node_4 18728916.10807599
Cbr34 netL34 node_4 -7.866302122786872e-24

* Branch 35
Rabr35 node_1 netRa35 -2077531.7880725777
Lbr35 netRa35 netL35 3.0966403483616347e-09
Rbbr35 netL35 node_4 5226126.709173862
Cbr35 netL35 node_4 2.852076074707e-22

* Branch 36
Rabr36 node_1 netRa36 2709269.7405383307
Lbr36 netRa36 netL36 3.327619057151884e-09
Rbbr36 netL36 node_4 -5619854.664174579
Cbr36 netL36 node_4 2.185537177680587e-22

* Branch 37
Rabr37 node_1 netRa37 7688.8259556667945
Lbr37 netRa37 netL37 2.5112017679503312e-09
Rbbr37 netL37 node_4 -536110943.4211978
Cbr37 netL37 node_4 6.099841697972077e-22

* Branch 38
Rabr38 node_1 netRa38 797662.5039661435
Lbr38 netRa38 netL38 2.6488397912188715e-09
Rbbr38 netL38 node_4 -6287672.917338242
Cbr38 netL38 node_4 5.28146620045198e-22

* Branch 39
Rabr39 node_1 netRa39 1190571.6100210813
Lbr39 netRa39 netL39 2.6856753467980347e-09
Rbbr39 netL39 node_4 -5690514.7328935275
Cbr39 netL39 node_4 3.964166885035633e-22

* Branch 40
Rabr40 node_1 netRa40 1208152.308509651
Lbr40 netRa40 netL40 2.9681256547685192e-09
Rbbr40 netL40 node_4 -5554792.328879182
Cbr40 netL40 node_4 4.422822417269749e-22

* Branch 41
Rabr41 node_1 netRa41 1510026.803326887
Lbr41 netRa41 netL41 2.6943348269288636e-09
Rbbr41 netL41 node_4 -5231226.231284848
Cbr41 netL41 node_4 3.4108991726707467e-22

* Branch 42
Rabr42 node_1 netRa42 1191216.695275895
Lbr42 netRa42 netL42 2.949110897328096e-09
Rbbr42 netL42 node_4 -5343292.8001565235
Cbr42 netL42 node_4 4.63340443916901e-22

* Branch 43
Rabr43 node_1 netRa43 1599621.5421481712
Lbr43 netRa43 netL43 2.7384029511308552e-09
Rbbr43 netL43 node_4 -5377867.121004925
Cbr43 netL43 node_4 3.18329092328065e-22

* Branch 44
Rabr44 node_1 netRa44 1068957.8664850455
Lbr44 netRa44 netL44 3.0068063511832434e-09
Rbbr44 netL44 node_4 -5652452.404023816
Cbr44 netL44 node_4 4.976461613390128e-22

* Branch 45
Rabr45 node_1 netRa45 1894419.2385197096
Lbr45 netRa45 netL45 2.7103592184347447e-09
Rbbr45 netL45 node_4 -5145965.7506793365
Cbr45 netL45 node_4 2.780291894389088e-22

* Branch 46
Rabr46 node_1 netRa46 1624470.8279339976
Lbr46 netRa46 netL46 2.621210212335642e-09
Rbbr46 netL46 node_4 -5311462.839334532
Cbr46 netL46 node_4 3.0379755222622995e-22

* Branch 47
Rabr47 node_1 netRa47 1103670.6014226824
Lbr47 netRa47 netL47 3.0457760154836533e-09
Rbbr47 netL47 node_4 -5439345.660109303
Cbr47 netL47 node_4 5.073728160380357e-22

* Branch 48
Rabr48 node_1 netRa48 1828525.673652638
Lbr48 netRa48 netL48 2.564591809309263e-09
Rbbr48 netL48 node_4 -5085845.766016468
Cbr48 netL48 node_4 2.7578017444404737e-22

* Branch 49
Rabr49 node_1 netRa49 892418.4949200155
Lbr49 netRa49 netL49 2.9267331458101264e-09
Rbbr49 netL49 node_4 -5599089.643875553
Cbr49 netL49 node_4 5.857600248514415e-22

* Branch 50
Rabr50 node_1 netRa50 2169432.0386737077
Lbr50 netRa50 netL50 2.6948741079858906e-09
Rbbr50 netL50 node_4 -5316387.243954852
Cbr50 netL50 node_4 2.336601066457336e-22

* Branch 51
Rabr51 node_1 netRa51 893571.1400545044
Lbr51 netRa51 netL51 3.0863267822549545e-09
Rbbr51 netL51 node_4 -5856198.745397623
Cbr51 netL51 node_4 5.8982468464588095e-22

* Branch 52
Rabr52 node_1 netRa52 742514.2842201982
Lbr52 netRa52 netL52 3.043534621837658e-09
Rbbr52 netL52 node_4 -6248730.940635418
Cbr52 netL52 node_4 6.560189274017426e-22

* Branch 53
Rabr53 node_1 netRa53 1601825.5626490144
Lbr53 netRa53 netL53 2.405693541432625e-09
Rbbr53 netL53 node_4 -5125265.398295923
Cbr53 netL53 node_4 2.930364493498315e-22

* Branch 54
Rabr54 node_1 netRa54 10967844.270469584
Lbr54 netRa54 netL54 -4.603463203782058e-09
Rbbr54 netL54 node_4 -14018963.44758674
Cbr54 netL54 node_4 -2.993944720870726e-23

* Branch 55
Rabr55 node_1 netRa55 645152.7316749261
Lbr55 netRa55 netL55 3.0357666743734664e-09
Rbbr55 netL55 node_4 -6613932.19044902
Cbr55 netL55 node_4 7.115235193478216e-22

* Branch 56
Rabr56 node_1 netRa56 1936959.4862555468
Lbr56 netRa56 netL56 2.4820328619562423e-09
Rbbr56 netL56 node_4 -5152430.9055768
Cbr56 netL56 node_4 2.487065892311864e-22

* Branch 57
Rabr57 node_1 netRa57 417459.75179047784
Lbr57 netRa57 netL57 2.9838783677602875e-09
Rbbr57 netL57 node_4 -8841465.50036364
Cbr57 netL57 node_4 8.085627929900453e-22

* Branch 58
Rabr58 node_1 netRa58 1635996.2555602528
Lbr58 netRa58 netL58 2.3536207913965183e-09
Rbbr58 netL58 node_4 -5182648.191887268
Cbr58 netL58 node_4 2.7760014120985307e-22

* Branch 59
Rabr59 node_1 netRa59 1936047.376711511
Lbr59 netRa59 netL59 2.353221835549177e-09
Rbbr59 netL59 node_4 -5038044.280630328
Cbr59 netL59 node_4 2.412693953505247e-22

* Branch 60
Rabr60 node_1 netRa60 2067174.8494030146
Lbr60 netRa60 netL60 2.402969624464676e-09
Rbbr60 netL60 node_4 -5201901.252583015
Cbr60 netL60 node_4 2.2347487130502137e-22

* Branch 61
Rabr61 node_1 netRa61 1660674.2917293597
Lbr61 netRa61 netL61 2.127851823616677e-09
Rbbr61 netL61 node_4 -4825003.007769393
Cbr61 netL61 node_4 2.6557381424004603e-22

* Branch 62
Rabr62 node_1 netRa62 2000834.6450047405
Lbr62 netRa62 netL62 2.26342320415114e-09
Rbbr62 netL62 node_4 -5072392.465027967
Cbr62 netL62 node_4 2.230326323697306e-22

* Branch 63
Rabr63 node_1 netRa63 1723211.58197449
Lbr63 netRa63 netL63 2.0239303042598715e-09
Rbbr63 netL63 node_4 -4669136.946066044
Cbr63 netL63 node_4 2.5157138788689267e-22

* Branch 64
Rabr64 node_1 netRa64 1245506.8133132663
Lbr64 netRa64 netL64 1.905453065215457e-09
Rbbr64 netL64 node_4 -4975785.197220528
Cbr64 netL64 node_4 3.075083033495433e-22

* Branch 65
Rabr65 node_1 netRa65 38247919.70771529
Lbr65 netRa65 netL65 7.136559842452163e-09
Rbbr65 netL65 node_4 -40598072.87277701
Cbr65 netL65 node_4 4.596051598428727e-24

* Branch 66
Rabr66 node_1 netRa66 1244778.40462945
Lbr66 netRa66 netL66 1.802897859749662e-09
Rbbr66 netL66 node_4 -4693259.069851086
Cbr66 netL66 node_4 3.086626178709646e-22

* Branch 67
Rabr67 node_1 netRa67 1352297.54685296
Lbr67 netRa67 netL67 1.8476349740213654e-09
Rbbr67 netL67 node_4 -4791068.91406231
Cbr67 netL67 node_4 2.8523071543968343e-22

* Branch 68
Rabr68 node_1 netRa68 336139.03645059426
Lbr68 netRa68 netL68 1.5030981618817e-09
Rbbr68 netL68 node_4 -9782631.373273533
Cbr68 netL68 node_4 4.575078916823466e-22

* Branch 69
Rabr69 node_1 netRa69 15054209.561699612
Lbr69 netRa69 netL69 5.665565733933249e-09
Rbbr69 netL69 node_4 -18518840.4507494
Cbr69 netL69 node_4 2.032401804216879e-23

* Branch 70
Rabr70 node_1 netRa70 -91671.72211460707
Lbr70 netRa70 netL70 1.4116338869467818e-09
Rbbr70 netL70 node_4 31407075.29107695
Cbr70 netL70 node_4 4.881124750682557e-22

* Branch 71
Rabr71 node_1 netRa71 12561619.100840924
Lbr71 netRa71 netL71 2.9287785718750848e-09
Rbbr71 netL71 node_4 -14077610.443971721
Cbr71 netL71 node_4 1.6563140804445002e-23

* Branch 72
Rabr72 node_1 netRa72 4057692.3209864805
Lbr72 netRa72 netL72 2.2652934856248463e-09
Rbbr72 netL72 node_4 -6474611.448316166
Cbr72 netL72 node_4 8.624098001290526e-23

* Branch 73
Rabr73 node_1 netRa73 1732053.9136387913
Lbr73 netRa73 netL73 2.3424385857577634e-09
Rbbr73 netL73 node_4 -6595526.177875991
Cbr73 netL73 node_4 2.0515144590411667e-22

* Branch 74
Rabr74 node_1 netRa74 -1443940.9113786118
Lbr74 netRa74 netL74 1.606162235440666e-09
Rbbr74 netL74 node_4 4106214.7755967914
Cbr74 netL74 node_4 2.7078040037207032e-22

* Branch 75
Rabr75 node_1 netRa75 1723341.6591822496
Lbr75 netRa75 netL75 1.5312098792387442e-09
Rbbr75 netL75 node_4 -4257067.773866086
Cbr75 netL75 node_4 2.0878838063238267e-22

* Branch 76
Rabr76 node_1 netRa76 2764513.2498609866
Lbr76 netRa76 netL76 2.8496029705173237e-09
Rbbr76 netL76 node_4 -8092001.707441625
Cbr76 netL76 node_4 1.274347802786421e-22

* Branch 77
Rabr77 node_1 netRa77 157566.41387785735
Lbr77 netRa77 netL77 9.132826306093527e-10
Rbbr77 netL77 node_4 -10833441.530096715
Cbr77 netL77 node_4 5.363536060061078e-22

* Branch 78
Rabr78 node_1 netRa78 631075.7445094535
Lbr78 netRa78 netL78 8.436463361128038e-10
Rbbr78 netL78 node_4 -3017403.2316000494
Cbr78 netL78 node_4 4.432985401072447e-22

* Branch 79
Rabr79 node_1 netRa79 509601.9463692469
Lbr79 netRa79 netL79 2.0644233530476403e-09
Rbbr79 netL79 node_4 -14904966.520630557
Cbr79 netL79 node_4 2.723398051540753e-22

* Branch 80
Rabr80 node_1 netRa80 -3172051.694265325
Lbr80 netRa80 netL80 1.1889551431764514e-09
Rbbr80 netL80 node_4 4091404.3998180456
Cbr80 netL80 node_4 9.159473445292443e-23

* Branch 81
Rabr81 node_1 netRa81 630613.0889490355
Lbr81 netRa81 netL81 8.339494329357347e-10
Rbbr81 netL81 node_4 -3022181.3419746766
Cbr81 netL81 node_4 4.378756568802338e-22

* Branch 82
Rabr82 node_1 netRa82 618241.8846442995
Lbr82 netRa82 netL82 7.208922177320569e-10
Rbbr82 netL82 node_4 -2576894.526815628
Cbr82 netL82 node_4 4.527958876181084e-22

* Branch 83
Rabr83 node_1 netRa83 -6205236.282997598
Lbr83 netRa83 netL83 1.5325567529060463e-09
Rbbr83 netL83 node_4 7353478.355959353
Cbr83 netL83 node_4 3.358176085132488e-23

* Branch 84
Rabr84 node_1 netRa84 676769.1650768865
Lbr84 netRa84 netL84 8.456093257855373e-10
Rbbr84 netL84 node_4 -3081247.8975758497
Cbr84 netL84 node_4 4.0580507095917956e-22

* Branch 85
Rabr85 node_1 netRa85 59051.45485179931
Lbr85 netRa85 netL85 1.0475067963916961e-09
Rbbr85 netL85 node_4 -36884907.457564786
Cbr85 netL85 node_4 4.860054831338219e-22

* Branch 86
Rabr86 node_1 netRa86 691687.0857756826
Lbr86 netRa86 netL86 6.999613218172635e-10
Rbbr86 netL86 node_4 -2420609.9092751658
Cbr86 netL86 node_4 4.18322251293343e-22

* Branch 87
Rabr87 node_1 netRa87 723353.722885445
Lbr87 netRa87 netL87 7.697817908794776e-10
Rbbr87 netL87 node_4 -2677115.6975121954
Cbr87 netL87 node_4 3.977770872273977e-22

* Branch 88
Rabr88 node_1 netRa88 -2649697.7675919146
Lbr88 netRa88 netL88 1.7942802823123467e-09
Rbbr88 netL88 node_4 4679504.836565366
Cbr88 netL88 node_4 1.4464136220561061e-22

* Branch 89
Rabr89 node_1 netRa89 -743852.0682643781
Lbr89 netRa89 netL89 5.672324978733773e-10
Rbbr89 netL89 node_4 2082408.8593627552
Cbr89 netL89 node_4 3.6597952495350228e-22

* Branch 90
Rabr90 node_1 netRa90 17931.82485625446
Lbr90 netRa90 netL90 4.46572750630918e-10
Rbbr90 netL90 node_4 -28406498.26494108
Cbr90 netL90 node_4 8.965658207526638e-22

* Branch 91
Rabr91 node_1 netRa91 -356524.1451733075
Lbr91 netRa91 netL91 3.7288955252490017e-10
Rbbr91 netL91 node_4 1587620.2027121913
Cbr91 netL91 node_4 6.58144684856771e-22

* Branch 92
Rabr92 node_1 netRa92 -91144.69725391743
Lbr92 netRa92 netL92 2.9619819896329683e-10
Rbbr92 netL92 node_4 2595148.079377876
Cbr92 netL92 node_4 1.2477283719828608e-21

* Branch 93
Rabr93 node_1 netRa93 -114758.49506859451
Lbr93 netRa93 netL93 2.9392785127510323e-10
Rbbr93 netL93 node_4 2533992.256791938
Cbr93 netL93 node_4 1.0076873053434576e-21

* Branch 94
Rabr94 node_1 netRa94 -247315.42477064914
Lbr94 netRa94 netL94 3.4501358326757653e-10
Rbbr94 netL94 node_4 1474021.618800555
Cbr94 netL94 node_4 9.447791708390938e-22

* Branch 95
Rabr95 node_1 netRa95 -316955.26021051407
Lbr95 netRa95 netL95 2.3814315340491517e-10
Rbbr95 netL95 node_4 904371.7090653612
Cbr95 netL95 node_4 8.294465927872829e-22

* Branch 96
Rabr96 node_1 netRa96 -89454.15553986085
Lbr96 netRa96 netL96 1.5576119644376803e-10
Rbbr96 netL96 node_4 810232.129163888
Cbr96 netL96 node_4 2.1406964615781944e-21

* Branch 97
Rabr97 node_1 netRa97 -573150.0933063151
Lbr97 netRa97 netL97 2.9648450026470134e-10
Rbbr97 netL97 node_4 1086135.3309084196
Cbr97 netL97 node_4 4.753962281591072e-22

* Branch 98
Rabr98 node_1 netRa98 140084.25795128747
Lbr98 netRa98 netL98 9.094336551240397e-11
Rbbr98 netL98 node_4 -300678.49872070405
Cbr98 netL98 node_4 2.1676290548444107e-21

* Branch 99
Rabr99 node_1 netRa99 -216534.59114695946
Lbr99 netRa99 netL99 7.550747596015935e-11
Rbbr99 netL99 node_4 306553.20170534
Cbr99 netL99 node_4 1.1297508684543246e-21

.ends


* Y'22
.subckt yp22 node_2 0
* Branch 0
Rabr0 node_2 netRa0 -31126.722783627214
Lbr0 netRa0 netL0 -2.2110341770271838e-11
Rbbr0 netL0 0 44981.268215747245
Cbr0 netL0 0 -1.6693519208422308e-20

* Branch 1
Rabr1 node_2 netRa1 -13647.32797262034
Lbr1 netRa1 netL1 -1.3917776502083044e-11
Rbbr1 netL1 0 26020.03202503799
Cbr1 netL1 0 -4.102990019861086e-20

* Branch 2
Rabr2 node_2 netRa2 -7977.72889578779
Lbr2 netRa2 netL2 6.243602076060146e-12
Rbbr2 netL2 0 25284.66001662448
Cbr2 netL2 0 3.0079883752355076e-20

* Branch 3
Rabr3 node_2 netRa3 -4818.99564672139
Lbr3 netRa3 netL3 5.6700536328939745e-12
Rbbr3 netL3 0 27851.095478736104
Cbr3 netL3 0 4.05042976461503e-20

* Branch 4
Rabr4 node_2 netRa4 14228.699023584213
Lbr4 netRa4 netL4 1.411924753752371e-11
Rbbr4 netL4 0 -23832.884821574913
Cbr4 netL4 0 4.2875247257943557e-20

* Branch 5
Rabr5 node_2 netRa5 17451.626678281496
Lbr5 netRa5 netL5 1.5545137292424016e-11
Rbbr5 netL5 0 -26891.588004222758
Cbr5 netL5 0 3.398424747493512e-20

* Branch 6
Rabr6 node_2 netRa6 9045509.902802862
Lbr6 netRa6 netL6 3.623378964022966e-10
Rbbr6 netL6 0 -9095028.840168996
Cbr6 netL6 0 4.408930208227926e-24

* Branch 7
Rabr7 node_2 netRa7 289619.5895417319
Lbr7 netRa7 netL7 -1.5741376627058912e-10
Rbbr7 netL7 0 -440511.43977968895
Cbr7 netL7 0 -1.2172595485822826e-21

* Branch 8
Rabr8 node_2 netRa8 -241434.4518808359
Lbr8 netRa8 netL8 8.040024988757858e-11
Rbbr8 netL8 0 319723.3116641046
Cbr8 netL8 0 1.033031451529498e-21

* Branch 9
Rabr9 node_2 netRa9 205645.10492818803
Lbr9 netRa9 netL9 4.774390391167928e-11
Rbbr9 netL9 0 -239554.66993198192
Cbr9 netL9 0 9.747343723184895e-22

* Branch 10
Rabr10 node_2 netRa10 -8419.375534421952
Lbr10 netRa10 netL10 -1.0434009269978508e-11
Rbbr10 netL10 0 19433.21183486891
Cbr10 netL10 0 -6.576285682361671e-20

* Branch 11
Rabr11 node_2 netRa11 3590543.9549645223
Lbr11 netRa11 netL11 3.491045941941169e-10
Rbbr11 netL11 0 -3680710.6630828334
Cbr11 netL11 0 2.6478476040902604e-23

* Branch 12
Rabr12 node_2 netRa12 2232714.6774916365
Lbr12 netRa12 netL12 -3.8983647775644206e-10
Rbbr12 netL12 0 -2369119.189353684
Cbr12 netL12 0 -7.338796513639682e-23

* Branch 13
Rabr13 node_2 netRa13 23026.56757238416
Lbr13 netRa13 netL13 2.7019023273773365e-11
Rbbr13 netL13 0 -107630.75413062218
Cbr13 netL13 0 1.1219858200112827e-20

* Branch 14
Rabr14 node_2 netRa14 29617.544006114742
Lbr14 netRa14 netL14 1.786972968205445e-11
Rbbr14 netL14 0 -36887.802449604445
Cbr14 netL14 0 1.6589616788873634e-20

* Branch 15
Rabr15 node_2 netRa15 25509.216668305064
Lbr15 netRa15 netL15 2.5158536295068254e-11
Rbbr15 netL15 0 -86367.0876609256
Cbr15 netL15 0 1.1686925247911864e-20

* Branch 16
Rabr16 node_2 netRa16 1093.02781621451
Lbr16 netRa16 netL16 5.733121572675713e-12
Rbbr16 netL16 0 -113238.18040096092
Cbr16 netL16 0 5.2567715653455955e-20

* Branch 17
Rabr17 node_2 netRa17 -69027.55443058934
Lbr17 netRa17 netL17 4.8863692882048845e-11
Rbbr17 netL17 0 153989.38251606288
Cbr17 netL17 0 4.525554917588804e-21

* Branch 18
Rabr18 node_2 netRa18 -15861.260252111175
Lbr18 netRa18 netL18 2.390091464280197e-11
Rbbr18 netL18 0 104797.26052340513
Cbr18 netL18 0 1.3917354750361618e-20

* Branch 19
Rabr19 node_2 netRa19 -278009.5469605858
Lbr19 netRa19 netL19 1.0566500203093206e-10
Rbbr19 netL19 0 350968.8423764065
Cbr19 netL19 0 1.0740234168618883e-21

* Branch 20
Rabr20 node_2 netRa20 90160.33698274646
Lbr20 netRa20 netL20 -2.3500698454294464e-11
Rbbr20 netL20 0 -110358.2691292007
Cbr20 netL20 0 -2.3491035255978775e-21

* Branch 21
Rabr21 node_2 netRa21 6386070.106806639
Lbr21 netRa21 netL21 -3.9644316017440353e-10
Rbbr21 netL21 0 -6456340.5261456575
Cbr21 netL21 0 -9.602834297095814e-24

* Branch 22
Rabr22 node_2 netRa22 215730.26756754916
Lbr22 netRa22 netL22 -1.222888426618367e-10
Rbbr22 netL22 0 -313049.0207104292
Cbr22 netL22 0 -1.7896457907531052e-21

* Branch 23
Rabr23 node_2 netRa23 2025754.614100569
Lbr23 netRa23 netL23 -3.279931087230927e-10
Rbbr23 netL23 0 -2133118.000881349
Cbr23 netL23 0 -7.565449957501851e-23

* Branch 24
Rabr24 node_2 netRa24 -107723.28190868397
Lbr24 netRa24 netL24 -7.165194600173611e-11
Rbbr24 netL24 0 171830.40291836875
Cbr24 netL24 0 -3.923615996901048e-21

* Branch 25
Rabr25 node_2 netRa25 -88043.71800502049
Lbr25 netRa25 netL25 5.2038555197357114e-11
Rbbr25 netL25 0 136066.78327083125
Cbr25 netL25 0 4.293940406514587e-21

* Branch 26
Rabr26 node_2 netRa26 6350.671327808842
Lbr26 netRa26 netL26 3.482734694369558e-11
Rbbr26 netL26 0 -382593.8975829844
Cbr26 netL26 0 1.6061138151280975e-20

* Branch 27
Rabr27 node_2 netRa27 1635677.148612561
Lbr27 netRa27 netL27 1.5588425811823267e-10
Rbbr27 netL27 0 -1676288.872890404
Cbr27 netL27 0 5.695901990676108e-23

* Branch 28
Rabr28 node_2 netRa28 104686.13496265377
Lbr28 netRa28 netL28 3.04171255678123e-11
Rbbr28 netL28 0 -110590.30630411353
Cbr28 netL28 0 2.6420992229146896e-21

* Branch 29
Rabr29 node_2 netRa29 -630621.6812225307
Lbr29 netRa29 netL29 1.5115422819732065e-10
Rbbr29 netL29 0 690978.5275935852
Cbr29 netL29 0 3.45305009802027e-22

* Branch 30
Rabr30 node_2 netRa30 -15732.812917343173
Lbr30 netRa30 netL30 2.0694695868259534e-11
Rbbr30 netL30 0 91340.4560445402
Cbr30 netL30 0 1.4052011583275188e-20

* Branch 31
Rabr31 node_2 netRa31 118153.76813473862
Lbr31 netRa31 netL31 6.640390806697029e-11
Rbbr31 netL31 0 -175015.93932280858
Cbr31 netL31 0 3.245056684131243e-21

* Branch 32
Rabr32 node_2 netRa32 211651.1368038956
Lbr32 netRa32 netL32 1.017244550980638e-10
Rbbr32 netL32 0 -293238.81944275537
Cbr32 netL32 0 1.6532385402968564e-21

* Branch 33
Rabr33 node_2 netRa33 -29252.290618934865
Lbr33 netRa33 netL33 4.365890224268558e-11
Rbbr33 netL33 0 138196.4471018774
Cbr33 netL33 0 1.053356898471309e-20

* Branch 34
Rabr34 node_2 netRa34 -30117.073489711118
Lbr34 netRa34 netL34 3.930869190977862e-11
Rbbr34 netL34 0 124146.82994363575
Cbr34 netL34 0 1.0286947452729746e-20

* Branch 35
Rabr35 node_2 netRa35 5242.687568844133
Lbr35 netRa35 netL35 3.793512277762576e-11
Rbbr35 netL35 0 -505070.8140363556
Cbr35 netL35 0 1.6210108628127063e-20

* Branch 36
Rabr36 node_2 netRa36 70996.43078846685
Lbr36 netRa36 netL36 4.546462054671932e-11
Rbbr36 netL36 0 -137517.592257891
Cbr36 netL36 0 4.705060229906082e-21

* Branch 37
Rabr37 node_2 netRa37 1138642.5744818747
Lbr37 netRa37 netL37 -3.6511441903087115e-10
Rbbr37 netL37 0 -1367065.4708951123
Cbr37 netL37 0 -2.333685635682965e-22

* Branch 38
Rabr38 node_2 netRa38 38328.82887908201
Lbr38 netRa38 netL38 5.2483540624228784e-11
Rbbr38 netL38 0 -197392.33008528786
Cbr38 netL38 0 7.08611031127771e-21

* Branch 39
Rabr39 node_2 netRa39 -2201754.6010060357
Lbr39 netRa39 netL39 -4.670218882473561e-10
Rbbr39 netL39 0 2355094.953924008
Cbr39 netL39 0 -9.036020012661909e-23

* Branch 40
Rabr40 node_2 netRa40 -5990530.4171849135
Lbr40 netRa40 netL40 2.30290711329908e-10
Rbbr40 netL40 0 5996054.904009057
Cbr40 netL40 0 6.407534337957581e-24

* Branch 41
Rabr41 node_2 netRa41 -1939297.601126092
Lbr41 netRa41 netL41 -1.6434844723376687e-10
Rbbr41 netL41 0 1947520.4072852265
Cbr41 netL41 0 -4.3571152876218827e-23

* Branch 42
Rabr42 node_2 netRa42 -27990.769861540404
Lbr42 netRa42 netL42 1.94923806336261e-11
Rbbr42 netL42 0 71389.93793751372
Cbr42 netL42 0 9.653412785053385e-21

* Branch 43
Rabr43 node_2 netRa43 35989.474881461225
Lbr43 netRa43 netL43 -6.475619708310072e-11
Rbbr43 netL43 0 -172850.02817904457
Cbr43 netL43 0 -1.0140284989053362e-20

* Branch 44
Rabr44 node_2 netRa44 -69174.02789355212
Lbr44 netRa44 netL44 3.381186612867519e-11
Rbbr44 netL44 0 121177.82830163295
Cbr44 netL44 0 4.006529765549788e-21

* Branch 45
Rabr45 node_2 netRa45 47370.989214229194
Lbr45 netRa45 netL45 4.479256156232327e-11
Rbbr45 netL45 0 -103080.30445799103
Cbr45 netL45 0 9.28843391562052e-21

* Branch 46
Rabr46 node_2 netRa46 -29880.350682769167
Lbr46 netRa46 netL46 3.5310744677458345e-11
Rbbr46 netL46 0 80554.84072170759
Cbr46 netL46 0 1.4454690375158363e-20

* Branch 47
Rabr47 node_2 netRa47 -29503.968586593284
Lbr47 netRa47 netL47 1.0590896229632808e-10
Rbbr47 netL47 0 919458.3021173957
Cbr47 netL47 0 3.7420248095813174e-21

* Branch 48
Rabr48 node_2 netRa48 -66152.60152253653
Lbr48 netRa48 netL48 3.0590237586828114e-11
Rbbr48 netL48 0 108268.08030393919
Cbr48 netL48 0 4.247472686039712e-21

* Branch 49
Rabr49 node_2 netRa49 -325165.3723599258
Lbr49 netRa49 netL49 8.858586368954969e-11
Rbbr49 netL49 0 389664.27286347374
Cbr49 netL49 0 6.9688158990436415e-22

* Branch 50
Rabr50 node_2 netRa50 -16147.492074012189
Lbr50 netRa50 netL50 3.75762568347664e-11
Rbbr50 netL50 0 131581.701466491
Cbr50 netL50 0 1.7221303132570612e-20

* Branch 51
Rabr51 node_2 netRa51 2809.2890005806535
Lbr51 netRa51 netL51 -2.7435507506144148e-11
Rbbr51 netL51 0 -843578.5863841209
Cbr51 netL51 0 -1.0411928617324907e-20

* Branch 52
Rabr52 node_2 netRa52 -19707.21812426017
Lbr52 netRa52 netL52 -1.8035575587809476e-11
Rbbr52 netL52 0 29055.61831013956
Cbr52 netL52 0 -3.18184442216756e-20

* Branch 53
Rabr53 node_2 netRa53 -14895.82149680941
Lbr53 netRa53 netL53 3.8381175790334363e-11
Rbbr53 netL53 0 157678.11985914095
Cbr53 netL53 0 1.589055385554629e-20

* Branch 54
Rabr54 node_2 netRa54 -89218.08795116251
Lbr54 netRa54 netL54 5.053732774679319e-11
Rbbr54 netL54 0 177462.87187576812
Cbr54 netL54 0 3.172676651914172e-21

* Branch 55
Rabr55 node_2 netRa55 -64152.863927894614
Lbr55 netRa55 netL55 6.127624764636462e-11
Rbbr55 netL55 0 147876.82028166926
Cbr55 netL55 0 6.394320727902977e-21

* Branch 56
Rabr56 node_2 netRa56 -40997.82278004625
Lbr56 netRa56 netL56 4.4143729292988836e-11
Rbbr56 netL56 0 93413.15289757452
Cbr56 netL56 0 1.1397858956704284e-20

* Branch 57
Rabr57 node_2 netRa57 -60307.07320968219
Lbr57 netRa57 netL57 5.593586133880517e-11
Rbbr57 netL57 0 180033.3608646875
Cbr57 netL57 0 5.1043291047855534e-21

* Branch 58
Rabr58 node_2 netRa58 -2821.7053612520895
Lbr58 netRa58 netL58 -1.0273374623659823e-11
Rbbr58 netL58 0 29602.23606359252
Cbr58 netL58 0 -1.2764433701337607e-19

* Branch 59
Rabr59 node_2 netRa59 -100441.6166712099
Lbr59 netRa59 netL59 7.238662822502002e-11
Rbbr59 netL59 0 244874.91671125256
Cbr59 netL59 0 2.922177470850534e-21

* Branch 60
Rabr60 node_2 netRa60 -18953.60731926855
Lbr60 netRa60 netL60 4.0904364637334075e-11
Rbbr60 netL60 0 184869.12049970767
Cbr60 netL60 0 1.142939941357146e-20

* Branch 61
Rabr61 node_2 netRa61 5337.184953607608
Lbr61 netRa61 netL61 3.8310823258473583e-11
Rbbr61 netL61 0 -418369.8549539818
Cbr61 netL61 0 1.8469185641962474e-20

* Branch 62
Rabr62 node_2 netRa62 16543.758962796768
Lbr62 netRa62 netL62 2.2446849767298644e-11
Rbbr62 netL62 0 -31518.63244474754
Cbr62 netL62 0 4.3604959447157824e-20

* Branch 63
Rabr63 node_2 netRa63 1317.453767924901
Lbr63 netRa63 netL63 -2.7481321495406002e-11
Rbbr63 netL63 0 -494632.7506275416
Cbr63 netL63 0 -3.562270563650581e-20

* Branch 64
Rabr64 node_2 netRa64 -17910130.37761763
Lbr64 netRa64 netL64 3.0796323346691744e-10
Rbbr64 netL64 0 17913591.590944704
Cbr64 netL64 0 9.597410830526673e-25

* Branch 65
Rabr65 node_2 netRa65 -295947.5045503996
Lbr65 netRa65 netL65 9.814938193967953e-11
Rbbr65 netL65 0 366442.1243051349
Cbr65 netL65 0 9.026894794951446e-22

* Branch 66
Rabr66 node_2 netRa66 4603.671982425594
Lbr66 netRa66 netL66 3.1521453680921435e-11
Rbbr66 netL66 0 -293953.1382565048
Cbr66 netL66 0 2.4608602611337437e-20

* Branch 67
Rabr67 node_2 netRa67 -5997.2978362877475
Lbr67 netRa67 netL67 3.955014378078254e-11
Rbbr67 netL67 0 121601.32611198742
Cbr67 netL67 0 5.163392300271903e-20

* Branch 68
Rabr68 node_2 netRa68 -503436.3142265462
Lbr68 netRa68 netL68 -3.061754200765954e-10
Rbbr68 netL68 0 583491.4901368925
Cbr68 netL68 0 -1.0468309283479075e-21

* Branch 69
Rabr69 node_2 netRa69 -76773.88142544877
Lbr69 netRa69 netL69 7.530764462094532e-11
Rbbr69 netL69 0 243271.14686323475
Cbr69 netL69 0 4.005221953177449e-21

* Branch 70
Rabr70 node_2 netRa70 -170632.96497293594
Lbr70 netRa70 netL70 9.200016279171206e-11
Rbbr70 netL70 0 288449.86972036184
Cbr70 netL70 0 1.8623831374475087e-21

* Branch 71
Rabr71 node_2 netRa71 -161702.4877933815
Lbr71 netRa71 netL71 8.05690658348632e-11
Rbbr71 netL71 0 270926.80200490815
Cbr71 netL71 0 1.833407167854537e-21

* Branch 72
Rabr72 node_2 netRa72 -228005.40324630606
Lbr72 netRa72 netL72 1.6391352096775465e-10
Rbbr72 netL72 0 280238.7967515339
Cbr72 netL72 0 2.5540853742202397e-21

* Branch 73
Rabr73 node_2 netRa73 -2336.8312139593495
Lbr73 netRa73 netL73 -2.1506310404309496e-11
Rbbr73 netL73 0 746671.8262605068
Cbr73 netL73 0 -1.304449206567612e-20

* Branch 74
Rabr74 node_2 netRa74 688400.5961358226
Lbr74 netRa74 netL74 -9.529054780215416e-11
Rbbr74 netL74 0 -695067.1698550556
Cbr74 netL74 0 -1.9899832375569606e-22

* Branch 75
Rabr75 node_2 netRa75 -5432.314404385455
Lbr75 netRa75 netL75 6.206262235770123e-11
Rbbr75 netL75 0 1424561.6708454604
Cbr75 netL75 0 7.600058837558146e-21

* Branch 76
Rabr76 node_2 netRa76 -1405.3960986194083
Lbr76 netRa76 netL76 -2.164147758418827e-11
Rbbr76 netL76 0 195994.01831476047
Cbr76 netL76 0 -8.484668295103408e-20

* Branch 77
Rabr77 node_2 netRa77 -6432062.703771918
Lbr77 netRa77 netL77 -5.428948801937841e-10
Rbbr77 netL77 0 6475025.5242295
Cbr77 netL77 0 -1.3040132730719889e-23

* Branch 78
Rabr78 node_2 netRa78 21136.2297004179
Lbr78 netRa78 netL78 2.6849718614261568e-11
Rbbr78 netL78 0 -61665.59228909743
Cbr78 netL78 0 2.0711768930433184e-20

* Branch 79
Rabr79 node_2 netRa79 342077.6474726639
Lbr79 netRa79 netL79 8.765860232209966e-11
Rbbr79 netL79 0 -366841.6054423627
Cbr79 netL79 0 6.991386046019321e-22

* Branch 80
Rabr80 node_2 netRa80 68085.68255053791
Lbr80 netRa80 netL80 -3.458814933190527e-11
Rbbr80 netL80 0 -77240.8674777992
Cbr80 netL80 0 -6.566117570528121e-21

* Branch 81
Rabr81 node_2 netRa81 -484144.8629502043
Lbr81 netRa81 netL81 1.1875582986619513e-10
Rbbr81 netL81 0 541540.9935829546
Cbr81 netL81 0 4.527066616844908e-22

* Branch 82
Rabr82 node_2 netRa82 -1854058.5766417035
Lbr82 netRa82 netL82 3.3482136160715625e-10
Rbbr82 netL82 0 1975886.5822371594
Cbr82 netL82 0 9.137506466587064e-23

* Branch 83
Rabr83 node_2 netRa83 -130258.60699924346
Lbr83 netRa83 netL83 2.3937496859400413e-10
Rbbr83 netL83 0 1035928.3917870374
Cbr83 netL83 0 1.770218749279439e-21

* Branch 84
Rabr84 node_2 netRa84 38292.56359112642
Lbr84 netRa84 netL84 -1.374340088067537e-10
Rbbr84 netL84 0 -401657.25827820343
Cbr84 netL84 0 -8.899516032996776e-21

* Branch 85
Rabr85 node_2 netRa85 37178.30078314124
Lbr85 netRa85 netL85 4.156371456489172e-11
Rbbr85 netL85 0 -90820.71406920487
Cbr85 netL85 0 1.2324675311691079e-20

* Branch 86
Rabr86 node_2 netRa86 96640.42822868044
Lbr86 netRa86 netL86 1.6499870662133844e-10
Rbbr86 netL86 0 -722935.536306947
Cbr86 netL86 0 2.3657443663798137e-21

* Branch 87
Rabr87 node_2 netRa87 -44854252.895660274
Lbr87 netRa87 netL87 1.4078864709183367e-09
Rbbr87 netL87 0 44988504.84217238
Cbr87 netL87 0 6.9767189241892715e-25

* Branch 88
Rabr88 node_2 netRa88 18706054.23737524
Lbr88 netRa88 netL88 6.112057224971898e-10
Rbbr88 netL88 0 -18724716.26088273
Cbr88 netL88 0 1.7449932680816087e-24

* Branch 89
Rabr89 node_2 netRa89 65946.31770013503
Lbr89 netRa89 netL89 -6.4992829616678e-11
Rbbr89 netL89 0 -117327.31958735122
Cbr89 netL89 0 -8.397606685202462e-21

* Branch 90
Rabr90 node_2 netRa90 114151.33924262803
Lbr90 netRa90 netL90 8.766019964600652e-11
Rbbr90 netL90 0 -179645.90724463342
Cbr90 netL90 0 4.27571947619857e-21

* Branch 91
Rabr91 node_2 netRa91 260523.4287458366
Lbr91 netRa91 netL91 1.0887176162077325e-10
Rbbr91 netL91 0 -300058.4136218363
Cbr91 netL91 0 1.3929226348914559e-21

* Branch 92
Rabr92 node_2 netRa92 1183610.360752553
Lbr92 netRa92 netL92 2.0794082976815175e-10
Rbbr92 netL92 0 -1214148.958327801
Cbr92 netL92 0 1.4470705185946979e-22

* Branch 93
Rabr93 node_2 netRa93 5728.649097471045
Lbr93 netRa93 netL93 -2.1841871926118228e-11
Rbbr93 netL93 0 -69297.75261382626
Cbr93 netL93 0 -5.492871762343111e-20

* Branch 94
Rabr94 node_2 netRa94 173282.3941068957
Lbr94 netRa94 netL94 1.0985074865271308e-10
Rbbr94 netL94 0 -236211.60157329726
Cbr94 netL94 0 2.6847301460720734e-21

* Branch 95
Rabr95 node_2 netRa95 19150.869851410447
Lbr95 netRa95 netL95 3.163377795733571e-11
Rbbr95 netL95 0 -73703.58360814072
Cbr95 netL95 0 2.2457501544934303e-20

* Branch 96
Rabr96 node_2 netRa96 26146.863614544585
Lbr96 netRa96 netL96 2.852086115630803e-11
Rbbr96 netL96 0 -59693.053873572004
Cbr96 netL96 0 1.8300603999541524e-20

* Branch 97
Rabr97 node_2 netRa97 54748.737638902945
Lbr97 netRa97 netL97 3.5176222496313846e-11
Rbbr97 netL97 0 -77477.01984003316
Cbr97 netL97 0 8.3032509743407e-21

* Branch 98
Rabr98 node_2 netRa98 17747.11567493235
Lbr98 netRa98 netL98 1.4434982790285555e-11
Rbbr98 netL98 0 -25733.21247103876
Cbr98 netL98 0 3.227926816194977e-20

* Branch 99
Rabr99 node_2 netRa99 -4164.52955107727
Lbr99 netRa99 netL99 5.771277601666088e-12
Rbbr99 netL99 0 31312.23619743734
Cbr99 netL99 0 4.193668733424415e-20

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 3855534.5390559984
Lbr0 netRa0 netL0 -2.768553400814807e-10
Rbbr0 netL0 node_3 -3917425.2189643895
Cbr0 netL0 node_3 -1.8241998161676092e-23

* Branch 1
Rabr1 node_2 netRa1 1027658.3883831204
Lbr1 netRa1 netL1 -1.7725718907512156e-10
Rbbr1 netL1 node_3 -1109492.1347499876
Cbr1 netL1 node_3 -1.5382498761586122e-22

* Branch 2
Rabr2 node_2 netRa2 3167441.900371965
Lbr2 netRa2 netL2 -2.429704489465672e-10
Rbbr2 netL2 node_3 -3226089.308057045
Cbr2 netL2 node_3 -2.3679303717293374e-23

* Branch 3
Rabr3 node_2 netRa3 787693.3157951123
Lbr3 netRa3 netL3 -1.496374951474356e-10
Rbbr3 netL3 node_3 -864734.4798609456
Cbr3 netL3 node_3 -2.1788836984273395e-22

* Branch 4
Rabr4 node_2 netRa4 3952085.959406826
Lbr4 netRa4 netL4 -2.6026399580672645e-10
Rbbr4 netL4 node_3 -4006989.497636566
Cbr4 netL4 node_3 -1.6393022004342992e-23

* Branch 5
Rabr5 node_2 netRa5 1434871.9871936047
Lbr5 netRa5 netL5 -1.659465066205275e-10
Rbbr5 netL5 node_3 -1494686.567534655
Cbr5 netL5 node_3 -7.703643609287871e-23

* Branch 6
Rabr6 node_2 netRa6 582590.1869176343
Lbr6 netRa6 netL6 -1.3299792038067792e-10
Rbbr6 netL6 node_3 -664157.8522063969
Cbr6 netL6 node_3 -3.413061251097782e-22

* Branch 7
Rabr7 node_2 netRa7 3869120.352397914
Lbr7 netRa7 netL7 -2.554861418103259e-10
Rbbr7 netL7 node_3 -3924639.346299186
Cbr7 netL7 node_3 -1.679206479547739e-23

* Branch 8
Rabr8 node_2 netRa8 264558.1823657107
Lbr8 netRa8 netL8 -2.6009861807648275e-10
Rbbr8 netL8 node_3 -510758.06398508063
Cbr8 netL8 node_3 -1.893296649294846e-21

* Branch 9
Rabr9 node_2 netRa9 282828.48315785377
Lbr9 netRa9 netL9 -2.538290250574165e-10
Rbbr9 netL9 node_3 -521008.9357704569
Cbr9 netL9 node_3 -1.6970571927185907e-21

* Branch 10
Rabr10 node_2 netRa10 246888.4241473142
Lbr10 netRa10 netL10 -2.6614854826144446e-10
Rbbr10 netL10 node_3 -500641.8018952006
Cbr10 netL10 node_3 -2.1154286487836445e-21

* Branch 11
Rabr11 node_2 netRa11 229127.92121926232
Lbr11 netRa11 netL11 -2.717920897143158e-10
Rbbr11 netL11 node_3 -490108.8974195187
Cbr11 netL11 node_3 -2.3753372887092207e-21

* Branch 12
Rabr12 node_2 netRa12 301737.68595835083
Lbr12 netRa12 netL12 -2.4767678384190585e-10
Rbbr12 netL12 node_3 -531834.814453682
Cbr12 netL12 node_3 -1.523764007066329e-21

* Branch 13
Rabr13 node_2 netRa13 211384.15103734194
Lbr13 netRa13 netL13 -2.772460764845006e-10
Rbbr13 netL13 node_3 -479465.1573590913
Cbr13 netL13 node_3 -2.6821180395974796e-21

* Branch 14
Rabr14 node_2 netRa14 369301.0076668889
Lbr14 netRa14 netL14 -1.553663631316704e-10
Rbbr14 netL14 node_3 -511462.583798412
Cbr14 netL14 node_3 -8.175334620857625e-22

* Branch 15
Rabr15 node_2 netRa15 193732.94383348597
Lbr15 netRa15 netL15 -2.8253074350374573e-10
Rbbr15 netL15 node_3 -468739.3105882432
Cbr15 netL15 node_3 -3.047119431073302e-21

* Branch 16
Rabr16 node_2 netRa16 176357.3298435496
Lbr16 netRa16 netL16 -2.8771473370486867e-10
Rbbr16 netL16 node_3 -458168.4823197428
Cbr16 netL16 node_3 -3.4823272025923484e-21

* Branch 17
Rabr17 node_2 netRa17 319417.818423598
Lbr17 netRa17 netL17 -2.421393283177458e-10
Rbbr17 netL17 node_3 -542382.959558406
Cbr17 netL17 node_3 -1.3832108325600326e-21

* Branch 18
Rabr18 node_2 netRa18 386381.71087692695
Lbr18 netRa18 netL18 -1.6633240506544715e-10
Rbbr18 netL18 node_3 -537566.0947137213
Cbr18 netL18 node_3 -7.961115745372088e-22

* Branch 19
Rabr19 node_2 netRa19 330921.15272071416
Lbr19 netRa19 netL19 -2.333124484472814e-10
Rbbr19 netL19 node_3 -546600.768701445
Cbr19 netL19 node_3 -1.2776059998611854e-21

* Branch 20
Rabr20 node_2 netRa20 159455.477760623
Lbr20 netRa20 netL20 -2.928591547828014e-10
Rbbr20 netL20 node_3 -447944.3148310389
Cbr20 netL20 node_3 -4.002604448310438e-21

* Branch 21
Rabr21 node_2 netRa21 359048.01186705113
Lbr21 netRa21 netL21 -2.2683272128421145e-10
Rbbr21 netL21 node_3 -561842.4301463082
Cbr21 netL21 node_3 -1.1154593268144343e-21

* Branch 22
Rabr22 node_2 netRa22 143322.38968107064
Lbr22 netRa22 netL22 -2.9845111796637146e-10
Rbbr22 netL22 node_3 -438150.714623575
Cbr22 netL22 node_3 -4.631574064489863e-21

* Branch 23
Rabr23 node_2 netRa23 428130.3573620831
Lbr23 netRa23 netL23 -1.406811441564591e-10
Rbbr23 netL23 node_3 -539436.8295403848
Cbr23 netL23 node_3 -6.070004633014185e-22

* Branch 24
Rabr24 node_2 netRa24 425766.9000862392
Lbr24 netRa24 netL24 -1.938872734304673e-10
Rbbr24 netL24 node_3 -593470.1740320129
Cbr24 netL24 node_3 -7.637527913518535e-22

* Branch 25
Rabr25 node_2 netRa25 577645.5311439473
Lbr25 netRa25 netL25 -1.5177106586279516e-10
Rbbr25 netL25 node_3 -678882.5569018935
Cbr25 netL25 node_3 -3.8599076929431346e-22

* Branch 26
Rabr26 node_2 netRa26 449870.05557774147
Lbr26 netRa26 netL26 -2.062259787979896e-10
Rbbr26 netL26 node_3 -618880.6831006706
Cbr26 netL26 node_3 -7.375299628252134e-22

* Branch 27
Rabr27 node_2 netRa27 462799.0566539518
Lbr27 netRa27 netL27 -1.879676997267184e-10
Rbbr27 netL27 node_3 -619744.2341229189
Cbr27 netL27 node_3 -6.528887349687967e-22

* Branch 28
Rabr28 node_2 netRa28 352456.5884110142
Lbr28 netRa28 netL28 -2.1466101337253622e-10
Rbbr28 netL28 node_3 -550339.1920615223
Cbr28 netL28 node_3 -1.1020928523841069e-21

* Branch 29
Rabr29 node_2 netRa29 392623.9518586359
Lbr29 netRa29 netL29 -2.0117413076552826e-10
Rbbr29 netL29 node_3 -561326.1328655308
Cbr29 netL29 node_3 -9.100501087513107e-22

* Branch 30
Rabr30 node_2 netRa30 -52544.517469585684
Lbr30 netRa30 netL30 -1.2318007256879038e-10
Rbbr30 netL30 node_3 889607.5752424805
Cbr30 netL30 node_3 -2.6562350316555968e-21

* Branch 31
Rabr31 node_2 netRa31 2329224.510360476
Lbr31 netRa31 netL31 -7.244784219028489e-10
Rbbr31 netL31 node_3 -3099784.4474394945
Cbr31 netL31 node_3 -1.002390858787466e-22

* Branch 32
Rabr32 node_2 netRa32 -369922.7012846304
Lbr32 netRa32 netL32 4.978672958222322e-09
Rbbr32 netL32 node_3 118402619.36997792
Cbr32 netL32 node_3 1.1341580892908091e-22

* Branch 33
Rabr33 node_2 netRa33 88966438.35063088
Lbr33 netRa33 netL33 -1.4455288866397744e-08
Rbbr33 netL33 node_3 -92675606.31615847
Cbr33 netL33 node_3 -1.7531797027924785e-24

* Branch 34
Rabr34 node_2 netRa34 43870579.70890216
Lbr34 netRa34 netL34 1.3758249721698125e-08
Rbbr34 netL34 node_3 -50882049.94343101
Cbr34 netL34 node_3 6.163631011122012e-24

* Branch 35
Rabr35 node_2 netRa35 -3085884.041819407
Lbr35 netRa35 netL35 3.1884807384133672e-09
Rbbr35 netL35 node_3 5333244.133426685
Cbr35 netL35 node_3 1.9373695547131401e-22

* Branch 36
Rabr36 node_2 netRa36 -349090.97783354914
Lbr36 netRa36 netL36 2.190688766568617e-09
Rbbr36 netL36 node_3 9323681.615786256
Cbr36 netL36 node_3 6.730578226480014e-22

* Branch 37
Rabr37 node_2 netRa37 2007489.68846769
Lbr37 netRa37 netL37 2.715710633688699e-09
Rbbr37 netL37 node_3 -4623737.303290927
Cbr37 netL37 node_3 2.9257542310799e-22

* Branch 38
Rabr38 node_2 netRa38 479439.4426093887
Lbr38 netRa38 netL38 2.183685625297156e-09
Rbbr38 netL38 node_3 -6687060.413569229
Cbr38 netL38 node_3 6.811234873563926e-22

* Branch 39
Rabr39 node_2 netRa39 1091353.3971643816
Lbr39 netRa39 netL39 2.3425967981611853e-09
Rbbr39 netL39 node_3 -4826294.543214483
Cbr39 netL39 node_3 4.44756051486576e-22

* Branch 40
Rabr40 node_2 netRa40 944503.9318710085
Lbr40 netRa40 netL40 2.5071338990818033e-09
Rbbr40 netL40 node_3 -4911494.21363433
Cbr40 netL40 node_3 5.404621356797844e-22

* Branch 41
Rabr41 node_2 netRa41 1401341.285934615
Lbr41 netRa41 netL41 2.3408038058099123e-09
Rbbr41 netL41 node_3 -4427906.404421294
Cbr41 netL41 node_3 3.7724853856906745e-22

* Branch 42
Rabr42 node_2 netRa42 983315.073033693
Lbr42 netRa42 netL42 2.4952763420734013e-09
Rbbr42 netL42 node_3 -4584275.026348359
Cbr42 netL42 node_3 5.535588266029944e-22

* Branch 43
Rabr43 node_2 netRa43 1465511.4024219331
Lbr43 netRa43 netL43 2.389813353665228e-09
Rbbr43 netL43 node_3 -4606391.822016031
Cbr43 netL43 node_3 3.540140433441577e-22

* Branch 44
Rabr44 node_2 netRa44 925420.6622445589
Lbr44 netRa44 netL44 2.589279818125671e-09
Rbbr44 netL44 node_3 -4851559.963910878
Cbr44 netL44 node_3 5.767291193925231e-22

* Branch 45
Rabr45 node_2 netRa45 1644384.8168230425
Lbr45 netRa45 netL45 2.320755260650893e-09
Rbbr45 netL45 node_3 -4390811.304929976
Cbr45 netL45 node_3 3.214317464655186e-22

* Branch 46
Rabr46 node_2 netRa46 1441793.4752737554
Lbr46 netRa46 netL46 2.2681755804515344e-09
Rbbr46 netL46 node_3 -4552301.333798611
Cbr46 netL46 node_3 3.4558321764981216e-22

* Branch 47
Rabr47 node_2 netRa47 961325.4372517179
Lbr47 netRa47 netL47 2.608183486584631e-09
Rbbr47 netL47 node_3 -4611449.278033066
Cbr47 netL47 node_3 5.883664815432448e-22

* Branch 48
Rabr48 node_2 netRa48 1536711.8033412956
Lbr48 netRa48 netL48 2.188710247331262e-09
Rbbr48 netL48 node_3 -4359708.811259575
Cbr48 netL48 node_3 3.267005643176893e-22

* Branch 49
Rabr49 node_2 netRa49 721488.8964303071
Lbr49 netRa49 netL49 2.473028948445933e-09
Rbbr49 netL49 node_3 -4878208.8469341975
Cbr49 netL49 node_3 7.0269788035873205e-22

* Branch 50
Rabr50 node_2 netRa50 1897197.165209718
Lbr50 netRa50 netL50 2.3258609313789153e-09
Rbbr50 netL50 node_3 -4577693.556633918
Cbr50 netL50 node_3 2.678153951502466e-22

* Branch 51
Rabr51 node_2 netRa51 778587.0849346998
Lbr51 netRa51 netL51 2.647629041838724e-09
Rbbr51 netL51 node_3 -4970086.467010761
Cbr51 netL51 node_3 6.842564699998781e-22

* Branch 52
Rabr52 node_2 netRa52 1380717.5433758474
Lbr52 netRa52 netL52 2.0839165521123845e-09
Rbbr52 netL52 node_3 -4448039.407266952
Cbr52 netL52 node_3 3.393309641848041e-22

* Branch 53
Rabr53 node_2 netRa53 648003.4095774479
Lbr53 netRa53 netL53 2.6031997948761862e-09
Rbbr53 netL53 node_3 -5263814.773948638
Cbr53 netL53 node_3 7.63264610023309e-22

* Branch 54
Rabr54 node_2 netRa54 1710765.625260427
Lbr54 netRa54 netL54 2.1481680525959527e-09
Rbbr54 netL54 node_3 -4437840.762732391
Cbr54 netL54 node_3 2.8295789909850904e-22

* Branch 55
Rabr55 node_2 netRa55 550569.2801013441
Lbr55 netRa55 netL55 2.586019704394363e-09
Rbbr55 netL55 node_3 -5626044.445816277
Cbr55 netL55 node_3 8.349795363080497e-22

* Branch 56
Rabr56 node_2 netRa56 343353.63490517554
Lbr56 netRa56 netL56 2.5334989363358064e-09
Rbbr56 netL56 node_3 -7727501.85363021
Cbr56 netL56 node_3 9.550875949720255e-22

* Branch 57
Rabr57 node_2 netRa57 1505846.2058002008
Lbr57 netRa57 netL57 2.074468162788595e-09
Rbbr57 netL57 node_3 -4499226.943622804
Cbr57 netL57 node_3 3.062026979338248e-22

* Branch 58
Rabr58 node_2 netRa58 1747018.8024539144
Lbr58 netRa58 netL58 2.053367986738068e-09
Rbbr58 netL58 node_3 -4364408.447326983
Cbr58 netL58 node_3 2.6931779219575105e-22

* Branch 59
Rabr59 node_2 netRa59 1979559.7612182528
Lbr59 netRa59 netL59 2.150746770249384e-09
Rbbr59 netL59 node_3 -4601905.013858145
Cbr59 netL59 node_3 2.3610553585880955e-22

* Branch 60
Rabr60 node_2 netRa60 1494903.3286826676
Lbr60 netRa60 netL60 1.8650157129811837e-09
Rbbr60 netL60 node_3 -4195363.400425619
Cbr60 netL60 node_3 2.973943548585079e-22

* Branch 61
Rabr61 node_2 netRa61 1934758.9510649901
Lbr61 netRa61 netL61 2.044781165556672e-09
Rbbr61 netL61 node_3 -4527179.31240751
Cbr61 netL61 node_3 2.334668493433883e-22

* Branch 62
Rabr62 node_2 netRa62 1861159.4834799173
Lbr62 netRa62 netL62 1.9106143092722695e-09
Rbbr62 netL62 node_3 -4291839.691925989
Cbr62 netL62 node_3 2.3921826060117515e-22

* Branch 63
Rabr63 node_2 netRa63 1141382.4457205487
Lbr63 netRa63 netL63 1.7219000784415024e-09
Rbbr63 netL63 node_3 -4465631.939696468
Cbr63 netL63 node_3 3.37900417669098e-22

* Branch 64
Rabr64 node_2 netRa64 983507.1191607948
Lbr64 netRa64 netL64 1.5574431378756315e-09
Rbbr64 netL64 node_3 -4240837.252960527
Cbr64 netL64 node_3 3.7351866191370035e-22

* Branch 65
Rabr65 node_2 netRa65 1326520.6061262705
Lbr65 netRa65 netL65 1.759021783500612e-09
Rbbr65 netL65 node_3 -4504043.626132469
Cbr65 netL65 node_3 2.944903001450727e-22

* Branch 66
Rabr66 node_2 netRa66 12462028.079880644
Lbr66 netRa66 netL66 3.7229248059730725e-09
Rbbr66 netL66 node_3 -14931203.342455462
Cbr66 netL66 node_3 2.0009127531240234e-23

* Branch 67
Rabr67 node_2 netRa67 -2987284.162942476
Lbr67 netRa67 netL67 5.876260986845167e-09
Rbbr67 netL67 node_3 20719718.347261954
Cbr67 netL67 node_3 9.488990513151711e-23

* Branch 68
Rabr68 node_2 netRa68 137205.39731743655
Lbr68 netRa68 netL68 1.3697620190809384e-09
Rbbr68 netL68 node_3 -19391704.064220272
Cbr68 netL68 node_3 5.16226992230503e-22

* Branch 69
Rabr69 node_2 netRa69 -106003315.51214011
Lbr69 netRa69 netL69 1.2115447224288041e-08
Rbbr69 netL69 node_3 108515147.08842807
Cbr69 netL69 node_3 1.0531984914032472e-24

* Branch 70
Rabr70 node_2 netRa70 -510329.0954567078
Lbr70 netRa70 netL70 1.381017457651597e-09
Rbbr70 netL70 node_3 5912783.631746653
Cbr70 netL70 node_3 4.571903257195756e-22

* Branch 71
Rabr71 node_2 netRa71 -86186.02952849404
Lbr71 netRa71 netL71 1.3870121689568124e-09
Rbbr71 netL71 node_3 42465112.97562415
Cbr71 netL71 node_3 3.764777691495025e-22

* Branch 72
Rabr72 node_2 netRa72 1259848.6795585344
Lbr72 netRa72 netL72 9.491363739795341e-10
Rbbr72 netL72 node_3 -2964929.1603205707
Cbr72 netL72 node_3 2.541753674746829e-22

* Branch 73
Rabr73 node_2 netRa73 -6671241.4715043185
Lbr73 netRa73 netL73 1.5628832189652903e-09
Rbbr73 netL73 node_3 7426719.349668604
Cbr73 netL73 node_3 3.154119038907224e-23

* Branch 74
Rabr74 node_2 netRa74 -2945917.151941861
Lbr74 netRa74 netL74 1.868529320334269e-09
Rbbr74 netL74 node_3 4712389.976357865
Cbr74 netL74 node_3 1.3455868712686758e-22

* Branch 75
Rabr75 node_2 netRa75 370179.947652826
Lbr75 netRa75 netL75 1.6035123951251582e-09
Rbbr75 netL75 node_3 -13329212.309634347
Cbr75 netL75 node_3 3.2563073421556625e-22

* Branch 76
Rabr76 node_2 netRa76 -15899565.386411382
Lbr76 netRa76 netL76 3.6512251583784633e-09
Rbbr76 netL76 node_3 17341131.53303639
Cbr76 netL76 node_3 1.324127265371399e-23

* Branch 77
Rabr77 node_2 netRa77 48525.32214687523
Lbr77 netRa77 netL77 2.9632211626902294e-10
Rbbr77 netL77 node_3 -5094828.717766966
Cbr77 netL77 node_3 1.2020791073409054e-21

* Branch 78
Rabr78 node_2 netRa78 239354.0775816776
Lbr78 netRa78 netL78 7.384959580993699e-10
Rbbr78 netL78 node_3 -5065285.569338296
Cbr78 netL78 node_3 6.100387649760147e-22

* Branch 79
Rabr79 node_2 netRa79 1488500.6773866029
Lbr79 netRa79 netL79 1.1464340800770814e-09
Rbbr79 netL79 node_3 -3545354.939562271
Cbr79 netL79 node_3 2.173225314267794e-22

* Branch 80
Rabr80 node_2 netRa80 405075.95576283056
Lbr80 netRa80 netL80 8.994594838547455e-10
Rbbr80 netL80 node_3 -4738597.825639897
Cbr80 netL80 node_3 4.691354993467326e-22

* Branch 81
Rabr81 node_2 netRa81 215188.55104226686
Lbr81 netRa81 netL81 5.994277871934296e-10
Rbbr81 netL81 node_3 -4389880.933561378
Cbr81 netL81 node_3 6.355868682112192e-22

* Branch 82
Rabr82 node_2 netRa82 283452.1749116106
Lbr82 netRa82 netL82 6.505287789352078e-10
Rbbr82 netL82 node_3 -3930399.4411686906
Cbr82 netL82 node_3 5.847035889578901e-22

* Branch 83
Rabr83 node_2 netRa83 -449951.40269297577
Lbr83 netRa83 netL83 8.700292652787997e-10
Rbbr83 netL83 node_3 3830894.9315097504
Cbr83 netL83 node_3 5.041623745149257e-22

* Branch 84
Rabr84 node_2 netRa84 320584.8878844723
Lbr84 netRa84 netL84 9.917713130861766e-10
Rbbr84 netL84 node_3 -7312863.071199759
Cbr84 netL84 node_3 4.239108590336992e-22

* Branch 85
Rabr85 node_2 netRa85 -22334.80162035066
Lbr85 netRa85 netL85 4.331685158318726e-10
Rbbr85 netL85 node_3 21646687.610892016
Cbr85 netL85 node_3 8.8331815508036e-22

* Branch 86
Rabr86 node_2 netRa86 69516.89791744157
Lbr86 netRa86 netL86 3.9763947971399883e-10
Rbbr86 netL86 node_3 -6166743.886979708
Cbr86 netL86 node_3 9.316219378111414e-22

* Branch 87
Rabr87 node_2 netRa87 -3560247775.9348598
Lbr87 netRa87 netL87 -5.1581270263057256e-08
Rbbr87 netL87 node_3 3561497483.472891
Cbr87 netL87 node_3 -4.068028341604966e-27

* Branch 88
Rabr88 node_2 netRa88 -3005082.173292533
Lbr88 netRa88 netL88 1.5176929978550263e-09
Rbbr88 netL88 node_3 4508321.386826736
Cbr88 netL88 node_3 1.1197778712151817e-22

* Branch 89
Rabr89 node_2 netRa89 152288.8947676521
Lbr89 netRa89 netL89 4.033150249391943e-10
Rbbr89 netL89 node_3 -3071414.4456206444
Cbr89 netL89 node_3 8.641980132767998e-22

* Branch 90
Rabr90 node_2 netRa90 -516764.85000088724
Lbr90 netRa90 netL90 3.195926035983202e-10
Rbbr90 netL90 node_3 1128448.3638646305
Cbr90 netL90 node_3 5.477408593898701e-22

* Branch 91
Rabr91 node_2 netRa91 -540121.792335998
Lbr91 netRa91 netL91 4.165082824504602e-10
Rbbr91 netL91 node_3 1359651.6677353804
Cbr91 netL91 node_3 5.667436170315324e-22

* Branch 92
Rabr92 node_2 netRa92 -367787.66984728305
Lbr92 netRa92 netL92 3.295286986701846e-10
Rbbr92 netL92 node_3 1262573.4609911193
Cbr92 netL92 node_3 7.089553989350902e-22

* Branch 93
Rabr93 node_2 netRa93 -1106117.7368315784
Lbr93 netRa93 netL93 3.585140442972381e-10
Rbbr93 netL93 node_3 1473222.6749426974
Cbr93 netL93 node_3 2.1992305848456177e-22

* Branch 94
Rabr94 node_2 netRa94 -2173861.853407239
Lbr94 netRa94 netL94 5.914698576739931e-10
Rbbr94 netL94 node_3 2652025.9196142564
Cbr94 netL94 node_3 1.0255501256821694e-22

* Branch 95
Rabr95 node_2 netRa95 -441587.3502911783
Lbr95 netRa95 netL95 -2.0435551775854026e-10
Rbbr95 netL95 node_3 717552.273126488
Cbr95 netL95 node_3 -6.454045318401307e-22

* Branch 96
Rabr96 node_2 netRa96 -579400.6942759637
Lbr96 netRa96 netL96 2.607713678812588e-10
Rbbr96 netL96 node_3 957521.2803437469
Cbr96 netL96 node_3 4.69656058798303e-22

* Branch 97
Rabr97 node_2 netRa97 -414168.1181710686
Lbr97 netRa97 netL97 1.7497396387417552e-10
Rbbr97 netL97 node_3 656794.0026029242
Cbr97 netL97 node_3 6.42133354354678e-22

* Branch 98
Rabr98 node_2 netRa98 -1071045.1723736257
Lbr98 netRa98 netL98 4.227972950930836e-10
Rbbr98 netL98 node_3 1628806.5140100012
Cbr98 netL98 node_3 2.4191617311932623e-22

* Branch 99
Rabr99 node_2 netRa99 -618411.6284749418
Lbr99 netRa99 netL99 1.0569682980674141e-10
Rbbr99 netL99 node_3 680203.1904983808
Cbr99 netL99 node_3 2.502073943700559e-22

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 -30466410.944484357
Lbr0 netRa0 netL0 1.3233921526444974e-09
Rbbr0 netL0 node_4 30649438.04998695
Cbr0 netL0 node_4 1.4116576194651862e-24

* Branch 1
Rabr1 node_2 netRa1 -6511171.773340995
Lbr1 netRa1 netL1 5.805768596815027e-10
Rbbr1 netL1 node_4 6676554.392247318
Cbr1 netL1 node_4 1.3275245942666466e-23

* Branch 2
Rabr2 node_2 netRa2 -5391718.015721327
Lbr2 netRa2 netL2 4.795127892275372e-10
Rbbr2 netL2 node_4 5530178.630683724
Cbr2 netL2 node_4 1.6009368517699303e-23

* Branch 3
Rabr3 node_2 netRa3 -17864986.220585603
Lbr3 netRa3 netL3 -1.4191904338299395e-09
Rbbr3 netL3 node_4 18176971.728143215
Cbr3 netL3 node_4 -4.386478358173587e-24

* Branch 4
Rabr4 node_2 netRa4 -156226349.66951025
Lbr4 netRa4 netL4 -4.121978919210532e-09
Rbbr4 netL4 node_4 156523924.70740333
Cbr4 netL4 node_4 -1.687506313923439e-25

* Branch 5
Rabr5 node_2 netRa5 -13084562.399622006
Lbr5 netRa5 netL5 1.2218155498764265e-09
Rbbr5 netL5 node_4 13387973.190621665
Cbr5 netL5 node_4 6.957231344891622e-24

* Branch 6
Rabr6 node_2 netRa6 -1351057.2922020878
Lbr6 netRa6 netL6 1.1369292069655015e-09
Rbbr6 netL6 node_4 2343838.443730517
Cbr6 netL6 node_4 3.534603487668042e-22

* Branch 7
Rabr7 node_2 netRa7 -1271349.7256911655
Lbr7 netRa7 netL7 1.1676021308122394e-09
Rbbr7 netL7 node_4 2297295.8732124427
Cbr7 netL7 node_4 3.9302339591816344e-22

* Branch 8
Rabr8 node_2 netRa8 -1189985.9389716536
Lbr8 netRa8 netL8 1.1970310871080097e-09
Rbbr8 netL8 node_4 2248131.641702523
Cbr8 netL8 node_4 4.393341751659991e-22

* Branch 9
Rabr9 node_2 netRa9 -1429893.3945939206
Lbr9 netRa9 netL9 1.1041436798674434e-09
Rbbr9 netL9 node_4 2387836.1326442114
Cbr9 netL9 node_4 3.1892408851894416e-22

* Branch 10
Rabr10 node_2 netRa10 -1108198.5364142624
Lbr10 netRa10 netL10 1.2254427161802515e-09
Rbbr10 netL10 node_4 2197424.702042168
Cbr10 netL10 node_4 4.934145217944108e-22

* Branch 11
Rabr11 node_2 netRa11 1589056.5773706196
Lbr11 netRa11 netL11 4.762088206613125e-10
Rbbr11 netL11 node_4 -2000933.7151926567
Cbr11 netL11 node_4 1.505731342291202e-22

* Branch 12
Rabr12 node_2 netRa12 -2373273.7923810505
Lbr12 netRa12 netL12 6.830746815494905e-10
Rbbr12 netL12 node_4 2830691.3267290257
Cbr12 netL12 node_4 1.0116174510864025e-22

* Branch 13
Rabr13 node_2 netRa13 -470196.1401692508
Lbr13 netRa13 netL13 2.2482345639164524e-10
Rbbr13 netL13 node_4 791480.2042989157
Cbr13 netL13 node_4 5.991417653093843e-22

* Branch 14
Rabr14 node_2 netRa14 -1584078.2574581997
Lbr14 netRa14 netL14 1.0362402907600725e-09
Rbbr14 netL14 node_4 2469184.4811572144
Cbr14 netL14 node_4 2.6204387387203576e-22

* Branch 15
Rabr15 node_2 netRa15 -1506002.3655001791
Lbr15 netRa15 netL15 1.0705716002739842e-09
Rbbr15 netL15 node_4 2428676.6072916556
Cbr15 netL15 node_4 2.8924862347234793e-22

* Branch 16
Rabr16 node_2 netRa16 -944852.3056571768
Lbr16 netRa16 netL16 1.2788277442354332e-09
Rbbr16 netL16 node_4 2092558.1304546185
Cbr16 netL16 node_4 6.329397758678595e-22

* Branch 17
Rabr17 node_2 netRa17 -546423.2064047065
Lbr17 netRa17 netL17 -1.1121024303206796e-10
Rbbr17 netL17 node_4 624235.7212685837
Cbr17 netL17 node_4 -3.271124483818616e-22

* Branch 18
Rabr18 node_2 netRa18 -1660030.2507433067
Lbr18 netRa18 netL18 1.0002955753389658e-09
Rbbr18 netL18 node_4 2505463.3299351344
Cbr18 netL18 node_4 2.3818891041904134e-22

* Branch 19
Rabr19 node_2 netRa19 -1025188.1481488342
Lbr19 netRa19 netL19 1.2526284152563006e-09
Rbbr19 netL19 node_4 2146149.5419245185
Cbr19 netL19 node_4 5.5840328844372755e-22

* Branch 20
Rabr20 node_2 netRa20 -2787547.3191727693
Lbr20 netRa20 netL20 6.735535088150372e-10
Rbbr20 netL20 node_4 3186360.575141405
Cbr20 netL20 node_4 7.554393958306905e-23

* Branch 21
Rabr21 node_2 netRa21 -2128781.3805550653
Lbr21 netRa21 netL21 7.2267388504948e-10
Rbbr21 netL21 node_4 2660398.668365024
Cbr21 netL21 node_4 1.2692591108459656e-22

* Branch 22
Rabr22 node_2 netRa22 -862916.5852273309
Lbr22 netRa22 netL22 1.303733751618403e-09
Rbbr22 netL22 node_4 2039927.0693804245
Cbr22 netL22 node_4 7.244614121590516e-22

* Branch 23
Rabr23 node_2 netRa23 -1908003.976523883
Lbr23 netRa23 netL23 8.972707922479019e-10
Rbbr23 netL23 node_4 2633492.799392165
Cbr23 netL23 node_4 1.773919614028944e-22

* Branch 24
Rabr24 node_2 netRa24 -1701855.9698251325
Lbr24 netRa24 netL24 9.576816858531935e-10
Rbbr24 netL24 node_4 2513022.550570571
Cbr24 netL24 node_4 2.222144519231954e-22

* Branch 25
Rabr25 node_2 netRa25 -703924.4286959218
Lbr25 netRa25 netL25 1.3527835176683052e-09
Rbbr25 netL25 node_4 1929861.3805630258
Cbr25 netL25 node_4 9.70884514219718e-22

* Branch 26
Rabr26 node_2 netRa26 -783020.9924179488
Lbr26 netRa26 netL26 1.3290826505676268e-09
Rbbr26 netL26 node_4 1986778.856728496
Cbr26 netL26 node_4 8.356126921223262e-22

* Branch 27
Rabr27 node_2 netRa27 -1791955.1741148976
Lbr27 netRa27 netL27 9.210820441525173e-10
Rbbr27 netL27 node_4 2551355.162490652
Cbr27 netL27 node_4 2.0021884508376565e-22

* Branch 28
Rabr28 node_2 netRa28 -1993532.8992951289
Lbr28 netRa28 netL28 7.601354145362605e-10
Rbbr28 netL28 node_4 2582837.898780145
Cbr28 netL28 node_4 1.469942320093176e-22

* Branch 29
Rabr29 node_2 netRa29 -1899709.0671039992
Lbr29 netRa29 netL29 8.29974129241606e-10
Rbbr29 netL29 node_4 2572348.2166063045
Cbr29 netL29 node_4 1.6903937606937991e-22

* Branch 30
Rabr30 node_2 netRa30 -1973819.7180749683
Lbr30 netRa30 netL30 7.379028559981042e-10
Rbbr30 netL30 node_4 2547344.5230855644
Cbr30 netL30 node_4 1.4631676804877715e-22

* Branch 31
Rabr31 node_2 netRa31 242056.493100406
Lbr31 netRa31 netL31 2.7307823008814915e-10
Rbbr31 netL31 node_4 -1298266.536412998
Cbr31 netL31 node_4 8.69791173363187e-22

* Branch 32
Rabr32 node_2 netRa32 5662902.025742724
Lbr32 netRa32 netL32 -8.431236287015741e-09
Rbbr32 netL32 node_4 -40641975.15095814
Cbr32 netL32 node_4 -3.661360977834618e-23

* Branch 33
Rabr33 node_2 netRa33 -345235610.1725302
Lbr33 netRa33 netL33 -2.6911198320138414e-08
Rbbr33 netL33 node_4 350958486.8499893
Cbr33 netL33 node_4 -2.221070615813687e-25

* Branch 34
Rabr34 node_2 netRa34 -4059939.1591132586
Lbr34 netRa34 netL34 1.1310677714092128e-08
Rbbr34 netL34 node_4 21978949.71311235
Cbr34 netL34 node_4 1.267489720273922e-22

* Branch 35
Rabr35 node_2 netRa35 -3834331.283400041
Lbr35 netRa35 netL35 1.169730518418951e-08
Rbbr35 netL35 node_4 23171986.048686434
Cbr35 netL35 node_4 1.3164806921081826e-22

* Branch 36
Rabr36 node_2 netRa36 -4938527.1423304705
Lbr36 netRa36 netL36 1.105685781261209e-08
Rbbr36 netL36 node_4 23325307.635701746
Cbr36 netL36 node_4 9.598320666587993e-23

* Branch 37
Rabr37 node_2 netRa37 -4307107.482164856
Lbr37 netRa37 netL37 1.1566468050361697e-08
Rbbr37 netL37 node_4 22821525.92740827
Cbr37 netL37 node_4 1.17667498507762e-22

* Branch 38
Rabr38 node_2 netRa38 -3777863.6116899042
Lbr38 netRa38 netL38 1.1711567880996978e-08
Rbbr38 netL38 node_4 22504583.862642866
Cbr38 netL38 node_4 1.3774755497963012e-22

* Branch 39
Rabr39 node_2 netRa39 -3292530.1265561865
Lbr39 netRa39 netL39 1.1531530201769491e-08
Rbbr39 netL39 node_4 23095681.672528
Cbr39 netL39 node_4 1.5164064718413523e-22

* Branch 40
Rabr40 node_2 netRa40 -3388301.559755474
Lbr40 netRa40 netL40 1.1979734506082254e-08
Rbbr40 netL40 node_4 23105281.007333495
Cbr40 netL40 node_4 1.5301873907062564e-22

* Branch 41
Rabr41 node_2 netRa41 -3209903.013462223
Lbr41 netRa41 netL41 1.1978239850358245e-08
Rbbr41 netL41 node_4 22936834.39158067
Cbr41 netL41 node_4 1.626896177084073e-22

* Branch 42
Rabr42 node_2 netRa42 -3017731.171792966
Lbr42 netRa42 netL42 1.1997226241293012e-08
Rbbr42 netL42 node_4 22945075.850792687
Cbr42 netL42 node_4 1.7326237624316085e-22

* Branch 43
Rabr43 node_2 netRa43 -4026362.8683694527
Lbr43 netRa43 netL43 1.1108300957819916e-08
Rbbr43 netL43 node_4 23153615.402816553
Cbr43 netL43 node_4 1.1915487532832945e-22

* Branch 44
Rabr44 node_2 netRa44 -2851214.5838467865
Lbr44 netRa44 netL44 1.2051289516901404e-08
Rbbr44 netL44 node_4 22967001.760464262
Cbr44 netL44 node_4 1.8403208632233356e-22

* Branch 45
Rabr45 node_2 netRa45 -4432624.81615963
Lbr45 netRa45 netL45 1.0805403669999168e-08
Rbbr45 netL45 node_4 23190574.94941176
Cbr45 netL45 node_4 1.0511566064995193e-22

* Branch 46
Rabr46 node_2 netRa46 -4170764.282920321
Lbr46 netRa46 netL46 1.1100511849041564e-08
Rbbr46 netL46 node_4 23457721.379769597
Cbr46 netL46 node_4 1.1345945480051689e-22

* Branch 47
Rabr47 node_2 netRa47 -4049767.256687188
Lbr47 netRa47 netL47 1.0779886869830452e-08
Rbbr47 netL47 node_4 23623908.71523079
Cbr47 netL47 node_4 1.1267614542811483e-22

* Branch 48
Rabr48 node_2 netRa48 -23870222.301651556
Lbr48 netRa48 netL48 1.73788761845442e-08
Rbbr48 netL48 node_4 43855926.35397312
Cbr48 netL48 node_4 1.6601076235329233e-23

* Branch 49
Rabr49 node_2 netRa49 -5281355.883439379
Lbr49 netRa49 netL49 -1.0420299009229634e-08
Rbbr49 netL49 node_4 22520972.72823902
Cbr49 netL49 node_4 -8.760965827018598e-23

* Branch 50
Rabr50 node_2 netRa50 -4110222.216370223
Lbr50 netRa50 netL50 -9.94483639033626e-09
Rbbr50 netL50 node_4 25085618.788870078
Cbr50 netL50 node_4 -9.64523808863654e-23

* Branch 51
Rabr51 node_2 netRa51 -6255134.81821525
Lbr51 netRa51 netL51 -1.0423022973510012e-08
Rbbr51 netL51 node_4 21983160.839259498
Cbr51 netL51 node_4 -7.580028669861968e-23

* Branch 52
Rabr52 node_2 netRa52 -3752235.1098200455
Lbr52 netRa52 netL52 -1.0161700291461953e-08
Rbbr52 netL52 node_4 25932031.530199908
Cbr52 netL52 node_4 -1.0443514112410551e-22

* Branch 53
Rabr53 node_2 netRa53 -5607205.870330318
Lbr53 netRa53 netL53 -1.0116045610255307e-08
Rbbr53 netL53 node_4 22763954.24458526
Cbr53 netL53 node_4 -7.925400527683633e-23

* Branch 54
Rabr54 node_2 netRa54 -4347882.911227475
Lbr54 netRa54 netL54 -9.442537513501884e-09
Rbbr54 netL54 node_4 24346455.79072345
Cbr54 netL54 node_4 -8.920339090505714e-23

* Branch 55
Rabr55 node_2 netRa55 -5093734.449642687
Lbr55 netRa55 netL55 -9.567735819046408e-09
Rbbr55 netL55 node_4 23262758.682862792
Cbr55 netL55 node_4 -8.074537193570553e-23

* Branch 56
Rabr56 node_2 netRa56 -10148965.20268624
Lbr56 netRa56 netL56 -1.2793684136834696e-08
Rbbr56 netL56 node_4 22632358.121565405
Cbr56 netL56 node_4 -5.569914266081724e-23

* Branch 57
Rabr57 node_2 netRa57 -4639811.623712021
Lbr57 netRa57 netL57 -9.286705256765514e-09
Rbbr57 netL57 node_4 24108988.879626963
Cbr57 netL57 node_4 -8.302136759282595e-23

* Branch 58
Rabr58 node_2 netRa58 -6016174.300974302
Lbr58 netRa58 netL58 -9.526050050781468e-09
Rbbr58 netL58 node_4 22374351.175313868
Cbr58 netL58 node_4 -7.076993041750089e-23

* Branch 59
Rabr59 node_2 netRa59 -6330637.147826051
Lbr59 netRa59 netL59 -9.573301853253383e-09
Rbbr59 netL59 node_4 22576930.290781427
Cbr59 netL59 node_4 -6.698186571353794e-23

* Branch 60
Rabr60 node_2 netRa60 -5759680.415064658
Lbr60 netRa60 netL60 -9.08277884785023e-09
Rbbr60 netL60 node_4 22382963.589835227
Cbr60 netL60 node_4 -7.045499963319096e-23

* Branch 61
Rabr61 node_2 netRa61 -6930223.813892478
Lbr61 netRa61 netL61 -9.446934866407116e-09
Rbbr61 netL61 node_4 22378108.818637606
Cbr61 netL61 node_4 -6.091576455156889e-23

* Branch 62
Rabr62 node_2 netRa62 -8674123.72757154
Lbr62 netRa62 netL62 -9.762356136062566e-09
Rbbr62 netL62 node_4 22289864.284828704
Cbr62 netL62 node_4 -5.0493128268558507e-23

* Branch 63
Rabr63 node_2 netRa63 -3621154.388827595
Lbr63 netRa63 netL63 -8.148990138026943e-09
Rbbr63 netL63 node_4 27086936.323101778
Cbr63 netL63 node_4 -8.308571202636995e-23

* Branch 64
Rabr64 node_2 netRa64 -4365128.834156615
Lbr64 netRa64 netL64 -8.205349572836066e-09
Rbbr64 netL64 node_4 24733260.72952908
Cbr64 netL64 node_4 -7.600649189398015e-23

* Branch 65
Rabr65 node_2 netRa65 -3469336.065414834
Lbr65 netRa65 netL65 -7.925322915697135e-09
Rbbr65 netL65 node_4 28130921.29492042
Cbr65 netL65 node_4 -8.121410625034458e-23

* Branch 66
Rabr66 node_2 netRa66 27093999.906352647
Lbr66 netRa66 netL66 -2.7726047135167362e-08
Rbbr66 netL66 node_4 -77182711.6819713
Cbr66 netL66 node_4 -1.3257770261730737e-23

* Branch 67
Rabr67 node_2 netRa67 -119942518.89790425
Lbr67 netRa67 netL67 -4.365447691066696e-08
Rbbr67 netL67 node_4 144328507.04280692
Cbr67 netL67 node_4 -2.521815816456246e-24

* Branch 68
Rabr68 node_2 netRa68 908497.8075783608
Lbr68 netRa68 netL68 -7.090500079924117e-09
Rbbr68 netL68 node_4 -78581687.48145443
Cbr68 netL68 node_4 -9.927021304269854e-23

* Branch 69
Rabr69 node_2 netRa69 -3141415.1699290606
Lbr69 netRa69 netL69 -2.6011417555667554e-08
Rbbr69 netL69 node_4 393921194.5282942
Cbr69 netL69 node_4 -2.103103096764716e-23

* Branch 70
Rabr70 node_2 netRa70 -27142241.938670967
Lbr70 netRa70 netL70 -1.0963839940216373e-08
Rbbr70 netL70 node_4 36509377.81195431
Cbr70 netL70 node_4 -1.106433256876405e-23

* Branch 71
Rabr71 node_2 netRa71 -19490824.197582483
Lbr71 netRa71 netL71 -7.944329191647346e-09
Rbbr71 netL71 node_4 27391761.99602221
Cbr71 netL71 node_4 -1.4880609948735563e-23

* Branch 72
Rabr72 node_2 netRa72 -63952726.83583501
Lbr72 netRa72 netL72 -2.1786154428279893e-08
Rbbr72 netL72 node_4 78138013.29686841
Cbr72 netL72 node_4 -4.35984435657539e-24

* Branch 73
Rabr73 node_2 netRa73 18795123.6793986
Lbr73 netRa73 netL73 -7.993094477929115e-09
Rbbr73 netL73 node_4 -25808476.21176373
Cbr73 netL73 node_4 -1.647749593782313e-23

* Branch 74
Rabr74 node_2 netRa74 4138641.7359855524
Lbr74 netRa74 netL74 -7.536844164170313e-09
Rbbr74 netL74 node_4 -23998304.881221212
Cbr74 netL74 node_4 -7.587197907773484e-23

* Branch 75
Rabr75 node_2 netRa75 -37970578.65698954
Lbr75 netRa75 netL75 -1.427088398307907e-08
Rbbr75 netL75 node_4 49882013.597473614
Cbr75 netL75 node_4 -7.534852962884358e-24

* Branch 76
Rabr76 node_2 netRa76 -6978897.802804712
Lbr76 netRa76 netL76 -1.7750989404647436e-08
Rbbr76 netL76 node_4 80370179.94536231
Cbr76 netL76 node_4 -3.165536074669481e-23

* Branch 77
Rabr77 node_2 netRa77 60540199.80020191
Lbr77 netRa77 netL77 -1.7670440766526757e-08
Rbbr77 netL77 node_4 -68228766.32631676
Cbr77 netL77 node_4 -4.277826084457246e-24

* Branch 78
Rabr78 node_2 netRa78 -10907750.980073584
Lbr78 netRa78 netL78 -7.167243792249469e-09
Rbbr78 netL78 node_4 21877060.781785063
Cbr78 netL78 node_4 -3.0037035635564667e-23

* Branch 79
Rabr79 node_2 netRa79 -11032256.250610644
Lbr79 netRa79 netL79 -6.990090512165609e-09
Rbbr79 netL79 node_4 21592378.154290423
Cbr79 netL79 node_4 -2.9345911265158235e-23

* Branch 80
Rabr80 node_2 netRa80 1664652.9485478895
Lbr80 netRa80 netL80 -5.1364449341462556e-09
Rbbr80 netL80 node_4 -33540255.87956872
Cbr80 netL80 node_4 -9.196178766521917e-23

* Branch 81
Rabr81 node_2 netRa81 -1414250.8295168334
Lbr81 netRa81 netL81 -3.2486619411196917e-09
Rbbr81 netL81 node_4 20905547.188229673
Cbr81 netL81 node_4 -1.0991105858429835e-22

* Branch 82
Rabr82 node_2 netRa82 -1513960.2246610655
Lbr82 netRa82 netL82 -8.306781536829013e-09
Rbbr82 netL82 node_4 86440352.73424678
Cbr82 netL82 node_4 -6.35191056207588e-23

* Branch 83
Rabr83 node_2 netRa83 -3342015.3573602745
Lbr83 netRa83 netL83 -3.5323283209311873e-09
Rbbr83 netL83 node_4 13309594.699455485
Cbr83 netL83 node_4 -7.942316310563631e-23

* Branch 84
Rabr84 node_2 netRa84 -3249890.598038159
Lbr84 netRa84 netL84 -5.4376503782212095e-09
Rbbr84 netL84 node_4 23949456.364382014
Cbr84 netL84 node_4 -6.987864699558951e-23

* Branch 85
Rabr85 node_2 netRa85 -2160004.49282962
Lbr85 netRa85 netL85 -4.04291885027409e-09
Rbbr85 netL85 node_4 21055518.05451795
Cbr85 netL85 node_4 -8.891719633893348e-23

* Branch 86
Rabr86 node_2 netRa86 -542959.3792949496
Lbr86 netRa86 netL86 -4.944592087766589e-09
Rbbr86 netL86 node_4 98272826.98484115
Cbr86 netL86 node_4 -9.278484576235964e-23

* Branch 87
Rabr87 node_2 netRa87 -535882.5214213397
Lbr87 netRa87 netL87 -3.426196600533215e-09
Rbbr87 netL87 node_4 56523422.33412436
Cbr87 netL87 node_4 -1.132189479521447e-22

* Branch 88
Rabr88 node_2 netRa88 42940329.062849514
Lbr88 netRa88 netL88 -1.3969919076170369e-08
Rbbr88 netL88 node_4 -50535985.91808368
Cbr88 netL88 node_4 -6.437341034234013e-24

* Branch 89
Rabr89 node_2 netRa89 4700908.923274555
Lbr89 netRa89 netL89 -6.672945997823232e-09
Rbbr89 netL89 node_4 -23275250.37407239
Cbr89 netL89 node_4 -6.097153756371585e-23

* Branch 90
Rabr90 node_2 netRa90 112217614.63351427
Lbr90 netRa90 netL90 -1.9452977601141283e-08
Rbbr90 netL90 node_4 -118011701.88482256
Cbr90 netL90 node_4 -1.4688762349237185e-24

* Branch 91
Rabr91 node_2 netRa91 1250396.371152221
Lbr91 netRa91 netL91 6.199231271517284e-10
Rbbr91 netL91 node_4 -2146260.0294714044
Cbr91 netL91 node_4 2.310329024512571e-22

* Branch 92
Rabr92 node_2 netRa92 1070599.0132815596
Lbr92 netRa92 netL92 -1.0508610705170485e-09
Rbbr92 netL92 node_4 -4328689.931389392
Cbr92 netL92 node_4 -2.2667348060946094e-22

* Branch 93
Rabr93 node_2 netRa93 970971.2178922022
Lbr93 netRa93 netL93 -1.111369067280754e-09
Rbbr93 netL93 node_4 -4907844.3184041735
Cbr93 netL93 node_4 -2.331095729424867e-22

* Branch 94
Rabr94 node_2 netRa94 23080.61359240005
Lbr94 netRa94 netL94 -8.965106028659421e-10
Rbbr94 netL94 node_4 -110395466.25206386
Cbr94 netL94 node_4 -3.459329844158729e-22

* Branch 95
Rabr95 node_2 netRa95 1726547.9452101972
Lbr95 netRa95 netL95 -1.1565257064762183e-09
Rbbr95 netL95 node_4 -4075789.0950855725
Cbr95 netL95 node_4 -1.6428213598644102e-22

* Branch 96
Rabr96 node_2 netRa96 568440.9851581651
Lbr96 netRa96 netL96 -8.668499598946665e-10
Rbbr96 netL96 node_4 -4911264.780967987
Cbr96 netL96 node_4 -3.1017636666473997e-22

* Branch 97
Rabr97 node_2 netRa97 3625214.9102907456
Lbr97 netRa97 netL97 -1.355442354793304e-09
Rbbr97 netL97 node_4 -5131088.39568002
Cbr97 netL97 node_4 -7.284765212771357e-23

* Branch 98
Rabr98 node_2 netRa98 2751506.0350268357
Lbr98 netRa98 netL98 -1.1721565226928377e-09
Rbbr98 netL98 node_4 -4426154.138051597
Cbr98 netL98 node_4 -9.621320631033389e-23

* Branch 99
Rabr99 node_2 netRa99 276769.85381548206
Lbr99 netRa99 netL99 1.2088011929045868e-10
Rbbr99 netL99 node_4 -462195.02764673607
Cbr99 netL99 node_4 9.522630092911428e-22

.ends


* Y'33
.subckt yp33 node_3 0
* Branch 0
Rabr0 node_3 netRa0 158578.78844908168
Lbr0 netRa0 netL0 1.1604213258789739e-11
Rbbr0 netL0 0 -161740.87857058368
Cbr0 netL0 0 4.596435062986448e-22

* Branch 1
Rabr1 node_3 netRa1 2575931.6667255647
Lbr1 netRa1 netL1 -4.619371586188315e-11
Rbbr1 netL1 0 -2578953.6411949587
Cbr1 netL1 0 -6.928893321394493e-24

* Branch 2
Rabr2 node_3 netRa2 251197.67480552706
Lbr2 netRa2 netL2 -1.4577602306424668e-11
Rbbr2 netL2 0 -254256.1636855531
Cbr2 netL2 0 -2.25719802787388e-22

* Branch 3
Rabr3 node_3 netRa3 23058.201735704417
Lbr3 netRa3 netL3 -4.838961060634758e-12
Rbbr3 netL3 0 -26615.524790605046
Cbr3 netL3 0 -7.60124660387465e-21

* Branch 4
Rabr4 node_3 netRa4 1559.3891658665386
Lbr4 netRa4 netL4 -2.400649180524659e-12
Rbbr4 netL4 0 -12350.603224570945
Cbr4 netL4 0 -1.012629166137997e-19

* Branch 5
Rabr5 node_3 netRa5 -2786010.4862513356
Lbr5 netRa5 netL5 4.540169537165732e-11
Rbbr5 netL5 0 2788625.788085845
Cbr5 netL5 0 5.8331637772889916e-24

* Branch 6
Rabr6 node_3 netRa6 95660.58587684298
Lbr6 netRa6 netL6 8.915371055084392e-12
Rbbr6 netL6 0 -98568.38119679174
Cbr6 netL6 0 9.524522823835222e-22

* Branch 7
Rabr7 node_3 netRa7 -95314.37112061627
Lbr7 netRa7 netL7 3.0045505027846537e-11
Rbbr7 netL7 0 102383.58696141449
Cbr7 netL7 0 3.008029339198452e-21

* Branch 8
Rabr8 node_3 netRa8 -279962.8219839038
Lbr8 netRa8 netL8 5.025555876333437e-11
Rbbr8 netL8 0 286802.8336156266
Cbr8 netL8 0 6.195084218979049e-22

* Branch 9
Rabr9 node_3 netRa9 5872.7701190928965
Lbr9 netRa9 netL9 -1.877670177979358e-12
Rbbr9 netL9 0 -7854.4067580579
Cbr9 netL9 0 -4.005961349254425e-20

* Branch 10
Rabr10 node_3 netRa10 -195.0193544342493
Lbr10 netRa10 netL10 7.813791413436548e-13
Rbbr10 netL10 0 8883.394521559872
Cbr10 netL10 0 3.7580694419998734e-19

* Branch 11
Rabr11 node_3 netRa11 -597192.102904898
Lbr11 netRa11 netL11 7.273053545611974e-11
Rbbr11 netL11 0 603945.6386405791
Cbr11 netL11 0 2.0066939251271628e-22

* Branch 12
Rabr12 node_3 netRa12 -187796.37377273006
Lbr12 netRa12 netL12 4.239882633319168e-11
Rbbr12 netL12 0 195064.6902503379
Cbr12 netL12 0 1.1492228207440448e-21

* Branch 13
Rabr13 node_3 netRa13 8728.594901200697
Lbr13 netRa13 netL13 3.2088772796192782e-12
Rbbr13 netL13 0 -12573.168856752422
Cbr13 netL13 0 2.9560641157570696e-20

* Branch 14
Rabr14 node_3 netRa14 -56131.49417076134
Lbr14 netRa14 netL14 2.496845202130014e-11
Rbbr14 netL14 0 64517.60982915474
Cbr14 netL14 0 6.813583429344935e-21

* Branch 15
Rabr15 node_3 netRa15 -2079.140840460049
Lbr15 netRa15 netL15 2.0851159773827588e-12
Rbbr15 netL15 0 8596.3734997697
Cbr15 netL15 0 1.1389292492170705e-19

* Branch 16
Rabr16 node_3 netRa16 5891.197142394252
Lbr16 netRa16 netL16 3.972691453004193e-12
Rbbr16 netL16 0 -12328.66649748826
Cbr16 netL16 0 5.560251048718977e-20

* Branch 17
Rabr17 node_3 netRa17 -91217.29397133666
Lbr17 netRa17 netL17 -2.1337140197779244e-11
Rbbr17 netL17 0 105161.6191982915
Cbr17 netL17 0 -2.2359288180040513e-21

* Branch 18
Rabr18 node_3 netRa18 -3126.272214274657
Lbr18 netRa18 netL18 -5.088068437117104e-12
Rbbr18 netL18 0 26265.253230318376
Cbr18 netL18 0 -6.412791758052675e-20

* Branch 19
Rabr19 node_3 netRa19 1993.8813941335436
Lbr19 netRa19 netL19 3.711374456444805e-12
Rbbr19 netL19 0 -16355.376565425351
Cbr19 netL19 0 1.1836021531269983e-19

* Branch 20
Rabr20 node_3 netRa20 7468757.997790704
Lbr20 netRa20 netL20 -1.6737842937780773e-10
Rbbr20 netL20 0 -7476406.904979644
Cbr20 netL20 0 -2.996125399616337e-24

* Branch 21
Rabr21 node_3 netRa21 732320.6153335628
Lbr21 netRa21 netL21 8.163617857124347e-11
Rbbr21 netL21 0 -745997.5650203739
Cbr21 netL21 0 1.4977175354381644e-22

* Branch 22
Rabr22 node_3 netRa22 3505.142755131921
Lbr22 netRa22 netL22 3.2992315191345208e-12
Rbbr22 netL22 0 -11537.26055783935
Cbr22 netL22 0 8.316114654062142e-20

* Branch 23
Rabr23 node_3 netRa23 -16075.36398957615
Lbr23 netRa23 netL23 7.320369699611945e-12
Rbbr23 netL23 0 25637.223481815377
Cbr23 netL23 0 1.7601280562963322e-20

* Branch 24
Rabr24 node_3 netRa24 -39781023.442396455
Lbr24 netRa24 netL24 3.7421130626353805e-10
Rbbr24 netL24 0 39791026.02679252
Cbr24 netL24 0 2.3636037829765255e-25

* Branch 25
Rabr25 node_3 netRa25 150626.5574586967
Lbr25 netRa25 netL25 7.35111519404987e-11
Rbbr25 netL25 0 -166193.601109506
Cbr25 netL25 0 2.9652279808740317e-21

* Branch 26
Rabr26 node_3 netRa26 49.23593918916588
Lbr26 netRa26 netL26 3.2736620097310137e-12
Rbbr26 netL26 0 1619419.8543332478
Cbr26 netL26 0 1.3251944519719618e-19

* Branch 27
Rabr27 node_3 netRa27 -3283.593380459264
Lbr27 netRa27 netL27 -6.457546067889811e-12
Rbbr27 netL27 0 13180.059162510795
Cbr27 netL27 0 -1.5517160165854286e-19

* Branch 28
Rabr28 node_3 netRa28 -22467.609429257922
Lbr28 netRa28 netL28 7.53072555304299e-12
Rbbr28 netL28 0 29901.2898736761
Cbr28 netL28 0 1.1137063080783075e-20

* Branch 29
Rabr29 node_3 netRa29 -2808.573831951331
Lbr29 netRa29 netL29 3.63887696501685e-12
Rbbr29 netL29 0 16685.651007657572
Cbr29 netL29 0 7.584420941137337e-20

* Branch 30
Rabr30 node_3 netRa30 3287.7799579285074
Lbr30 netRa30 netL30 5.487878796188966e-12
Rbbr30 netL30 0 -28277.60350546281
Cbr30 netL30 0 6.089227728885919e-20

* Branch 31
Rabr31 node_3 netRa31 -851.153423074731
Lbr31 netRa31 netL31 4.510110332083225e-12
Rbbr31 netL31 0 43333.902834106586
Cbr31 netL31 0 1.1148363860679828e-19

* Branch 32
Rabr32 node_3 netRa32 1583.5839589080974
Lbr32 netRa32 netL32 5.73695247303987e-12
Rbbr32 netL32 0 -34261.58213357986
Cbr32 netL32 0 1.1315071496074936e-19

* Branch 33
Rabr33 node_3 netRa33 2021.4295469233564
Lbr33 netRa33 netL33 5.891427760479398e-12
Rbbr33 netL33 0 -50212.60984761112
Cbr33 netL33 0 6.125723465569233e-20

* Branch 34
Rabr34 node_3 netRa34 26016.71666965969
Lbr34 netRa34 netL34 1.2404275353681495e-11
Rbbr34 netL34 0 -35600.86271109856
Cbr34 netL34 0 1.3507969550319113e-20

* Branch 35
Rabr35 node_3 netRa35 5499.212049654715
Lbr35 netRa35 netL35 5.5555288179064605e-12
Rbbr35 netL35 0 -15785.661927801111
Cbr35 netL35 0 6.516672268183971e-20

* Branch 36
Rabr36 node_3 netRa36 -11690.448645797895
Lbr36 netRa36 netL36 8.575360201789855e-12
Rbbr36 netL36 0 23533.96624281871
Cbr36 netL36 0 3.07754796923508e-20

* Branch 37
Rabr37 node_3 netRa37 19281.478861475352
Lbr37 netRa37 netL37 -8.882609093652382e-12
Rbbr37 netL37 0 -29065.70560959121
Cbr37 netL37 0 -1.5724113353845405e-20

* Branch 38
Rabr38 node_3 netRa38 -2892.030794349789
Lbr38 netRa38 netL38 7.564116677084057e-12
Rbbr38 netL38 0 32647.47304986946
Cbr38 netL38 0 7.664817726815059e-20

* Branch 39
Rabr39 node_3 netRa39 -140975.9473962051
Lbr39 netRa39 netL39 4.693605742740925e-11
Rbbr39 netL39 0 164830.74191636412
Cbr39 netL39 0 2.0085186280831735e-21

* Branch 40
Rabr40 node_3 netRa40 -29033.783452278753
Lbr40 netRa40 netL40 1.730983829303055e-11
Rbbr40 netL40 0 43306.55010275982
Cbr40 netL40 0 1.362944296754028e-20

* Branch 41
Rabr41 node_3 netRa41 -2260.078653895273
Lbr41 netRa41 netL41 4.042406530806126e-12
Rbbr41 netL41 0 23827.20307521676
Cbr41 netL41 0 7.286893947671248e-20

* Branch 42
Rabr42 node_3 netRa42 -5621.123993076366
Lbr42 netRa42 netL42 4.841255549662144e-12
Rbbr42 netL42 0 18520.77235634791
Cbr42 netL42 0 4.5845920531238436e-20

* Branch 43
Rabr43 node_3 netRa43 3898.583134665484
Lbr43 netRa43 netL43 5.738898172922286e-12
Rbbr43 netL43 0 -18665.41388988826
Cbr43 netL43 0 8.079995519538533e-20

* Branch 44
Rabr44 node_3 netRa44 -2043.7140358139063
Lbr44 netRa44 netL44 7.086506153001264e-12
Rbbr44 netL44 0 35499.70574478686
Cbr44 netL44 0 9.290718839456844e-20

* Branch 45
Rabr45 node_3 netRa45 -164992.81178170728
Lbr45 netRa45 netL45 4.3354097869840725e-11
Rbbr45 netL45 0 186095.99278160755
Cbr45 netL45 0 1.4065535248154093e-21

* Branch 46
Rabr46 node_3 netRa46 5329.887365218566
Lbr46 netRa46 netL46 8.82245322691585e-12
Rbbr46 netL46 0 -22364.771671151495
Cbr46 netL46 0 7.582930541812145e-20

* Branch 47
Rabr47 node_3 netRa47 74726.70901850876
Lbr47 netRa47 netL47 1.5357341924800797e-11
Rbbr47 netL47 0 -81377.49269964412
Cbr47 netL47 0 2.5327341281499588e-21

* Branch 48
Rabr48 node_3 netRa48 -20399.096849076603
Lbr48 netRa48 netL48 1.0185549964888438e-11
Rbbr48 netL48 0 32969.533645351825
Cbr48 netL48 0 1.5040996306537425e-20

* Branch 49
Rabr49 node_3 netRa49 -16531.63463194507
Lbr49 netRa49 netL49 1.4374816885532614e-11
Rbbr49 netL49 0 37136.42481994655
Cbr49 netL49 0 2.314205772536723e-20

* Branch 50
Rabr50 node_3 netRa50 3917.9264553793596
Lbr50 netRa50 netL50 5.7146395470021e-12
Rbbr50 netL50 0 -15232.201798366434
Cbr50 netL50 0 9.764979351981128e-20

* Branch 51
Rabr51 node_3 netRa51 -351773.56109460164
Lbr51 netRa51 netL51 -6.987195397632547e-11
Rbbr51 netL51 0 382682.63468502613
Cbr51 netL51 0 -5.203938635236151e-22

* Branch 52
Rabr52 node_3 netRa52 25973.962790590536
Lbr52 netRa52 netL52 3.711872312770738e-11
Rbbr52 netL52 0 -82450.65786981826
Cbr52 netL52 0 1.7641403742481808e-20

* Branch 53
Rabr53 node_3 netRa53 804051.5764701905
Lbr53 netRa53 netL53 1.6131729899606437e-10
Rbbr53 netL53 0 -848378.3475621922
Cbr53 netL53 0 2.3706783331454107e-22

* Branch 54
Rabr54 node_3 netRa54 566.3950148058491
Lbr54 netRa54 netL54 -1.6670623090085387e-11
Rbbr54 netL54 0 -635864.6094211424
Cbr54 netL54 0 -3.481006455673002e-20

* Branch 55
Rabr55 node_3 netRa55 19657.447574867336
Lbr55 netRa55 netL55 -1.0620714900093147e-11
Rbbr55 netL55 0 -32018.52828818707
Cbr55 netL55 0 -1.6773965148785555e-20

* Branch 56
Rabr56 node_3 netRa56 -82125.77790582311
Lbr56 netRa56 netL56 -4.567529204825584e-11
Rbbr56 netL56 0 123670.53856281265
Cbr56 netL56 0 -4.524046225009588e-21

* Branch 57
Rabr57 node_3 netRa57 819521.4165067065
Lbr57 netRa57 netL57 -1.592609752573372e-10
Rbbr57 netL57 0 -857719.8980309363
Cbr57 netL57 0 -2.261025195760367e-22

* Branch 58
Rabr58 node_3 netRa58 -94338.28564999424
Lbr58 netRa58 netL58 2.5181722266963944e-11
Rbbr58 netL58 0 109559.91890533347
Cbr58 netL58 0 2.4295645355637234e-21

* Branch 59
Rabr59 node_3 netRa59 -1908.3400757853994
Lbr59 netRa59 netL59 6.3110755395601624e-12
Rbbr59 netL59 0 26598.529717797348
Cbr59 netL59 0 1.202113484233824e-19

* Branch 60
Rabr60 node_3 netRa60 -55646.8706501063
Lbr60 netRa60 netL60 2.602556274245664e-11
Rbbr60 netL60 0 77021.02937237329
Cbr60 netL60 0 6.0432319213262036e-21

* Branch 61
Rabr61 node_3 netRa61 -5574.461770290588
Lbr61 netRa61 netL61 6.270097055532567e-12
Rbbr61 netL61 0 14700.334136050498
Cbr61 netL61 0 7.565058988189338e-20

* Branch 62
Rabr62 node_3 netRa62 -208854270.0200669
Lbr62 netRa62 netL62 -1.1244627317067904e-09
Rbbr62 netL62 0 208866834.318225
Cbr62 netL62 0 -2.5778335458683116e-26

* Branch 63
Rabr63 node_3 netRa63 19658.292150439323
Lbr63 netRa63 netL63 -7.809969819697452e-12
Rbbr63 netL63 0 -27629.978021287712
Cbr63 netL63 0 -1.432382679796094e-20

* Branch 64
Rabr64 node_3 netRa64 -113.21817609194218
Lbr64 netRa64 netL64 4.416857368617736e-12
Rbbr64 netL64 0 271952.0135065887
Cbr64 netL64 0 1.0524494622820523e-19

* Branch 65
Rabr65 node_3 netRa65 660.0951179218108
Lbr65 netRa65 netL65 9.166401219420345e-12
Rbbr65 netL65 0 -117928.08522334769
Cbr65 netL65 0 1.3510409117075225e-19

* Branch 66
Rabr66 node_3 netRa66 -22425.1967646291
Lbr66 netRa66 netL66 -2.4754772333535382e-11
Rbbr66 netL66 0 72374.23007215871
Cbr66 netL66 0 -1.53808008818351e-20

* Branch 67
Rabr67 node_3 netRa67 -52200.564463879266
Lbr67 netRa67 netL67 2.9752643245771814e-11
Rbbr67 netL67 0 73748.82003750395
Cbr67 netL67 0 7.699069746436306e-21

* Branch 68
Rabr68 node_3 netRa68 -4178.08803981318
Lbr68 netRa68 netL68 1.1874219440110635e-11
Rbbr68 netL68 0 35190.643083431
Cbr68 netL68 0 7.928968697926669e-20

* Branch 69
Rabr69 node_3 netRa69 4102.799262823536
Lbr69 netRa69 netL69 1.1946613006380417e-11
Rbbr69 netL69 0 -33704.622509612775
Cbr69 netL69 0 8.802575970824901e-20

* Branch 70
Rabr70 node_3 netRa70 -3331.662960864198
Lbr70 netRa70 netL70 -1.12199432763327e-11
Rbbr70 netL70 0 22792.10917358626
Cbr70 netL70 0 -1.508871483378072e-19

* Branch 71
Rabr71 node_3 netRa71 -7779.313270344974
Lbr71 netRa71 netL71 -3.902332994233708e-11
Rbbr71 netL71 0 95796.45368421468
Cbr71 netL71 0 -5.3998341843266715e-20

* Branch 72
Rabr72 node_3 netRa72 -126563.2457594983
Lbr72 netRa72 netL72 6.76113300059472e-11
Rbbr72 netL72 0 168176.80581797892
Cbr72 netL72 0 3.167685025705919e-21

* Branch 73
Rabr73 node_3 netRa73 5908.948472817667
Lbr73 netRa73 netL73 -2.3773391008376168e-11
Rbbr73 netL73 0 -91521.67500798537
Cbr73 netL73 0 -4.307367971723066e-20

* Branch 74
Rabr74 node_3 netRa74 -11664.789129295415
Lbr74 netRa74 netL74 -1.9830052402407867e-11
Rbbr74 netL74 0 94861.8685555186
Cbr74 netL74 0 -1.8064564114236003e-20

* Branch 75
Rabr75 node_3 netRa75 -1430.613144241863
Lbr75 netRa75 netL75 -1.5633559686599608e-11
Rbbr75 netL75 0 87575.8694076096
Cbr75 netL75 0 -1.3102081645931242e-19

* Branch 76
Rabr76 node_3 netRa76 -11132.37565677436
Lbr76 netRa76 netL76 1.969473520918201e-11
Rbbr76 netL76 0 52455.38835457896
Cbr76 netL76 0 3.352158311922477e-20

* Branch 77
Rabr77 node_3 netRa77 -1882.9896568015572
Lbr77 netRa77 netL77 -2.5772489168066096e-11
Rbbr77 netL77 0 170898.39459224924
Cbr77 netL77 0 -8.37663188319879e-20

* Branch 78
Rabr78 node_3 netRa78 4648.095999603221
Lbr78 netRa78 netL78 1.34240059915759e-11
Rbbr78 netL78 0 -42565.914464047586
Cbr78 netL78 0 6.845729910249711e-20

* Branch 79
Rabr79 node_3 netRa79 -10620.901617244976
Lbr79 netRa79 netL79 -1.0009919077059451e-11
Rbbr79 netL79 0 35797.25757714302
Cbr79 netL79 0 -2.6403973662787268e-20

* Branch 80
Rabr80 node_3 netRa80 -140.4679155477281
Lbr80 netRa80 netL80 1.861225430919012e-11
Rbbr80 netL80 0 1907252.463671945
Cbr80 netL80 0 4.979971588657969e-20

* Branch 81
Rabr81 node_3 netRa81 -33897.11797217289
Lbr81 netRa81 netL81 -3.201543002346992e-11
Rbbr81 netL81 0 52860.562935525195
Cbr81 netL81 0 -1.7910492153647747e-20

* Branch 82
Rabr82 node_3 netRa82 -382.406190286069
Lbr82 netRa82 netL82 1.1601397685903915e-11
Rbbr82 netL82 0 372423.4535382531
Cbr82 netL82 0 7.732149741717385e-20

* Branch 83
Rabr83 node_3 netRa83 1934.091124950324
Lbr83 netRa83 netL83 8.639959878470396e-12
Rbbr83 netL83 0 -42031.13404790651
Cbr83 netL83 0 1.068491897021234e-19

* Branch 84
Rabr84 node_3 netRa84 2843.0958678666925
Lbr84 netRa84 netL84 9.008188412711379e-12
Rbbr84 netL84 0 -21655.403127165413
Cbr84 netL84 0 1.468364382010058e-19

* Branch 85
Rabr85 node_3 netRa85 61261.194863667595
Lbr85 netRa85 netL85 -3.499511568970905e-11
Rbbr85 netL85 0 -113536.01313145409
Cbr85 netL85 0 -5.030344898620775e-21

* Branch 86
Rabr86 node_3 netRa86 -2278.3305575901504
Lbr86 netRa86 netL86 -7.2526398365032086e-12
Rbbr86 netL86 0 14490.931180150208
Cbr86 netL86 0 -2.199147966904981e-19

* Branch 87
Rabr87 node_3 netRa87 10051.122254621238
Lbr87 netRa87 netL87 -4.59205462225021e-11
Rbbr87 netL87 0 -454101.53511619766
Cbr87 netL87 0 -1.0055928165456472e-20

* Branch 88
Rabr88 node_3 netRa88 9178.743961793825
Lbr88 netRa88 netL88 1.426834310794739e-11
Rbbr88 netL88 0 -31459.081111149637
Cbr88 netL88 0 4.941918055812379e-20

* Branch 89
Rabr89 node_3 netRa89 1582.7605512986404
Lbr89 netRa89 netL89 1.7410753890702335e-11
Rbbr89 netL89 0 -110625.06139283841
Cbr89 netL89 0 9.991975878799869e-20

* Branch 90
Rabr90 node_3 netRa90 41979.60182451287
Lbr90 netRa90 netL90 2.8620141452113847e-11
Rbbr90 netL90 0 -58903.46279760889
Cbr90 netL90 0 1.1578561568850634e-20

* Branch 91
Rabr91 node_3 netRa91 12382.788787657506
Lbr91 netRa91 netL91 2.3611596422814582e-11
Rbbr91 netL91 0 -38592.4890423961
Cbr91 netL91 0 4.9479114805544884e-20

* Branch 92
Rabr92 node_3 netRa92 -1256.7615372715763
Lbr92 netRa92 netL92 -4.9990835855938634e-12
Rbbr92 netL92 0 12226.308798935861
Cbr92 netL92 0 -3.2634314314645883e-19

* Branch 93
Rabr93 node_3 netRa93 279.0439405965204
Lbr93 netRa93 netL93 -1.2197596409177502e-11
Rbbr93 netL93 0 -310496.40278486995
Cbr93 netL93 0 -1.3581575122835072e-19

* Branch 94
Rabr94 node_3 netRa94 1144925.478269048
Lbr94 netRa94 netL94 1.7374706625993656e-10
Rbbr94 netL94 0 -1163025.8708796403
Cbr94 netL94 0 1.305138084100681e-22

* Branch 95
Rabr95 node_3 netRa95 22864.24556372943
Lbr95 netRa95 netL95 1.6456949622476627e-11
Rbbr95 netL95 0 -33491.43751522078
Cbr95 netL95 0 2.1516607533347882e-20

* Branch 96
Rabr96 node_3 netRa96 15.543059276235578
Lbr96 netRa96 netL96 5.021526753311332e-12
Rbbr96 netL96 0 -2719924.3512697928
Cbr96 netL96 0 3.0827590511612208e-19

* Branch 97
Rabr97 node_3 netRa97 39283.76018709307
Lbr97 netRa97 netL97 -3.0148021789651094e-11
Rbbr97 netL97 0 -55897.18137790201
Cbr97 netL97 0 -1.3700086679410992e-20

* Branch 98
Rabr98 node_3 netRa98 7414.9420292956875
Lbr98 netRa98 netL98 7.757962886310703e-12
Rbbr98 netL98 0 -13675.123244706172
Cbr98 netL98 0 7.758030553577455e-20

* Branch 99
Rabr99 node_3 netRa99 265131.98460130545
Lbr99 netRa99 netL99 1.530772114988819e-11
Rbbr99 netL99 0 -268403.6373007013
Cbr99 netL99 0 2.177785711855199e-22

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 398873.51095929305
Lbr0 netRa0 netL0 3.0471979664180646e-10
Rbbr0 netL0 node_4 -1110984.8600571295
Cbr0 netL0 node_4 1.2904029766764939e-21

* Branch 1
Rabr1 node_3 netRa1 509175.37508513365
Lbr1 netRa1 netL1 2.9782390508305445e-10
Rbbr1 netL1 node_4 -952404.7146118778
Cbr1 netL1 node_4 9.40993145085153e-22

* Branch 2
Rabr2 node_3 netRa2 715762.7696505741
Lbr2 netRa2 netL2 2.90100202930894e-10
Rbbr2 netL2 node_4 -976039.9262727405
Cbr2 netL2 node_4 5.369417836802333e-22

* Branch 3
Rabr3 node_3 netRa3 2564016.3312233565
Lbr3 netRa3 netL3 4.4125793614753385e-10
Rbbr3 netL3 node_4 -2709461.954818928
Cbr3 netL3 node_4 6.917837080579137e-23

* Branch 4
Rabr4 node_3 netRa4 6423881.0710014505
Lbr4 netRa4 netL4 -5.38585098168983e-10
Rbbr4 netL4 node_4 -6503196.017466893
Cbr4 netL4 node_4 -1.2556520592107094e-23

* Branch 5
Rabr5 node_3 netRa5 74876.36814222953
Lbr5 netRa5 netL5 2.212586124472378e-11
Rbbr5 netL5 node_4 -92145.38382049455
Cbr5 netL5 node_4 3.2568288421072078e-21

* Branch 6
Rabr6 node_3 netRa6 12292468.142260674
Lbr6 netRa6 netL6 -3.77621417671764e-10
Rbbr6 netL6 node_4 -12318919.537490837
Cbr6 netL6 node_4 -2.4898476719488232e-24

* Branch 7
Rabr7 node_3 netRa7 495833.0826537779
Lbr7 netRa7 netL7 6.149421440391361e-11
Rbbr7 netL7 node_4 -514961.0062789791
Cbr7 netL7 node_4 2.4230668383780152e-22

* Branch 8
Rabr8 node_3 netRa8 272649.4845222537
Lbr8 netRa8 netL8 4.085431809826263e-11
Rbbr8 netL8 node_4 -288373.3882229852
Cbr8 netL8 node_4 5.218533824667615e-22

* Branch 9
Rabr9 node_3 netRa9 -2193.727382116148
Lbr9 netRa9 netL9 4.298727538352144e-12
Rbbr9 netL9 node_4 27879.95297578737
Cbr9 netL9 node_4 6.772097450990663e-20

* Branch 10
Rabr10 node_3 netRa10 275093.4351310532
Lbr10 netRa10 netL10 -7.086990598454968e-11
Rbbr10 netL10 node_4 -311815.7816703982
Cbr10 netL10 node_4 -8.222866066968945e-22

* Branch 11
Rabr11 node_3 netRa11 8580.110924122346
Lbr11 netRa11 netL11 5.565910456507448e-12
Rbbr11 netL11 node_4 -20014.85896897255
Cbr11 netL11 node_4 3.274719071570707e-20

* Branch 12
Rabr12 node_3 netRa12 243.19188730024086
Lbr12 netRa12 netL12 6.584869592189017e-12
Rbbr12 netL12 node_4 -888276.1369028292
Cbr12 netL12 node_4 5.200831946692793e-20

* Branch 13
Rabr13 node_3 netRa13 524004.2623636852
Lbr13 netRa13 netL13 -1.0593180120807677e-10
Rbbr13 netL13 node_4 -536039.5485405279
Cbr13 netL13 node_4 -3.7606380886884904e-22

* Branch 14
Rabr14 node_3 netRa14 1660.7021422382948
Lbr14 netRa14 netL14 -1.0516130075762118e-11
Rbbr14 netL14 node_4 -32398.777419211427
Cbr14 netL14 node_4 -1.7949605186922491e-19

* Branch 15
Rabr15 node_3 netRa15 49617.69888148072
Lbr15 netRa15 netL15 2.764640559712018e-11
Rbbr15 netL15 node_4 -57133.07918446901
Cbr15 netL15 node_4 9.828032901544308e-21

* Branch 16
Rabr16 node_3 netRa16 -3495.1884184949768
Lbr16 netRa16 netL16 1.276027598377326e-11
Rbbr16 netL16 node_4 27599.053002068882
Cbr16 netL16 node_4 1.260267568186679e-19

* Branch 17
Rabr17 node_3 netRa17 987.9794209512057
Lbr17 netRa17 netL17 3.68666247333919e-12
Rbbr17 netL17 node_4 -47680.50473649565
Cbr17 netL17 node_4 8.236754992266197e-20

* Branch 18
Rabr18 node_3 netRa18 -338690.09813419764
Lbr18 netRa18 netL18 -7.092236825315624e-11
Rbbr18 netL18 node_4 346466.6775132901
Cbr18 netL18 node_4 -6.060745753089306e-22

* Branch 19
Rabr19 node_3 netRa19 1281.9001012930257
Lbr19 netRa19 netL19 1.0758899513792765e-11
Rbbr19 netL19 node_4 -48364.27225090489
Cbr19 netL19 node_4 1.9467537910880487e-19

* Branch 20
Rabr20 node_3 netRa20 -19403.159416359566
Lbr20 netRa20 netL20 2.0867594027442174e-11
Rbbr20 netL20 node_4 29277.06837158221
Cbr20 netL20 node_4 3.623169964494696e-20

* Branch 21
Rabr21 node_3 netRa21 -42855.89777553581
Lbr21 netRa21 netL21 -4.270380194750108e-11
Rbbr21 netL21 node_4 61308.370383406975
Cbr21 netL21 node_4 -1.646422952288311e-20

* Branch 22
Rabr22 node_3 netRa22 -22116.4080317273
Lbr22 netRa22 netL22 2.2126958150120703e-11
Rbbr22 netL22 node_4 35409.9670172713
Cbr22 netL22 node_4 2.790081381578753e-20

* Branch 23
Rabr23 node_3 netRa23 1410.3333640102555
Lbr23 netRa23 netL23 3.781132155480797e-12
Rbbr23 netL23 node_4 -35910.06907400714
Cbr23 netL23 node_4 7.721243098941418e-20

* Branch 24
Rabr24 node_3 netRa24 -5038.856914069673
Lbr24 netRa24 netL24 -1.0056907641047006e-11
Rbbr24 netL24 node_4 17081.83153497011
Cbr24 netL24 node_4 -1.1973255375315392e-19

* Branch 25
Rabr25 node_3 netRa25 8614.724809446521
Lbr25 netRa25 netL25 6.2365786432750524e-12
Rbbr25 netL25 node_4 -20713.086526036106
Cbr25 netL25 node_4 3.5241966886442524e-20

* Branch 26
Rabr26 node_3 netRa26 132542933.33255747
Lbr26 netRa26 netL26 1.351386063711215e-09
Rbbr26 netL26 node_4 -132554793.16046108
Cbr26 netL26 node_4 7.692673677210955e-26

* Branch 27
Rabr27 node_3 netRa27 1484.745186210315
Lbr27 netRa27 netL27 3.817603655007603e-12
Rbbr27 netL27 node_4 -35419.80124414502
Cbr27 netL27 node_4 7.474233268573572e-20

* Branch 28
Rabr28 node_3 netRa28 120145.35257173398
Lbr28 netRa28 netL28 -5.548368736269874e-11
Rbbr28 netL28 node_4 -166878.53130856575
Cbr28 netL28 node_4 -2.754937779930646e-21

* Branch 29
Rabr29 node_3 netRa29 2024931.471376494
Lbr29 netRa29 netL29 -2.4842508828510915e-10
Rbbr29 netL29 node_4 -2054301.5666315367
Cbr29 netL29 node_4 -5.96493787332627e-23

* Branch 30
Rabr30 node_3 netRa30 1070.796325972997
Lbr30 netRa30 netL30 3.3317806489190504e-12
Rbbr30 netL30 node_4 -38384.80700087095
Cbr30 netL30 node_4 8.349741834952923e-20

* Branch 31
Rabr31 node_3 netRa31 1515.1487812813766
Lbr31 netRa31 netL31 4.251938150150052e-12
Rbbr31 netL31 node_4 -43447.10598519222
Cbr31 netL31 node_4 6.627885808515303e-20

* Branch 32
Rabr32 node_3 netRa32 697821729.7256773
Lbr32 netRa32 netL32 2.29281298144487e-09
Rbbr32 netL32 node_4 -697840213.4934381
Cbr32 netL32 node_4 4.7084828515703244e-27

* Branch 33
Rabr33 node_3 netRa33 -29195.32485675603
Lbr33 netRa33 netL33 -3.678059925527537e-11
Rbbr33 netL33 node_4 62566.74991976428
Cbr33 netL33 node_4 -2.0356891160583648e-20

* Branch 34
Rabr34 node_3 netRa34 -13231.357612945154
Lbr34 netRa34 netL34 -2.3658818595159732e-11
Rbbr34 netL34 node_4 42362.62488514695
Cbr34 netL34 node_4 -4.285972144542088e-20

* Branch 35
Rabr35 node_3 netRa35 -23939.329311732952
Lbr35 netRa35 netL35 -2.5228903089080825e-11
Rbbr35 netL35 node_4 41350.57620020239
Cbr35 netL35 node_4 -2.5711542197493006e-20

* Branch 36
Rabr36 node_3 netRa36 654618.2869528811
Lbr36 netRa36 netL36 -9.186523982536468e-11
Rbbr36 netL36 node_4 -683093.7429735843
Cbr36 netL36 node_4 -2.052217563325504e-22

* Branch 37
Rabr37 node_3 netRa37 -23361.793585376596
Lbr37 netRa37 netL37 -1.6895107697558555e-11
Rbbr37 netL37 node_4 32938.30937567782
Cbr37 netL37 node_4 -2.20724442041864e-20

* Branch 38
Rabr38 node_3 netRa38 53292.693849614894
Lbr38 netRa38 netL38 -4.67926987553795e-11
Rbbr38 netL38 node_4 -119633.22150282018
Cbr38 netL38 node_4 -7.294432112729523e-21

* Branch 39
Rabr39 node_3 netRa39 92762.36381696186
Lbr39 netRa39 netL39 -5.174787463116433e-11
Rbbr39 netL39 node_4 -143777.69134448515
Cbr39 netL39 node_4 -3.865054435262009e-21

* Branch 40
Rabr40 node_3 netRa40 27716.477212673923
Lbr40 netRa40 netL40 -4.136928439319189e-11
Rbbr40 netL40 node_4 -119183.06822015706
Cbr40 netL40 node_4 -1.241138979584921e-20

* Branch 41
Rabr41 node_3 netRa41 5771.040187209096
Lbr41 netRa41 netL41 4.176161248333406e-12
Rbbr41 netL41 node_4 -15115.438078521494
Cbr41 netL41 node_4 4.8075185673421956e-20

* Branch 42
Rabr42 node_3 netRa42 5645.294996995056
Lbr42 netRa42 netL42 3.920875304022036e-12
Rbbr42 netL42 node_4 -13737.382451488284
Cbr42 netL42 node_4 5.074834662887189e-20

* Branch 43
Rabr43 node_3 netRa43 -72087.87863001708
Lbr43 netRa43 netL43 2.1277990914476275e-11
Rbbr43 netL43 node_4 77596.18423850488
Cbr43 netL43 node_4 3.798103290822077e-21

* Branch 44
Rabr44 node_3 netRa44 2165.1398517606685
Lbr44 netRa44 netL44 9.791138356684313e-12
Rbbr44 netL44 node_4 -39917.993143950924
Cbr44 netL44 node_4 1.1544516768169423e-19

* Branch 45
Rabr45 node_3 netRa45 184295.2886668266
Lbr45 netRa45 netL45 -3.697920406003781e-11
Rbbr45 netL45 node_4 -189942.07318922837
Cbr45 netL45 node_4 -1.0555697412987648e-21

* Branch 46
Rabr46 node_3 netRa46 9754.181377097533
Lbr46 netRa46 netL46 5.241401067101355e-12
Rbbr46 netL46 node_4 -18280.943846151913
Cbr46 netL46 node_4 2.944919681018293e-20

* Branch 47
Rabr47 node_3 netRa47 -18377.15634269512
Lbr47 netRa47 netL47 1.8498329896191705e-11
Rbbr47 netL47 node_4 33354.09187589462
Cbr47 netL47 node_4 3.007496145176829e-20

* Branch 48
Rabr48 node_3 netRa48 -3734.5688229240964
Lbr48 netRa48 netL48 9.293120383094528e-12
Rbbr48 netL48 node_4 25329.591761174426
Cbr48 netL48 node_4 9.743810798940386e-20

* Branch 49
Rabr49 node_3 netRa49 -21169.18096298078
Lbr49 netRa49 netL49 -2.820611519119663e-11
Rbbr49 netL49 node_4 61432.994749974205
Cbr49 netL49 node_4 -2.177523283079867e-20

* Branch 50
Rabr50 node_3 netRa50 4241.83067495296
Lbr50 netRa50 netL50 -3.423337090291511e-11
Rbbr50 netL50 node_4 -349515.5823397453
Cbr50 netL50 node_4 -2.2594327640467378e-20

* Branch 51
Rabr51 node_3 netRa51 -21434.991561725088
Lbr51 netRa51 netL51 1.4589400033823132e-11
Rbbr51 netL51 node_4 30444.76593993226
Cbr51 netL51 node_4 2.2318077433876522e-20

* Branch 52
Rabr52 node_3 netRa52 -11384.585658977176
Lbr52 netRa52 netL52 -3.1124547655246094e-11
Rbbr52 netL52 node_4 111528.7093614051
Cbr52 netL52 node_4 -2.459007226691069e-20

* Branch 53
Rabr53 node_3 netRa53 12284.181467956614
Lbr53 netRa53 netL53 -3.618843209357563e-11
Rbbr53 netL53 node_4 -159017.44189639678
Cbr53 netL53 node_4 -1.8479669983163484e-20

* Branch 54
Rabr54 node_3 netRa54 70489.09814877166
Lbr54 netRa54 netL54 1.5418251363587192e-11
Rbbr54 netL54 node_4 -79675.48703749845
Cbr54 netL54 node_4 2.7455981732936963e-21

* Branch 55
Rabr55 node_3 netRa55 -107204.78779992055
Lbr55 netRa55 netL55 3.701987648700255e-11
Rbbr55 netL55 node_4 120612.56785692832
Cbr55 netL55 node_4 2.862592461146932e-21

* Branch 56
Rabr56 node_3 netRa56 51014.48161637029
Lbr56 netRa56 netL56 3.862528953269832e-11
Rbbr56 netL56 node_4 -69313.99292013203
Cbr56 netL56 node_4 1.0927112715880154e-20

* Branch 57
Rabr57 node_3 netRa57 25272.709745342712
Lbr57 netRa57 netL57 -3.487691575940704e-11
Rbbr57 netL57 node_4 -59556.177192734816
Cbr57 netL57 node_4 -2.316298042558738e-20

* Branch 58
Rabr58 node_3 netRa58 -48615.872496697666
Lbr58 netRa58 netL58 -5.084874214563481e-11
Rbbr58 netL58 node_4 83325.98452996476
Cbr58 netL58 node_4 -1.2552392067982533e-20

* Branch 59
Rabr59 node_3 netRa59 -23011.434987593515
Lbr59 netRa59 netL59 -4.745754631662135e-11
Rbbr59 netL59 node_4 89769.83058026701
Cbr59 netL59 node_4 -2.297402634739324e-20

* Branch 60
Rabr60 node_3 netRa60 942158.7778856627
Lbr60 netRa60 netL60 1.7803341363010597e-10
Rbbr60 netL60 node_4 -1024235.8599664782
Cbr60 netL60 node_4 1.8449223878401925e-22

* Branch 61
Rabr61 node_3 netRa61 512970.9066020212
Lbr61 netRa61 netL61 1.1183059956603572e-10
Rbbr61 netL61 node_4 -567102.3960245315
Cbr61 netL61 node_4 3.8442430116653935e-22

* Branch 62
Rabr62 node_3 netRa62 537835.1593188948
Lbr62 netRa62 netL62 1.457426433217764e-10
Rbbr62 netL62 node_4 -631988.2264533435
Cbr62 netL62 node_4 4.287798238996737e-22

* Branch 63
Rabr63 node_3 netRa63 -6671021.709745062
Lbr63 netRa63 netL63 3.611204482414208e-10
Rbbr63 netL63 node_4 6692975.517662771
Cbr63 netL63 node_4 8.087962897304813e-24

* Branch 64
Rabr64 node_3 netRa64 410699.82377465186
Lbr64 netRa64 netL64 9.863156826276637e-11
Rbbr64 netL64 node_4 -464568.8080753436
Cbr64 netL64 node_4 5.169507271491398e-22

* Branch 65
Rabr65 node_3 netRa65 377111.271814994
Lbr65 netRa65 netL65 9.711908434449062e-11
Rbbr65 netL65 node_4 -435356.07002251246
Cbr65 netL65 node_4 5.915604062236626e-22

* Branch 66
Rabr66 node_3 netRa66 342298.20365583524
Lbr66 netRa66 netL66 1.1167486249375908e-10
Rbbr66 netL66 node_4 -419350.71878545824
Cbr66 netL66 node_4 7.78010761650798e-22

* Branch 67
Rabr67 node_3 netRa67 276906.42727754073
Lbr67 netRa67 netL67 1.1180937086895681e-10
Rbbr67 netL67 node_4 -374760.532636597
Cbr67 netL67 node_4 1.0774739761796668e-21

* Branch 68
Rabr68 node_3 netRa68 309169.2133928326
Lbr68 netRa68 netL68 1.0230290953272195e-10
Rbbr68 netL68 node_4 -379003.00370530476
Cbr68 netL68 node_4 8.730961830925534e-22

* Branch 69
Rabr69 node_3 netRa69 175553.75227333463
Lbr69 netRa69 netL69 6.760964488688484e-11
Rbbr69 netL69 node_4 -240545.89893478324
Cbr69 netL69 node_4 1.6010955243795738e-21

* Branch 70
Rabr70 node_3 netRa70 218650.09567356197
Lbr70 netRa70 netL70 9.922142834354813e-11
Rbbr70 netL70 node_4 -306954.23265744175
Cbr70 netL70 node_4 1.47843425414758e-21

* Branch 71
Rabr71 node_3 netRa71 210918.5082505645
Lbr71 netRa71 netL71 8.916094195405268e-11
Rbbr71 netL71 node_4 -286743.43603422795
Cbr71 netL71 node_4 1.4742977591404908e-21

* Branch 72
Rabr72 node_3 netRa72 210316.34545173383
Lbr72 netRa72 netL72 9.523316589686982e-11
Rbbr72 netL72 node_4 -290605.4250817536
Cbr72 netL72 node_4 1.5582300663936295e-21

* Branch 73
Rabr73 node_3 netRa73 186106.56485570467
Lbr73 netRa73 netL73 8.439144998651033e-11
Rbbr73 netL73 node_4 -259244.75584979297
Cbr73 netL73 node_4 1.7492337177182227e-21

* Branch 74
Rabr74 node_3 netRa74 107995.44860486622
Lbr74 netRa74 netL74 8.765914524832566e-11
Rbbr74 netL74 node_4 -230233.0484148678
Cbr74 netL74 node_4 3.525847472618752e-21

* Branch 75
Rabr75 node_3 netRa75 89881.2032073671
Lbr75 netRa75 netL75 8.501001556719727e-11
Rbbr75 netL75 node_4 -231825.32494699612
Cbr75 netL75 node_4 4.0802556449455675e-21

* Branch 76
Rabr76 node_3 netRa76 119374.44842097013
Lbr76 netRa76 netL76 8.232450470416709e-11
Rbbr76 netL76 node_4 -222324.68204436311
Cbr76 netL76 node_4 3.102161531736158e-21

* Branch 77
Rabr77 node_3 netRa77 98410.98211400138
Lbr77 netRa77 netL77 8.360575879677054e-11
Rbbr77 netL77 node_4 -217115.24268218837
Cbr77 netL77 node_4 3.913313626677332e-21

* Branch 78
Rabr78 node_3 netRa78 54100.31259037732
Lbr78 netRa78 netL78 7.599123304828912e-11
Rbbr78 netL78 node_4 -222732.59579688127
Cbr78 netL78 node_4 6.307461612768345e-21

* Branch 79
Rabr79 node_3 netRa79 62890.066583488995
Lbr79 netRa79 netL79 7.147306999016274e-11
Rbbr79 netL79 node_4 -194902.9226389134
Cbr79 netL79 node_4 5.83180940261499e-21

* Branch 80
Rabr80 node_3 netRa80 48207.499174950484
Lbr80 netRa80 netL80 7.593427195512755e-11
Rbbr80 netL80 node_4 -231814.2986386258
Cbr80 netL80 node_4 6.796234746973914e-21

* Branch 81
Rabr81 node_3 netRa81 77220.30048117049
Lbr81 netRa81 netL81 1.6491380617645e-11
Rbbr81 netL81 node_4 -87023.58582649032
Cbr81 netL81 node_4 2.4541466452961468e-21

* Branch 82
Rabr82 node_3 netRa82 19722.497536335286
Lbr82 netRa82 netL82 7.38931175141661e-11
Rbbr82 netL82 node_4 -432611.68367477844
Cbr82 netL82 node_4 8.664750337008412e-21

* Branch 83
Rabr83 node_3 netRa83 8808.00880405428
Lbr83 netRa83 netL83 8.218968771853252e-11
Rbbr83 netL83 node_4 -1120028.3369449924
Cbr83 netL83 node_4 8.341434322623781e-21

* Branch 84
Rabr84 node_3 netRa84 2124.570616696067
Lbr84 netRa84 netL84 8.38111795327403e-11
Rbbr84 netL84 node_4 -4669360.187064798
Cbr84 netL84 node_4 8.492711345010413e-21

* Branch 85
Rabr85 node_3 netRa85 -45463.604946781175
Lbr85 netRa85 netL85 8.440490742718242e-11
Rbbr85 netL85 node_4 258856.45104117243
Cbr85 netL85 node_4 7.170248178996232e-21

* Branch 86
Rabr86 node_3 netRa86 -74650.12498596187
Lbr86 netRa86 netL86 9.080593220015899e-11
Rbbr86 netL86 node_4 220493.9924343179
Cbr86 netL86 node_4 5.515844609646017e-21

* Branch 87
Rabr87 node_3 netRa87 -90702.82774915396
Lbr87 netRa87 netL87 8.772753687711933e-11
Rbbr87 netL87 node_4 199266.0614439805
Cbr87 netL87 node_4 4.8531220867975245e-21

* Branch 88
Rabr88 node_3 netRa88 -127167.1605608218
Lbr88 netRa88 netL88 8.49427645051907e-11
Rbbr88 netL88 node_4 197485.00496164666
Cbr88 netL88 node_4 3.3819692636210225e-21

* Branch 89
Rabr89 node_3 netRa89 -135937.3235273126
Lbr89 netRa89 netL89 8.199337529211157e-11
Rbbr89 netL89 node_4 195270.80891566753
Cbr89 netL89 node_4 3.0885663286575346e-21

* Branch 90
Rabr90 node_3 netRa90 -860715.4975286638
Lbr90 netRa90 netL90 9.941972729687376e-11
Rbbr90 netL90 node_4 873186.3467041356
Cbr90 netL90 node_4 1.3228050973578626e-22

* Branch 91
Rabr91 node_3 netRa91 -1681808.1526301135
Lbr91 netRa91 netL91 8.79395061745071e-11
Rbbr91 netL91 node_4 1686320.6027827559
Cbr91 netL91 node_4 3.100716564568507e-23

* Branch 92
Rabr92 node_3 netRa92 -108974.07929851423
Lbr92 netRa92 netL92 5.189145395808948e-11
Rbbr92 netL92 node_4 137662.4658472718
Cbr92 netL92 node_4 3.458601443344144e-21

* Branch 93
Rabr93 node_3 netRa93 33542.14519769747
Lbr93 netRa93 netL93 3.25003081757222e-11
Rbbr93 netL93 node_4 -113961.00016846429
Cbr93 netL93 node_4 8.504680250035516e-21

* Branch 94
Rabr94 node_3 netRa94 37190.354799685345
Lbr94 netRa94 netL94 1.5374949690212623e-11
Rbbr94 netL94 node_4 -53777.00759676526
Cbr94 netL94 node_4 7.688523069177367e-21

* Branch 95
Rabr95 node_3 netRa95 -128543.1133111197
Lbr95 netRa95 netL95 3.296309800481551e-11
Rbbr95 netL95 node_4 137108.56563399688
Cbr95 netL95 node_4 1.8700302607711464e-21

* Branch 96
Rabr96 node_3 netRa96 -5693.3813067416795
Lbr96 netRa96 netL96 3.1859018007724233e-12
Rbbr96 netL96 node_4 12061.447652388835
Cbr96 netL96 node_4 4.6357774996466774e-20

* Branch 97
Rabr97 node_3 netRa97 9252.579120649105
Lbr97 netRa97 netL97 5.719163261429887e-12
Rbbr97 netL97 node_4 -19310.681553862516
Cbr97 netL97 node_4 3.203786506577267e-20

* Branch 98
Rabr98 node_3 netRa98 13535.876587169132
Lbr98 netRa98 netL98 4.789417705286661e-12
Rbbr98 netL98 node_4 -18045.076009456643
Cbr98 netL98 node_4 1.9619294923814327e-20

* Branch 99
Rabr99 node_3 netRa99 5868.200222483408
Lbr99 netRa99 netL99 3.198375168263396e-12
Rbbr99 netL99 node_4 -10922.38438248265
Cbr99 netL99 node_4 4.9987815229893056e-20

.ends


* Y'44
.subckt yp44 node_4 0
* Branch 0
Rabr0 node_4 netRa0 6583.987242104647
Lbr0 netRa0 netL0 4.739774817202493e-12
Rbbr0 netL0 0 -20068.60648842926
Cbr0 netL0 0 3.9640257743112337e-20

* Branch 1
Rabr1 node_4 netRa1 12973.509376221087
Lbr1 netRa1 netL1 5.796916700699978e-12
Rbbr1 netL1 0 -22712.97991604763
Cbr1 netL1 0 2.0764998272464022e-20

* Branch 2
Rabr2 node_4 netRa2 51091.70889514828
Lbr2 netRa2 netL2 1.0393082849354237e-11
Rbbr2 netL2 0 -58743.41256169984
Cbr2 netL2 0 3.537910566961956e-21

* Branch 3
Rabr3 node_4 netRa3 1255529.0758797515
Lbr3 netRa3 netL3 5.765942741269628e-11
Rbbr3 netL3 0 -1264883.1114508263
Cbr3 netL3 0 3.6479956679279904e-23

* Branch 4
Rabr4 node_4 netRa4 590.7854034989957
Lbr4 netRa4 netL4 -2.2474131433288803e-12
Rbbr4 netL4 0 -24128.4267982664
Cbr4 netL4 0 -1.2473066230325413e-19

* Branch 5
Rabr5 node_4 netRa5 1853.2796124957524
Lbr5 netRa5 netL5 2.487798314929067e-12
Rbbr5 netL5 0 -14153.737173731275
Cbr5 netL5 0 1.0225426051790698e-19

* Branch 6
Rabr6 node_4 netRa6 -1783.0412057021463
Lbr6 netRa6 netL6 -5.3480988076578514e-12
Rbbr6 netL6 0 14042.027334836837
Cbr6 netL6 0 -2.4998087185773173e-19

* Branch 7
Rabr7 node_4 netRa7 -234249.90051575587
Lbr7 netRa7 netL7 -6.255762107407988e-11
Rbbr7 netL7 0 246338.8071766063
Cbr7 netL7 0 -1.0939865119393986e-21

* Branch 8
Rabr8 node_4 netRa8 -415445.6012042646
Lbr8 netRa8 netL8 -8.91077350783523e-11
Rbbr8 netL8 0 429226.0784617746
Cbr8 netL8 0 -5.03006802066108e-22

* Branch 9
Rabr9 node_4 netRa9 -24851.01152332764
Lbr9 netRa9 netL9 -1.924151738845028e-11
Rbbr9 netL9 0 35491.18810061074
Cbr9 netL9 0 -2.2332531107242027e-20

* Branch 10
Rabr10 node_4 netRa10 -9007.271700902653
Lbr10 netRa10 netL10 -9.160529520325525e-12
Rbbr10 netL10 0 43365.60639496546
Cbr10 netL10 0 -2.415602189215633e-20

* Branch 11
Rabr11 node_4 netRa11 -211523.65183563763
Lbr11 netRa11 netL11 -7.083026983916647e-11
Rbbr11 netL11 0 228620.53979755315
Cbr11 netL11 0 -1.478674342937133e-21

* Branch 12
Rabr12 node_4 netRa12 135001.52433323502
Lbr12 netRa12 netL12 1.3478129370278057e-11
Rbbr12 netL12 0 -139430.28058706078
Cbr12 netL12 0 7.180137664350316e-22

* Branch 13
Rabr13 node_4 netRa13 -9034.082852155105
Lbr13 netRa13 netL13 3.4466945501763126e-12
Rbbr13 netL13 0 13276.637802049232
Cbr13 netL13 0 2.84389571206957e-20

* Branch 14
Rabr14 node_4 netRa14 -4475673.672604358
Lbr14 netRa14 netL14 3.432614126895429e-10
Rbbr14 netL14 0 4494492.75163125
Cbr14 netL14 0 1.70315886651873e-23

* Branch 15
Rabr15 node_4 netRa15 39924.53905839212
Lbr15 netRa15 netL15 1.091834646015091e-11
Rbbr15 netL15 0 -48790.13761501761
Cbr15 netL15 0 5.641090801184219e-21

* Branch 16
Rabr16 node_4 netRa16 -1881.2718830240792
Lbr16 netRa16 netL16 4.266012901659271e-12
Rbbr16 netL16 0 25192.23939292238
Cbr16 netL16 0 8.551250292571003e-20

* Branch 17
Rabr17 node_4 netRa17 25415.156841730295
Lbr17 netRa17 netL17 -4.209152754579472e-11
Rbbr17 netL17 0 -152559.62922739872
Cbr17 netL17 0 -1.046868070559649e-20

* Branch 18
Rabr18 node_4 netRa18 12755.846554504882
Lbr18 netRa18 netL18 5.3187045948400984e-12
Rbbr18 netL18 0 -19054.323097895118
Cbr18 netL18 0 2.2085703336850904e-20

* Branch 19
Rabr19 node_4 netRa19 -27767.987681117593
Lbr19 netRa19 netL19 -2.722517933456497e-11
Rbbr19 netL19 0 74970.9474841553
Cbr19 netL19 0 -1.3366353957140455e-20

* Branch 20
Rabr20 node_4 netRa20 1835.981368398053
Lbr20 netRa20 netL20 9.282094697349891e-12
Rbbr20 netL20 0 -99488.43793454861
Cbr20 netL20 0 5.701506129457493e-20

* Branch 21
Rabr21 node_4 netRa21 -3660.0975967302998
Lbr21 netRa21 netL21 4.7923456656255466e-12
Rbbr21 netL21 0 18743.50060159011
Cbr21 netL21 0 6.794612279553338e-20

* Branch 22
Rabr22 node_4 netRa22 -117973.14644454901
Lbr22 netRa22 netL22 2.975849472182388e-11
Rbbr22 netL22 0 130102.69640274662
Cbr22 netL22 0 1.928675243816373e-21

* Branch 23
Rabr23 node_4 netRa23 16959.93793300939
Lbr23 netRa23 netL23 1.4246307546730734e-11
Rbbr23 netL23 0 -42085.75118279785
Cbr23 netL23 0 2.0307365012771684e-20

* Branch 24
Rabr24 node_4 netRa24 127266.3249839229
Lbr24 netRa24 netL24 2.123224128544568e-11
Rbbr24 netL24 0 -137479.09128074546
Cbr24 netL24 0 1.2176277311611946e-21

* Branch 25
Rabr25 node_4 netRa25 1011.0926496444109
Lbr25 netRa25 netL25 4.832914781364911e-12
Rbbr25 netL25 0 -67141.20521410108
Cbr25 netL25 0 7.863288465921565e-20

* Branch 26
Rabr26 node_4 netRa26 4028.505305268646
Lbr26 netRa26 netL26 1.278393173751902e-11
Rbbr26 netL26 0 -77613.0424461148
Cbr26 netL26 0 4.359365453765586e-20

* Branch 27
Rabr27 node_4 netRa27 2021.0111824692308
Lbr27 netRa27 netL27 1.0540268090130244e-11
Rbbr27 netL27 0 -97387.02407233047
Cbr27 netL27 0 5.96087625755398e-20

* Branch 28
Rabr28 node_4 netRa28 -8648.813234984584
Lbr28 netRa28 netL28 1.0585957066236164e-11
Rbbr28 netL28 0 31555.441287462945
Cbr28 netL28 0 3.788974897409559e-20

* Branch 29
Rabr29 node_4 netRa29 23872.29542017824
Lbr29 netRa29 netL29 -4.112573883672943e-11
Rbbr29 netL29 0 -133317.2192923009
Cbr29 netL29 0 -1.2504860683258348e-20

* Branch 30
Rabr30 node_4 netRa30 589.8771396095946
Lbr30 netRa30 netL30 2.879680760828251e-12
Rbbr30 netL30 0 -43502.39949520429
Cbr30 netL30 0 1.2390900682318876e-19

* Branch 31
Rabr31 node_4 netRa31 27818.777496833773
Lbr31 netRa31 netL31 -1.1668688153936435e-11
Rbbr31 netL31 0 -42435.63472221702
Cbr31 netL31 0 -9.806200443514643e-21

* Branch 32
Rabr32 node_4 netRa32 333.77507272058796
Lbr32 netRa32 netL32 4.252877626834164e-12
Rbbr32 netL32 0 -168920.52247021068
Cbr32 netL32 0 9.912971740051912e-20

* Branch 33
Rabr33 node_4 netRa33 3368.0285750001613
Lbr33 netRa33 netL33 4.9104228254630135e-12
Rbbr33 netL33 0 -22872.29248695531
Cbr33 netL33 0 6.551492637045396e-20

* Branch 34
Rabr34 node_4 netRa34 43098.15573314111
Lbr34 netRa34 netL34 -2.0845431020917184e-11
Rbbr34 netL34 0 -69937.4272183029
Cbr34 netL34 0 -6.854546222884e-21

* Branch 35
Rabr35 node_4 netRa35 -1690.3872432635112
Lbr35 netRa35 netL35 -9.624271401078086e-12
Rbbr35 netL35 0 71023.83751757327
Cbr35 netL35 0 -8.956527328883939e-20

* Branch 36
Rabr36 node_4 netRa36 -247287.09259293866
Lbr36 netRa36 netL36 3.9941797911281956e-11
Rbbr36 netL36 0 255510.69766334747
Cbr36 netL36 0 6.302929490449411e-22

* Branch 37
Rabr37 node_4 netRa37 1276.5013581761739
Lbr37 netRa37 netL37 3.0384124971301054e-12
Rbbr37 netL37 0 -24667.018311171123
Cbr37 netL37 0 1.0073562761530406e-19

* Branch 38
Rabr38 node_4 netRa38 -7506.885604714724
Lbr38 netRa38 netL38 -2.556706021449299e-11
Rbbr38 netL38 0 141907.76925434376
Cbr38 netL38 0 -2.5523365615290248e-20

* Branch 39
Rabr39 node_4 netRa39 -16893.078900044344
Lbr39 netRa39 netL39 1.2709879852533702e-11
Rbbr39 netL39 0 31279.045921497967
Cbr39 netL39 0 2.37423618682013e-20

* Branch 40
Rabr40 node_4 netRa40 -79928.80828509369
Lbr40 netRa40 netL40 -2.599619343188379e-11
Rbbr40 netL40 0 91543.95890498221
Cbr40 netL40 0 -3.572985313787726e-21

* Branch 41
Rabr41 node_4 netRa41 -164576.77663255247
Lbr41 netRa41 netL41 -3.88109460767844e-11
Rbbr41 netL41 0 170264.59843556775
Cbr41 netL41 0 -1.3905941550884937e-21

* Branch 42
Rabr42 node_4 netRa42 2129.095031616663
Lbr42 netRa42 netL42 -1.4692442246073525e-11
Rbbr42 netL42 0 -116262.34590138505
Cbr42 netL42 0 -5.330279508522681e-20

* Branch 43
Rabr43 node_4 netRa43 -69700.63200680552
Lbr43 netRa43 netL43 2.75917272270792e-11
Rbbr43 netL43 0 88874.0404653333
Cbr43 netL43 0 4.426130230147391e-21

* Branch 44
Rabr44 node_4 netRa44 -449341.4472530656
Lbr44 netRa44 netL44 -5.075559933822884e-11
Rbbr44 netL44 0 455333.3697700256
Cbr44 netL44 0 -2.485148734064224e-22

* Branch 45
Rabr45 node_4 netRa45 5449.634577112965
Lbr45 netRa45 netL45 7.516525908426203e-12
Rbbr45 netL45 0 -29071.965871632525
Cbr45 netL45 0 4.849734886829201e-20

* Branch 46
Rabr46 node_4 netRa46 14329.67939838028
Lbr46 netRa46 netL46 1.9785783820239797e-11
Rbbr46 netL46 0 -48275.85299161379
Cbr46 netL46 0 2.923127921265169e-20

* Branch 47
Rabr47 node_4 netRa47 -14945.76575260177
Lbr47 netRa47 netL47 1.3717793833335356e-11
Rbbr47 netL47 0 29728.481133438334
Cbr47 netL47 0 3.045440924635308e-20

* Branch 48
Rabr48 node_4 netRa48 -11799.988533361546
Lbr48 netRa48 netL48 8.167946555924931e-12
Rbbr48 netL48 0 24745.09358570478
Cbr48 netL48 0 2.7693682221736894e-20

* Branch 49
Rabr49 node_4 netRa49 -2112.411996376652
Lbr49 netRa49 netL49 1.145593114371418e-11
Rbbr49 netL49 0 77474.61889911068
Cbr49 netL49 0 6.487504473981757e-20

* Branch 50
Rabr50 node_4 netRa50 -6739.635923207433
Lbr50 netRa50 netL50 1.3780768871685644e-11
Rbbr50 netL50 0 52274.076904806374
Cbr50 netL50 0 3.802086621725646e-20

* Branch 51
Rabr51 node_4 netRa51 -879765.6723762706
Lbr51 netRa51 netL51 -8.369719786173988e-11
Rbbr51 netL51 0 899160.9856336433
Cbr51 netL51 0 -1.0594319680163885e-22

* Branch 52
Rabr52 node_4 netRa52 -419388.7825890099
Lbr52 netRa52 netL52 5.735841044261531e-11
Rbbr52 netL52 0 434504.1098181054
Cbr52 netL52 0 3.142307671192001e-22

* Branch 53
Rabr53 node_4 netRa53 -21230.058819487662
Lbr53 netRa53 netL53 -1.0981872669439281e-11
Rbbr53 netL53 0 26598.59173493996
Cbr53 netL53 0 -1.9573302863944192e-20

* Branch 54
Rabr54 node_4 netRa54 -51281.99413896908
Lbr54 netRa54 netL54 1.7217361902675117e-11
Rbbr54 netL54 0 66977.63434151986
Cbr54 netL54 0 4.9923128350831615e-21

* Branch 55
Rabr55 node_4 netRa55 2193.536221040108
Lbr55 netRa55 netL55 7.329853208161114e-12
Rbbr55 netL55 0 -55697.68457042498
Cbr55 netL55 0 6.253139034228073e-20

* Branch 56
Rabr56 node_4 netRa56 42754.650298636894
Lbr56 netRa56 netL56 2.2405328460595256e-11
Rbbr56 netL56 0 -66425.22759116592
Cbr56 netL56 0 7.938159782534159e-21

* Branch 57
Rabr57 node_4 netRa57 -22443.11720259371
Lbr57 netRa57 netL57 -1.9666269164272696e-11
Rbbr57 netL57 0 78460.45770946465
Cbr57 netL57 0 -1.1281830094048545e-20

* Branch 58
Rabr58 node_4 netRa58 12533.727020846787
Lbr58 netRa58 netL58 2.1094052674343014e-11
Rbbr58 netL58 0 -52508.034698770476
Cbr58 netL58 0 3.26796979008193e-20

* Branch 59
Rabr59 node_4 netRa59 238054.92059610086
Lbr59 netRa59 netL59 6.806221875602215e-11
Rbbr59 netL59 0 -264360.0323904482
Cbr59 netL59 0 1.0850042471231398e-21

* Branch 60
Rabr60 node_4 netRa60 4496.608334511572
Lbr60 netRa60 netL60 -3.431238653744719e-11
Rbbr60 netL60 0 -517282.83050749596
Cbr60 netL60 0 -1.3603268892424715e-20

* Branch 61
Rabr61 node_4 netRa61 -107438.77292430287
Lbr61 netRa61 netL61 4.018997013086564e-11
Rbbr61 netL61 0 129681.09492469356
Cbr61 netL61 0 2.8729330145909907e-21

* Branch 62
Rabr62 node_4 netRa62 -35404.076790169776
Lbr62 netRa62 netL62 1.4632498027248958e-11
Rbbr62 netL62 0 38108.21822100449
Cbr62 netL62 0 1.0797282795004548e-20

* Branch 63
Rabr63 node_4 netRa63 -64952.567719276405
Lbr63 netRa63 netL63 2.9094566513638744e-11
Rbbr63 netL63 0 79941.31779522709
Cbr63 netL63 0 5.5764562252495126e-21

* Branch 64
Rabr64 node_4 netRa64 1255.3995119624358
Lbr64 netRa64 netL64 1.458747353062083e-11
Rbbr64 netL64 0 -275783.75691257766
Cbr64 netL64 0 4.761811538236182e-20

* Branch 65
Rabr65 node_4 netRa65 21031.023994646144
Lbr65 netRa65 netL65 -1.5631533730995015e-11
Rbbr65 netL65 0 -32864.426303699096
Cbr65 netL65 0 -2.2455667432059e-20

* Branch 66
Rabr66 node_4 netRa66 -1549.2297583901243
Lbr66 netRa66 netL66 6.95091327945037e-12
Rbbr66 netL66 0 30363.723032117254
Cbr66 netL66 0 1.4203788890918575e-19

* Branch 67
Rabr67 node_4 netRa67 21865.49362818384
Lbr67 netRa67 netL67 2.4598611120067192e-11
Rbbr67 netL67 0 -49573.51151406437
Cbr67 netL67 0 2.2890701710706348e-20

* Branch 68
Rabr68 node_4 netRa68 66492.1228549849
Lbr68 netRa68 netL68 -3.4582686461877554e-11
Rbbr68 netL68 0 -109329.86392133795
Cbr68 netL68 0 -4.738669806214553e-21

* Branch 69
Rabr69 node_4 netRa69 28376.943013653414
Lbr69 netRa69 netL69 -2.8986737776245375e-11
Rbbr69 netL69 0 -121364.13780868675
Cbr69 netL69 0 -8.353123853886388e-21

* Branch 70
Rabr70 node_4 netRa70 -2825.9778099138907
Lbr70 netRa70 netL70 1.4100126989759385e-11
Rbbr70 netL70 0 75690.12250204194
Cbr70 netL70 0 6.360281993295868e-20

* Branch 71
Rabr71 node_4 netRa71 -6084.428556783807
Lbr71 netRa71 netL71 1.772931220625962e-11
Rbbr71 netL71 0 76810.96552910603
Cbr71 netL71 0 3.718983658024498e-20

* Branch 72
Rabr72 node_4 netRa72 43858.790835005915
Lbr72 netRa72 netL72 2.4460579183433133e-11
Rbbr72 netL72 0 -52181.33382088737
Cbr72 netL72 0 1.0727897202357432e-20

* Branch 73
Rabr73 node_4 netRa73 265916.27854448836
Lbr73 netRa73 netL73 -7.740758035268489e-11
Rbbr73 netL73 0 -280060.9860779035
Cbr73 netL73 0 -1.0375020886975298e-21

* Branch 74
Rabr74 node_4 netRa74 4661.6957672572835
Lbr74 netRa74 netL74 -7.948682681937406e-12
Rbbr74 netL74 0 -46343.82574461143
Cbr74 netL74 0 -3.6435137773671986e-20

* Branch 75
Rabr75 node_4 netRa75 16937.43422153307
Lbr75 netRa75 netL75 -1.554116226767728e-11
Rbbr75 netL75 0 -24025.985738992746
Cbr75 netL75 0 -3.800400863013686e-20

* Branch 76
Rabr76 node_4 netRa76 35660.24750001943
Lbr76 netRa76 netL76 -2.0559750706713304e-11
Rbbr76 netL76 0 -45728.717126199655
Cbr76 netL76 0 -1.2573083797782451e-20

* Branch 77
Rabr77 node_4 netRa77 -77371.6360715283
Lbr77 netRa77 netL77 3.175562680847532e-11
Rbbr77 netL77 0 106827.96298282339
Cbr77 netL77 0 3.83450416418799e-21

* Branch 78
Rabr78 node_4 netRa78 15178.019132857455
Lbr78 netRa78 netL78 -1.4591883445492636e-11
Rbbr78 netL78 0 -27543.91087262819
Cbr78 netL78 0 -3.4755320541294923e-20

* Branch 79
Rabr79 node_4 netRa79 -466751.8128261811
Lbr79 netRa79 netL79 6.945402107355461e-11
Rbbr79 netL79 0 487101.20570374344
Cbr79 netL79 0 3.0531744314566126e-22

* Branch 80
Rabr80 node_4 netRa80 9905808.586125344
Lbr80 netRa80 netL80 2.5285402200854355e-10
Rbbr80 netL80 0 -9910499.67440356
Cbr80 netL80 0 2.5758780082433907e-24

* Branch 81
Rabr81 node_4 netRa81 13855.495387134326
Lbr81 netRa81 netL81 1.3443505758215308e-11
Rbbr81 netL81 0 -21606.186414023723
Cbr81 netL81 0 4.506715876995093e-20

* Branch 82
Rabr82 node_4 netRa82 -210124.0115425735
Lbr82 netRa82 netL82 -5.770738078914535e-11
Rbbr82 netL82 0 244597.37503251727
Cbr82 netL82 0 -1.123912292801167e-21

* Branch 83
Rabr83 node_4 netRa83 14768.320954426696
Lbr83 netRa83 netL83 3.8173971794269804e-11
Rbbr83 netL83 0 -91544.8868130036
Cbr83 netL83 0 2.844957573249831e-20

* Branch 84
Rabr84 node_4 netRa84 12295.40974668843
Lbr84 netRa84 netL84 -1.2322158408223876e-11
Rbbr84 netL84 0 -23571.74878038637
Cbr84 netL84 0 -4.239964629037699e-20

* Branch 85
Rabr85 node_4 netRa85 -57725.41052199303
Lbr85 netRa85 netL85 -3.01681517364931e-11
Rbbr85 netL85 0 89604.68054781794
Cbr85 netL85 0 -5.840650544536636e-21

* Branch 86
Rabr86 node_4 netRa86 -9812.347921766219
Lbr86 netRa86 netL86 -1.4183312777439214e-11
Rbbr86 netL86 0 72571.99760213151
Cbr86 netL86 0 -1.9975147614330152e-20

* Branch 87
Rabr87 node_4 netRa87 -2182396.6602932015
Lbr87 netRa87 netL87 -2.621636905453018e-10
Rbbr87 netL87 0 2247418.2200013194
Cbr87 netL87 0 -5.3461563385667e-23

* Branch 88
Rabr88 node_4 netRa88 57039.37855761017
Lbr88 netRa88 netL88 -4.22842155699699e-11
Rbbr88 netL88 0 -73446.75893469203
Cbr88 netL88 0 -1.0088098492217338e-20

* Branch 89
Rabr89 node_4 netRa89 -66056.25859530955
Lbr89 netRa89 netL89 6.651989631598042e-11
Rbbr89 netL89 0 214628.90122965194
Cbr89 netL89 0 4.689295539308462e-21

* Branch 90
Rabr90 node_4 netRa90 12536824.25982155
Lbr90 netRa90 netL90 6.109239218492826e-10
Rbbr90 netL90 0 -12553478.221591031
Cbr90 netL90 0 3.881889230210436e-24

* Branch 91
Rabr91 node_4 netRa91 27510.0506560281
Lbr91 netRa91 netL91 -2.0145482539347498e-11
Rbbr91 netL91 0 -34603.05317904223
Cbr91 netL91 0 -2.115792527770017e-20

* Branch 92
Rabr92 node_4 netRa92 29558.911837019587
Lbr92 netRa92 netL92 2.00493080813763e-11
Rbbr92 netL92 0 -40433.37316716726
Cbr92 netL92 0 1.6795446220680614e-20

* Branch 93
Rabr93 node_4 netRa93 -7023.115190768252
Lbr93 netRa93 netL93 -3.880927722794312e-11
Rbbr93 netL93 0 102602.98693754563
Cbr93 netL93 0 -5.483496136586425e-20

* Branch 94
Rabr94 node_4 netRa94 193407.12484489483
Lbr94 netRa94 netL94 3.769236154993731e-11
Rbbr94 netL94 0 -199448.83053053642
Cbr94 netL94 0 9.782165730422935e-22

* Branch 95
Rabr95 node_4 netRa95 3896.10762464434
Lbr95 netRa95 netL95 -6.8637601085153925e-12
Rbbr95 netL95 0 -11072.198845395047
Cbr95 netL95 0 -1.5718077093787152e-19

* Branch 96
Rabr96 node_4 netRa96 -692.8988680765785
Lbr96 netRa96 netL96 6.622425726433268e-12
Rbbr96 netL96 0 42055.16311251523
Cbr96 netL96 0 2.079443663440712e-19

* Branch 97
Rabr97 node_4 netRa97 134907.61524519167
Lbr97 netRa97 netL97 2.6827534579618972e-11
Rbbr97 netL97 0 -137349.93949048597
Cbr97 netL97 0 1.4510642472752264e-21

* Branch 98
Rabr98 node_4 netRa98 -5537.440199654416
Lbr98 netRa98 netL98 1.6444840277860103e-11
Rbbr98 netL98 0 26979.67728144098
Cbr98 netL98 0 9.95212469572332e-20

* Branch 99
Rabr99 node_4 netRa99 59410.06410167461
Lbr99 netRa99 netL99 1.1520976674682975e-11
Rbbr99 netL99 0 -67480.18384197226
Cbr99 netL99 0 2.9337773577211572e-21

.ends


.end
